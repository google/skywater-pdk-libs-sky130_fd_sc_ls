* File: sky130_fd_sc_ls__sdfrbp_1.pxi.spice
* Created: Wed Sep  2 11:26:54 2020
* 
x_PM_SKY130_FD_SC_LS__SDFRBP_1%A_27_74# N_A_27_74#_M1032_s N_A_27_74#_M1026_s
+ N_A_27_74#_M1008_g N_A_27_74#_c_304_n N_A_27_74#_M1019_g N_A_27_74#_c_299_n
+ N_A_27_74#_c_300_n N_A_27_74#_c_301_n N_A_27_74#_c_302_n N_A_27_74#_c_306_n
+ N_A_27_74#_c_303_n N_A_27_74#_c_307_n N_A_27_74#_c_308_n
+ PM_SKY130_FD_SC_LS__SDFRBP_1%A_27_74#
x_PM_SKY130_FD_SC_LS__SDFRBP_1%SCE N_SCE_M1032_g N_SCE_c_387_n N_SCE_c_388_n
+ N_SCE_M1026_g N_SCE_c_389_n N_SCE_c_390_n N_SCE_M1037_g N_SCE_M1022_g
+ N_SCE_c_376_n N_SCE_c_377_n N_SCE_c_378_n N_SCE_c_379_n N_SCE_c_380_n
+ N_SCE_c_381_n SCE SCE SCE N_SCE_c_382_n N_SCE_c_383_n N_SCE_c_384_n
+ N_SCE_c_385_n SCE N_SCE_c_386_n PM_SKY130_FD_SC_LS__SDFRBP_1%SCE
x_PM_SKY130_FD_SC_LS__SDFRBP_1%D N_D_M1012_g N_D_c_473_n N_D_c_477_n N_D_M1014_g
+ D N_D_c_474_n N_D_c_475_n PM_SKY130_FD_SC_LS__SDFRBP_1%D
x_PM_SKY130_FD_SC_LS__SDFRBP_1%SCD N_SCD_M1023_g N_SCD_M1016_g N_SCD_c_519_n
+ N_SCD_c_523_n SCD SCD N_SCD_c_521_n PM_SKY130_FD_SC_LS__SDFRBP_1%SCD
x_PM_SKY130_FD_SC_LS__SDFRBP_1%CLK N_CLK_c_560_n N_CLK_c_561_n N_CLK_c_562_n
+ N_CLK_M1025_g N_CLK_c_563_n N_CLK_M1024_g N_CLK_c_564_n N_CLK_c_569_n CLK
+ N_CLK_c_565_n N_CLK_c_566_n CLK PM_SKY130_FD_SC_LS__SDFRBP_1%CLK
x_PM_SKY130_FD_SC_LS__SDFRBP_1%A_1034_392# N_A_1034_392#_M1033_d
+ N_A_1034_392#_M1028_d N_A_1034_392#_c_642_n N_A_1034_392#_c_643_n
+ N_A_1034_392#_M1039_g N_A_1034_392#_c_621_n N_A_1034_392#_M1000_g
+ N_A_1034_392#_c_623_n N_A_1034_392#_M1020_g N_A_1034_392#_c_624_n
+ N_A_1034_392#_c_625_n N_A_1034_392#_c_645_n N_A_1034_392#_M1015_g
+ N_A_1034_392#_c_646_n N_A_1034_392#_c_626_n N_A_1034_392#_c_627_n
+ N_A_1034_392#_c_628_n N_A_1034_392#_c_629_n N_A_1034_392#_c_647_n
+ N_A_1034_392#_c_630_n N_A_1034_392#_c_631_n N_A_1034_392#_c_632_n
+ N_A_1034_392#_c_657_p N_A_1034_392#_c_687_p N_A_1034_392#_c_633_n
+ N_A_1034_392#_c_634_n N_A_1034_392#_c_635_n N_A_1034_392#_c_636_n
+ N_A_1034_392#_c_649_n N_A_1034_392#_c_637_n N_A_1034_392#_c_638_n
+ N_A_1034_392#_c_639_n N_A_1034_392#_c_640_n N_A_1034_392#_c_641_n
+ PM_SKY130_FD_SC_LS__SDFRBP_1%A_1034_392#
x_PM_SKY130_FD_SC_LS__SDFRBP_1%A_1367_93# N_A_1367_93#_M1030_d
+ N_A_1367_93#_M1040_d N_A_1367_93#_M1021_g N_A_1367_93#_M1034_g
+ N_A_1367_93#_c_839_n N_A_1367_93#_c_840_n N_A_1367_93#_c_841_n
+ N_A_1367_93#_c_842_n N_A_1367_93#_c_843_n N_A_1367_93#_c_844_n
+ N_A_1367_93#_c_845_n N_A_1367_93#_c_846_n
+ PM_SKY130_FD_SC_LS__SDFRBP_1%A_1367_93#
x_PM_SKY130_FD_SC_LS__SDFRBP_1%RESET_B N_RESET_B_M1036_g N_RESET_B_M1038_g
+ N_RESET_B_c_950_n N_RESET_B_c_951_n N_RESET_B_c_959_n N_RESET_B_c_960_n
+ N_RESET_B_M1011_g N_RESET_B_c_961_n N_RESET_B_M1004_g N_RESET_B_c_953_n
+ N_RESET_B_M1005_g N_RESET_B_M1027_g N_RESET_B_c_963_n N_RESET_B_c_955_n
+ N_RESET_B_c_956_n N_RESET_B_c_964_n N_RESET_B_c_965_n N_RESET_B_c_966_n
+ N_RESET_B_c_967_n N_RESET_B_c_968_n N_RESET_B_c_969_n RESET_B
+ N_RESET_B_c_971_n N_RESET_B_c_972_n N_RESET_B_c_973_n N_RESET_B_c_974_n
+ N_RESET_B_c_975_n N_RESET_B_c_957_n PM_SKY130_FD_SC_LS__SDFRBP_1%RESET_B
x_PM_SKY130_FD_SC_LS__SDFRBP_1%A_1234_119# N_A_1234_119#_M1035_d
+ N_A_1234_119#_M1039_d N_A_1234_119#_M1004_d N_A_1234_119#_M1030_g
+ N_A_1234_119#_c_1206_n N_A_1234_119#_M1040_g N_A_1234_119#_c_1207_n
+ N_A_1234_119#_c_1199_n N_A_1234_119#_c_1200_n N_A_1234_119#_c_1209_n
+ N_A_1234_119#_c_1210_n N_A_1234_119#_c_1201_n N_A_1234_119#_c_1202_n
+ N_A_1234_119#_c_1203_n N_A_1234_119#_c_1204_n N_A_1234_119#_c_1212_n
+ N_A_1234_119#_c_1281_n N_A_1234_119#_c_1213_n N_A_1234_119#_c_1214_n
+ N_A_1234_119#_c_1205_n PM_SKY130_FD_SC_LS__SDFRBP_1%A_1234_119#
x_PM_SKY130_FD_SC_LS__SDFRBP_1%A_835_98# N_A_835_98#_M1025_s N_A_835_98#_M1024_s
+ N_A_835_98#_c_1346_n N_A_835_98#_M1028_g N_A_835_98#_c_1336_n
+ N_A_835_98#_M1033_g N_A_835_98#_c_1347_n N_A_835_98#_c_1348_n
+ N_A_835_98#_c_1349_n N_A_835_98#_c_1337_n N_A_835_98#_c_1338_n
+ N_A_835_98#_M1035_g N_A_835_98#_M1010_g N_A_835_98#_c_1351_n
+ N_A_835_98#_c_1352_n N_A_835_98#_c_1353_n N_A_835_98#_M1013_g
+ N_A_835_98#_c_1339_n N_A_835_98#_c_1340_n N_A_835_98#_M1009_g
+ N_A_835_98#_c_1357_n N_A_835_98#_c_1363_n N_A_835_98#_c_1342_n
+ N_A_835_98#_c_1343_n N_A_835_98#_c_1344_n N_A_835_98#_c_1345_n
+ PM_SKY130_FD_SC_LS__SDFRBP_1%A_835_98#
x_PM_SKY130_FD_SC_LS__SDFRBP_1%A_2008_48# N_A_2008_48#_M1007_d
+ N_A_2008_48#_M1027_d N_A_2008_48#_M1003_g N_A_2008_48#_c_1516_n
+ N_A_2008_48#_c_1523_n N_A_2008_48#_c_1524_n N_A_2008_48#_M1017_g
+ N_A_2008_48#_c_1517_n N_A_2008_48#_c_1526_n N_A_2008_48#_c_1527_n
+ N_A_2008_48#_c_1528_n N_A_2008_48#_c_1529_n N_A_2008_48#_c_1518_n
+ N_A_2008_48#_c_1530_n N_A_2008_48#_c_1519_n N_A_2008_48#_c_1520_n
+ N_A_2008_48#_c_1532_n N_A_2008_48#_c_1521_n
+ PM_SKY130_FD_SC_LS__SDFRBP_1%A_2008_48#
x_PM_SKY130_FD_SC_LS__SDFRBP_1%A_1747_74# N_A_1747_74#_M1020_d
+ N_A_1747_74#_M1013_d N_A_1747_74#_c_1651_n N_A_1747_74#_M1007_g
+ N_A_1747_74#_c_1652_n N_A_1747_74#_c_1653_n N_A_1747_74#_c_1663_n
+ N_A_1747_74#_M1041_g N_A_1747_74#_c_1664_n N_A_1747_74#_c_1665_n
+ N_A_1747_74#_M1002_g N_A_1747_74#_c_1654_n N_A_1747_74#_M1006_g
+ N_A_1747_74#_c_1655_n N_A_1747_74#_c_1656_n N_A_1747_74#_c_1668_n
+ N_A_1747_74#_c_1669_n N_A_1747_74#_M1029_g N_A_1747_74#_M1001_g
+ N_A_1747_74#_c_1670_n N_A_1747_74#_c_1658_n N_A_1747_74#_c_1678_n
+ N_A_1747_74#_c_1681_n N_A_1747_74#_c_1672_n N_A_1747_74#_c_1673_n
+ N_A_1747_74#_c_1659_n N_A_1747_74#_c_1660_n N_A_1747_74#_c_1661_n
+ N_A_1747_74#_c_1662_n PM_SKY130_FD_SC_LS__SDFRBP_1%A_1747_74#
x_PM_SKY130_FD_SC_LS__SDFRBP_1%A_2513_424# N_A_2513_424#_M1001_s
+ N_A_2513_424#_M1029_s N_A_2513_424#_M1031_g N_A_2513_424#_c_1832_n
+ N_A_2513_424#_M1018_g N_A_2513_424#_c_1833_n N_A_2513_424#_c_1837_n
+ N_A_2513_424#_c_1834_n N_A_2513_424#_c_1835_n
+ PM_SKY130_FD_SC_LS__SDFRBP_1%A_2513_424#
x_PM_SKY130_FD_SC_LS__SDFRBP_1%VPWR N_VPWR_M1026_d N_VPWR_M1023_d N_VPWR_M1024_d
+ N_VPWR_M1034_d N_VPWR_M1040_s N_VPWR_M1017_d N_VPWR_M1041_d N_VPWR_M1029_d
+ N_VPWR_c_1882_n N_VPWR_c_1883_n N_VPWR_c_1884_n N_VPWR_c_1885_n
+ N_VPWR_c_1886_n N_VPWR_c_1887_n N_VPWR_c_1888_n N_VPWR_c_1998_n
+ N_VPWR_c_1889_n N_VPWR_c_1890_n N_VPWR_c_1891_n N_VPWR_c_1892_n
+ N_VPWR_c_1893_n N_VPWR_c_1894_n N_VPWR_c_1895_n N_VPWR_c_1896_n VPWR
+ N_VPWR_c_1897_n N_VPWR_c_1898_n N_VPWR_c_1899_n N_VPWR_c_1900_n
+ N_VPWR_c_1901_n N_VPWR_c_1902_n N_VPWR_c_1881_n N_VPWR_c_1904_n
+ N_VPWR_c_1905_n N_VPWR_c_1906_n N_VPWR_c_1907_n N_VPWR_c_1908_n
+ PM_SKY130_FD_SC_LS__SDFRBP_1%VPWR
x_PM_SKY130_FD_SC_LS__SDFRBP_1%A_409_81# N_A_409_81#_M1012_d N_A_409_81#_M1035_s
+ N_A_409_81#_M1014_d N_A_409_81#_M1038_d N_A_409_81#_M1039_s
+ N_A_409_81#_c_2085_n N_A_409_81#_c_2067_n N_A_409_81#_c_2107_n
+ N_A_409_81#_c_2068_n N_A_409_81#_c_2076_n N_A_409_81#_c_2077_n
+ N_A_409_81#_c_2078_n N_A_409_81#_c_2069_n N_A_409_81#_c_2070_n
+ N_A_409_81#_c_2079_n N_A_409_81#_c_2071_n N_A_409_81#_c_2072_n
+ N_A_409_81#_c_2080_n N_A_409_81#_c_2081_n N_A_409_81#_c_2073_n
+ N_A_409_81#_c_2083_n N_A_409_81#_c_2074_n N_A_409_81#_c_2116_n
+ N_A_409_81#_c_2084_n PM_SKY130_FD_SC_LS__SDFRBP_1%A_409_81#
x_PM_SKY130_FD_SC_LS__SDFRBP_1%Q_N N_Q_N_M1006_d N_Q_N_M1002_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N PM_SKY130_FD_SC_LS__SDFRBP_1%Q_N
x_PM_SKY130_FD_SC_LS__SDFRBP_1%Q N_Q_M1031_d N_Q_M1018_d Q Q Q Q Q Q Q
+ N_Q_c_2265_n PM_SKY130_FD_SC_LS__SDFRBP_1%Q
x_PM_SKY130_FD_SC_LS__SDFRBP_1%VGND N_VGND_M1032_d N_VGND_M1036_d N_VGND_M1025_d
+ N_VGND_M1011_d N_VGND_M1003_d N_VGND_M1006_s N_VGND_M1001_d N_VGND_c_2283_n
+ N_VGND_c_2284_n N_VGND_c_2285_n N_VGND_c_2286_n N_VGND_c_2287_n
+ N_VGND_c_2288_n N_VGND_c_2289_n N_VGND_c_2290_n VGND N_VGND_c_2291_n
+ N_VGND_c_2292_n N_VGND_c_2293_n N_VGND_c_2294_n N_VGND_c_2295_n
+ N_VGND_c_2296_n N_VGND_c_2297_n N_VGND_c_2298_n N_VGND_c_2299_n
+ N_VGND_c_2300_n N_VGND_c_2301_n N_VGND_c_2302_n N_VGND_c_2303_n
+ PM_SKY130_FD_SC_LS__SDFRBP_1%VGND
x_PM_SKY130_FD_SC_LS__SDFRBP_1%noxref_25 N_noxref_25_M1008_s N_noxref_25_M1016_d
+ N_noxref_25_c_2421_n N_noxref_25_c_2422_n N_noxref_25_c_2423_n
+ N_noxref_25_c_2424_n PM_SKY130_FD_SC_LS__SDFRBP_1%noxref_25
cc_1 VNB N_A_27_74#_M1008_g 0.0249134f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_2 VNB N_A_27_74#_c_299_n 0.0280153f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_3 VNB N_A_27_74#_c_300_n 0.0167958f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.05
cc_4 VNB N_A_27_74#_c_301_n 0.0201543f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_5 VNB N_A_27_74#_c_302_n 0.0460387f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_6 VNB N_A_27_74#_c_303_n 0.018224f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.145
cc_7 VNB N_SCE_M1032_g 0.0718805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_SCE_c_376_n 0.00457743f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.145
cc_9 VNB N_SCE_c_377_n 0.0145309f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_10 VNB N_SCE_c_378_n 0.0106899f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_11 VNB N_SCE_c_379_n 0.0120788f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_12 VNB N_SCE_c_380_n 0.00504066f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.135
cc_13 VNB N_SCE_c_381_n 0.0294595f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.145
cc_14 VNB N_SCE_c_382_n 0.0181262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_SCE_c_383_n 0.0212614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_SCE_c_384_n 0.0117716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_SCE_c_385_n 0.00943038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_SCE_c_386_n 0.001771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_D_M1012_g 0.0189319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_D_c_473_n 0.0243074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_D_c_474_n 0.0348012f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_22 VNB N_D_c_475_n 0.00645951f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.98
cc_23 VNB N_SCD_M1016_g 0.0413981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_SCD_c_519_n 0.00371437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB SCD 0.00358981f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_26 VNB N_SCD_c_521_n 0.0154984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_CLK_c_560_n 0.0269396f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_28 VNB N_CLK_c_561_n 0.0142627f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=2.32
cc_29 VNB N_CLK_c_562_n 0.0155002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_CLK_c_563_n 0.00452949f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.98
cc_31 VNB N_CLK_c_564_n 0.00972297f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_32 VNB N_CLK_c_565_n 0.0411335f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.31
cc_33 VNB N_CLK_c_566_n 0.00603566f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.05
cc_34 VNB CLK 0.00675705f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_35 VNB N_A_1034_392#_c_621_n 0.0113969f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_36 VNB N_A_1034_392#_M1000_g 0.0378998f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_37 VNB N_A_1034_392#_c_623_n 0.0165921f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.31
cc_38 VNB N_A_1034_392#_c_624_n 0.0218458f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_39 VNB N_A_1034_392#_c_625_n 0.007436f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_40 VNB N_A_1034_392#_c_626_n 0.00991314f $X=-0.19 $Y=-0.245 $X2=2.53
+ $Y2=1.995
cc_41 VNB N_A_1034_392#_c_627_n 6.30651e-19 $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_42 VNB N_A_1034_392#_c_628_n 0.0329865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1034_392#_c_629_n 0.00321642f $X=-0.19 $Y=-0.245 $X2=2.53
+ $Y2=2.135
cc_44 VNB N_A_1034_392#_c_630_n 0.00171326f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.98
cc_45 VNB N_A_1034_392#_c_631_n 0.00375765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1034_392#_c_632_n 8.50976e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1034_392#_c_633_n 0.00661626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1034_392#_c_634_n 0.00224396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1034_392#_c_635_n 0.00148299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1034_392#_c_636_n 0.0026896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1034_392#_c_637_n 4.42537e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1034_392#_c_638_n 0.00766144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1034_392#_c_639_n 0.0334285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1034_392#_c_640_n 0.00544115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1034_392#_c_641_n 0.0114218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1367_93#_M1021_g 0.030989f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_57 VNB N_A_1367_93#_c_839_n 0.00389529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1367_93#_c_840_n 0.0235983f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.31
cc_59 VNB N_A_1367_93#_c_841_n 4.58327e-19 $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_60 VNB N_A_1367_93#_c_842_n 0.00227583f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_61 VNB N_A_1367_93#_c_843_n 0.00765404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1367_93#_c_844_n 0.00268284f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.135
cc_63 VNB N_A_1367_93#_c_845_n 0.00673626f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.512
cc_64 VNB N_A_1367_93#_c_846_n 0.00219559f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.995
cc_65 VNB N_RESET_B_M1036_g 0.0468959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_RESET_B_c_950_n 0.272222f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_67 VNB N_RESET_B_c_951_n 0.012806f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_68 VNB N_RESET_B_M1011_g 0.0265319f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_69 VNB N_RESET_B_c_953_n 0.018981f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.145
cc_70 VNB N_RESET_B_M1005_g 0.0341606f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_71 VNB N_RESET_B_c_955_n 0.0294537f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=2.135
cc_72 VNB N_RESET_B_c_956_n 0.0234009f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_73 VNB N_RESET_B_c_957_n 0.0158526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1234_119#_M1030_g 0.0272516f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_75 VNB N_A_1234_119#_c_1199_n 0.0028857f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.145
cc_76 VNB N_A_1234_119#_c_1200_n 0.00422204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1234_119#_c_1201_n 6.72487e-19 $X=-0.19 $Y=-0.245 $X2=0.89
+ $Y2=2.512
cc_78 VNB N_A_1234_119#_c_1202_n 0.00192123f $X=-0.19 $Y=-0.245 $X2=2.53
+ $Y2=1.995
cc_79 VNB N_A_1234_119#_c_1203_n 0.00653818f $X=-0.19 $Y=-0.245 $X2=2.5
+ $Y2=1.995
cc_80 VNB N_A_1234_119#_c_1204_n 0.00301796f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.145
cc_81 VNB N_A_1234_119#_c_1205_n 0.0401207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_835_98#_c_1336_n 0.0155098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_835_98#_c_1337_n 0.0316811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_835_98#_c_1338_n 0.0159407f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.05
cc_85 VNB N_A_835_98#_c_1339_n 0.0216126f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_86 VNB N_A_835_98#_c_1340_n 0.00443907f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_87 VNB N_A_835_98#_M1009_g 0.0503748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_835_98#_c_1342_n 0.00128593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_835_98#_c_1343_n 0.00385897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_835_98#_c_1344_n 0.00150962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_835_98#_c_1345_n 0.0545089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2008_48#_M1003_g 0.0424527f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_93 VNB N_A_2008_48#_c_1516_n 0.0184816f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.245
cc_94 VNB N_A_2008_48#_c_1517_n 0.00245359f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.31
cc_95 VNB N_A_2008_48#_c_1518_n 0.00907094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_2008_48#_c_1519_n 6.5078e-19 $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.512
cc_97 VNB N_A_2008_48#_c_1520_n 0.00160142f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_98 VNB N_A_2008_48#_c_1521_n 0.00658078f $X=-0.19 $Y=-0.245 $X2=2.53
+ $Y2=2.135
cc_99 VNB N_A_1747_74#_c_1651_n 0.0180751f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.98
cc_100 VNB N_A_1747_74#_c_1652_n 0.031848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1747_74#_c_1653_n 0.0157622f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.245
cc_102 VNB N_A_1747_74#_c_1654_n 0.0240396f $X=-0.19 $Y=-0.245 $X2=0.365
+ $Y2=1.145
cc_103 VNB N_A_1747_74#_c_1655_n 0.0485723f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.145
cc_104 VNB N_A_1747_74#_c_1656_n 0.0663668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1747_74#_M1001_g 0.0405544f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.512
cc_106 VNB N_A_1747_74#_c_1658_n 0.00927852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1747_74#_c_1659_n 0.00242934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1747_74#_c_1660_n 0.00130137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1747_74#_c_1661_n 0.0147798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_1747_74#_c_1662_n 0.020816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_2513_424#_M1031_g 0.0280908f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.615
cc_112 VNB N_A_2513_424#_c_1832_n 0.0352088f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.245
cc_113 VNB N_A_2513_424#_c_1833_n 0.0126466f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=0.58
cc_114 VNB N_A_2513_424#_c_1834_n 0.00835153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2513_424#_c_1835_n 4.48326e-19 $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=1.145
cc_116 VNB N_VPWR_c_1881_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_409_81#_c_2067_n 0.0224999f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.31
cc_118 VNB N_A_409_81#_c_2068_n 0.00429144f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.145
cc_119 VNB N_A_409_81#_c_2069_n 9.90482e-19 $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.512
cc_120 VNB N_A_409_81#_c_2070_n 0.00159941f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_121 VNB N_A_409_81#_c_2071_n 0.00510468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_409_81#_c_2072_n 0.00161453f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.145
cc_123 VNB N_A_409_81#_c_2073_n 0.0025068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_409_81#_c_2074_n 0.00442165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB Q_N 0.0123064f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.98
cc_126 VNB Q 0.0267037f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_127 VNB Q 0.0127641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_Q_c_2265_n 0.0251085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2283_n 0.0135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2284_n 0.0123151f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.512
cc_131 VNB N_VGND_c_2285_n 0.0124127f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.512
cc_132 VNB N_VGND_c_2286_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2287_n 0.0363017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2288_n 0.0097163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2289_n 0.0217694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2290_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2291_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2292_n 0.0636389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2293_n 0.0552549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2294_n 0.060941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2295_n 0.0284194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2296_n 0.0193554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2297_n 0.727914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2298_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2299_n 0.0038619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2300_n 0.0140821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2301_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2302_n 0.0153005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2303_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_noxref_25_c_2421_n 0.00349162f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.615
cc_151 VNB N_noxref_25_c_2422_n 0.0131102f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.245
cc_152 VNB N_noxref_25_c_2423_n 0.0039073f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_153 VNB N_noxref_25_c_2424_n 0.00408915f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.64
cc_154 VPB N_A_27_74#_c_304_n 0.0501659f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.245
cc_155 VPB N_A_27_74#_c_300_n 0.0237442f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.05
cc_156 VPB N_A_27_74#_c_306_n 0.0219674f $X=-0.19 $Y=1.66 $X2=2.365 $Y2=2.135
cc_157 VPB N_A_27_74#_c_307_n 0.064305f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.512
cc_158 VPB N_A_27_74#_c_308_n 0.00653951f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_159 VPB N_SCE_c_387_n 0.021095f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_SCE_c_388_n 0.0272472f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_161 VPB N_SCE_c_389_n 0.0141937f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.245
cc_162 VPB N_SCE_c_390_n 0.0211539f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_163 VPB N_SCE_c_376_n 0.0130807f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.145
cc_164 VPB N_SCE_c_380_n 0.00304854f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.135
cc_165 VPB N_SCE_c_382_n 0.0215244f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_SCE_c_383_n 0.0217946f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_SCE_c_386_n 0.00321268f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_D_c_473_n 0.0303197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_D_c_477_n 0.0214973f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_170 VPB N_SCD_c_519_n 0.0318475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_SCD_c_523_n 0.0328892f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.245
cc_172 VPB SCD 0.00353896f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_173 VPB N_CLK_c_563_n 0.00946373f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_174 VPB N_CLK_c_569_n 0.0254998f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_175 VPB N_A_1034_392#_c_642_n 0.0152883f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_176 VPB N_A_1034_392#_c_643_n 0.0194827f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_177 VPB N_A_1034_392#_c_621_n 0.012785f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_178 VPB N_A_1034_392#_c_645_n 0.0616091f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_179 VPB N_A_1034_392#_c_646_n 0.00243629f $X=-0.19 $Y=1.66 $X2=1.055
+ $Y2=2.135
cc_180 VPB N_A_1034_392#_c_647_n 0.00144418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_1034_392#_c_630_n 0.0019321f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_182 VPB N_A_1034_392#_c_649_n 0.00535343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_1034_392#_c_641_n 0.0175819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1367_93#_M1034_g 0.0381305f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_185 VPB N_A_1367_93#_c_839_n 0.00183672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1367_93#_c_840_n 0.0212319f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.31
cc_187 VPB N_A_1367_93#_c_844_n 0.00432622f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.135
cc_188 VPB N_RESET_B_M1036_g 0.0077857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_RESET_B_c_959_n 0.0402652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_RESET_B_c_960_n 0.0302463f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.245
cc_191 VPB N_RESET_B_c_961_n 0.017445f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_192 VPB N_RESET_B_c_953_n 0.00842104f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.145
cc_193 VPB N_RESET_B_c_963_n 0.0216309f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_194 VPB N_RESET_B_c_964_n 0.0117494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_RESET_B_c_965_n 0.0274905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_RESET_B_c_966_n 0.0180958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_RESET_B_c_967_n 0.00158938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_RESET_B_c_968_n 0.0138407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_RESET_B_c_969_n 0.0117419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB RESET_B 0.00207862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_RESET_B_c_971_n 0.00810558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_RESET_B_c_972_n 0.0686527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_RESET_B_c_973_n 0.00775347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_RESET_B_c_974_n 0.0307002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_RESET_B_c_975_n 0.0048181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_RESET_B_c_957_n 0.00104493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_1234_119#_c_1206_n 0.0164664f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.98
cc_208 VPB N_A_1234_119#_c_1207_n 0.00486281f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_1234_119#_c_1200_n 0.00354403f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_1234_119#_c_1209_n 0.00182206f $X=-0.19 $Y=1.66 $X2=1.055
+ $Y2=2.135
cc_211 VPB N_A_1234_119#_c_1210_n 0.00814204f $X=-0.19 $Y=1.66 $X2=0.24
+ $Y2=1.145
cc_212 VPB N_A_1234_119#_c_1201_n 0.00255881f $X=-0.19 $Y=1.66 $X2=0.89
+ $Y2=2.512
cc_213 VPB N_A_1234_119#_c_1212_n 8.22498e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1234_119#_c_1213_n 0.00316104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_1234_119#_c_1214_n 0.00122086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1234_119#_c_1205_n 0.0234566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_835_98#_c_1346_n 0.0162235f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_218 VPB N_A_835_98#_c_1347_n 0.0722913f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.98
cc_219 VPB N_A_835_98#_c_1348_n 0.0567222f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.58
cc_220 VPB N_A_835_98#_c_1349_n 0.0123764f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_221 VPB N_A_835_98#_M1010_g 0.0386451f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_835_98#_c_1351_n 0.186472f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.135
cc_223 VPB N_A_835_98#_c_1352_n 0.00753678f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.512
cc_224 VPB N_A_835_98#_c_1353_n 0.0145726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_835_98#_M1013_g 0.00889026f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_226 VPB N_A_835_98#_c_1339_n 0.0212414f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_227 VPB N_A_835_98#_c_1340_n 0.00362133f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_228 VPB N_A_835_98#_c_1357_n 0.00749069f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_229 VPB N_A_835_98#_c_1344_n 0.00872141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_835_98#_c_1345_n 0.028132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_2008_48#_c_1516_n 0.0363084f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.245
cc_232 VPB N_A_2008_48#_c_1523_n 0.0157644f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_233 VPB N_A_2008_48#_c_1524_n 0.0216925f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_234 VPB N_A_2008_48#_c_1517_n 0.00554437f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.31
cc_235 VPB N_A_2008_48#_c_1526_n 0.00200572f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_236 VPB N_A_2008_48#_c_1527_n 0.00188008f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_237 VPB N_A_2008_48#_c_1528_n 0.0030033f $X=-0.19 $Y=1.66 $X2=2.365 $Y2=2.135
cc_238 VPB N_A_2008_48#_c_1529_n 0.00272239f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.512
cc_239 VPB N_A_2008_48#_c_1530_n 0.00910875f $X=-0.19 $Y=1.66 $X2=0.89 $Y2=2.465
cc_240 VPB N_A_2008_48#_c_1519_n 0.00102188f $X=-0.19 $Y=1.66 $X2=1.055
+ $Y2=2.512
cc_241 VPB N_A_2008_48#_c_1532_n 0.00510966f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_242 VPB N_A_1747_74#_c_1663_n 0.0156363f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_243 VPB N_A_1747_74#_c_1664_n 0.0266893f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_244 VPB N_A_1747_74#_c_1665_n 0.0200685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_1747_74#_c_1655_n 0.0295508f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_246 VPB N_A_1747_74#_c_1656_n 0.0208636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_1747_74#_c_1668_n 0.0185739f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.135
cc_248 VPB N_A_1747_74#_c_1669_n 0.0280061f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.145
cc_249 VPB N_A_1747_74#_c_1670_n 0.0189178f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_250 VPB N_A_1747_74#_c_1658_n 0.00103641f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_1747_74#_c_1672_n 0.00533426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_A_1747_74#_c_1673_n 0.00295698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_A_1747_74#_c_1660_n 0.00536747f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_A_2513_424#_c_1832_n 0.0293072f $X=-0.19 $Y=1.66 $X2=2.485
+ $Y2=2.245
cc_255 VPB N_A_2513_424#_c_1837_n 0.00679439f $X=-0.19 $Y=1.66 $X2=0.365
+ $Y2=1.145
cc_256 VPB N_VPWR_c_1882_n 0.00653637f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.145
cc_257 VPB N_VPWR_c_1883_n 0.00662228f $X=-0.19 $Y=1.66 $X2=0.89 $Y2=2.465
cc_258 VPB N_VPWR_c_1884_n 0.00396467f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_259 VPB N_VPWR_c_1885_n 0.0157581f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_260 VPB N_VPWR_c_1886_n 0.0177109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1887_n 0.0169757f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1888_n 0.0142672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1889_n 0.0141486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1890_n 0.0338628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1891_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1892_n 0.0352503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1893_n 0.00601569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1894_n 0.0551755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1895_n 0.00317016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1896_n 5.16032e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1897_n 0.0436019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1898_n 0.0270975f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1899_n 0.0505955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1900_n 0.020722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1901_n 0.0343043f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1902_n 0.0189057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1881_n 0.135885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1904_n 0.00614151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1905_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1906_n 0.0066101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_1907_n 0.00853483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_1908_n 0.00535984f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_409_81#_c_2068_n 0.00666589f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_284 VPB N_A_409_81#_c_2076_n 8.30015e-19 $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.135
cc_285 VPB N_A_409_81#_c_2077_n 0.00843413f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.145
cc_286 VPB N_A_409_81#_c_2078_n 0.00361747f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.512
cc_287 VPB N_A_409_81#_c_2079_n 0.00289353f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=2.135
cc_288 VPB N_A_409_81#_c_2080_n 0.00543975f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_289 VPB N_A_409_81#_c_2081_n 0.001897f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_290 VPB N_A_409_81#_c_2073_n 0.00484787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_291 VPB N_A_409_81#_c_2083_n 0.00256678f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_A_409_81#_c_2084_n 0.00836287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB Q_N 0.0164214f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_294 VPB Q 0.0100975f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.245
cc_295 VPB Q 0.0417421f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.512
cc_296 VPB N_Q_c_2265_n 0.00779891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 N_A_27_74#_c_299_n N_SCE_M1032_g 0.00834942f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_298 N_A_27_74#_c_300_n N_SCE_M1032_g 0.017345f $X=0.2 $Y=2.05 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_301_n N_SCE_M1032_g 0.0301676f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_302_n N_SCE_M1032_g 0.00651386f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_301 N_A_27_74#_c_306_n N_SCE_c_387_n 0.00485819f $X=2.365 $Y=2.135 $X2=0
+ $Y2=0
cc_302 N_A_27_74#_c_307_n N_SCE_c_387_n 0.00322075f $X=1.055 $Y=2.512 $X2=0
+ $Y2=0
cc_303 N_A_27_74#_c_306_n N_SCE_c_388_n 0.00822995f $X=2.365 $Y=2.135 $X2=0
+ $Y2=0
cc_304 N_A_27_74#_c_307_n N_SCE_c_388_n 0.014007f $X=1.055 $Y=2.512 $X2=0 $Y2=0
cc_305 N_A_27_74#_c_306_n N_SCE_c_389_n 0.00663467f $X=2.365 $Y=2.135 $X2=0
+ $Y2=0
cc_306 N_A_27_74#_c_306_n N_SCE_c_390_n 0.00943326f $X=2.365 $Y=2.135 $X2=0
+ $Y2=0
cc_307 N_A_27_74#_c_307_n N_SCE_c_390_n 7.55381e-19 $X=1.055 $Y=2.512 $X2=0
+ $Y2=0
cc_308 N_A_27_74#_c_307_n N_SCE_c_376_n 0.0185427f $X=1.055 $Y=2.512 $X2=0 $Y2=0
cc_309 N_A_27_74#_c_304_n N_SCE_c_379_n 5.18235e-19 $X=2.485 $Y=2.245 $X2=0
+ $Y2=0
cc_310 N_A_27_74#_c_306_n N_SCE_c_379_n 0.0226621f $X=2.365 $Y=2.135 $X2=0 $Y2=0
cc_311 N_A_27_74#_c_308_n N_SCE_c_379_n 0.00221846f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_312 N_A_27_74#_c_304_n N_SCE_c_380_n 9.36519e-19 $X=2.485 $Y=2.245 $X2=0
+ $Y2=0
cc_313 N_A_27_74#_c_308_n N_SCE_c_380_n 0.024597f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_314 N_A_27_74#_c_304_n N_SCE_c_381_n 0.0176236f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_315 N_A_27_74#_c_308_n N_SCE_c_381_n 3.89e-19 $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_316 N_A_27_74#_c_301_n N_SCE_c_382_n 0.00418014f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_317 N_A_27_74#_c_301_n N_SCE_c_383_n 3.70862e-19 $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_318 N_A_27_74#_c_302_n N_SCE_c_383_n 0.0219042f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_319 N_A_27_74#_c_306_n N_SCE_c_383_n 0.00313888f $X=2.365 $Y=2.135 $X2=0
+ $Y2=0
cc_320 N_A_27_74#_c_300_n N_SCE_c_385_n 0.0195247f $X=0.2 $Y=2.05 $X2=0 $Y2=0
cc_321 N_A_27_74#_c_301_n N_SCE_c_385_n 0.0626128f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_322 N_A_27_74#_c_302_n N_SCE_c_385_n 0.00563186f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_323 N_A_27_74#_c_307_n N_SCE_c_385_n 0.0467278f $X=1.055 $Y=2.512 $X2=0 $Y2=0
cc_324 N_A_27_74#_c_306_n N_SCE_c_386_n 0.0467278f $X=2.365 $Y=2.135 $X2=0 $Y2=0
cc_325 N_A_27_74#_c_308_n N_SCE_c_386_n 0.00165158f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_326 N_A_27_74#_M1008_g N_D_M1012_g 0.0255023f $X=1.485 $Y=0.615 $X2=0 $Y2=0
cc_327 N_A_27_74#_c_304_n N_D_c_473_n 0.0212855f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_328 N_A_27_74#_c_306_n N_D_c_473_n 0.00760671f $X=2.365 $Y=2.135 $X2=0 $Y2=0
cc_329 N_A_27_74#_c_308_n N_D_c_473_n 0.0013236f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_330 N_A_27_74#_c_304_n N_D_c_477_n 0.0137871f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_331 N_A_27_74#_c_306_n N_D_c_477_n 0.00916304f $X=2.365 $Y=2.135 $X2=0 $Y2=0
cc_332 N_A_27_74#_c_301_n N_D_c_474_n 2.658e-19 $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_333 N_A_27_74#_c_302_n N_D_c_474_n 0.0150607f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_334 N_A_27_74#_M1008_g N_D_c_475_n 0.00642636f $X=1.485 $Y=0.615 $X2=0 $Y2=0
cc_335 N_A_27_74#_c_301_n N_D_c_475_n 0.0286966f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_336 N_A_27_74#_c_302_n N_D_c_475_n 7.30413e-19 $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_337 N_A_27_74#_c_304_n N_SCD_c_519_n 0.0194764f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_338 N_A_27_74#_c_308_n N_SCD_c_519_n 0.00373007f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_339 N_A_27_74#_c_304_n N_SCD_c_523_n 0.0283894f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_340 N_A_27_74#_c_304_n SCD 3.55393e-19 $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_341 N_A_27_74#_c_308_n SCD 0.0195522f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_342 N_A_27_74#_c_306_n N_VPWR_c_1882_n 0.0234317f $X=2.365 $Y=2.135 $X2=0
+ $Y2=0
cc_343 N_A_27_74#_c_307_n N_VPWR_c_1882_n 0.0251436f $X=1.055 $Y=2.512 $X2=0
+ $Y2=0
cc_344 N_A_27_74#_c_304_n N_VPWR_c_1883_n 0.00124994f $X=2.485 $Y=2.245 $X2=0
+ $Y2=0
cc_345 N_A_27_74#_c_307_n N_VPWR_c_1890_n 0.0408917f $X=1.055 $Y=2.512 $X2=0
+ $Y2=0
cc_346 N_A_27_74#_c_304_n N_VPWR_c_1897_n 0.00294132f $X=2.485 $Y=2.245 $X2=0
+ $Y2=0
cc_347 N_A_27_74#_c_304_n N_VPWR_c_1881_n 0.00362058f $X=2.485 $Y=2.245 $X2=0
+ $Y2=0
cc_348 N_A_27_74#_c_307_n N_VPWR_c_1881_n 0.0345127f $X=1.055 $Y=2.512 $X2=0
+ $Y2=0
cc_349 N_A_27_74#_c_304_n N_A_409_81#_c_2085_n 0.00451918f $X=2.485 $Y=2.245
+ $X2=0 $Y2=0
cc_350 N_A_27_74#_c_308_n N_A_409_81#_c_2085_n 0.00895554f $X=2.5 $Y=1.995 $X2=0
+ $Y2=0
cc_351 N_A_27_74#_c_304_n N_A_409_81#_c_2083_n 0.0176784f $X=2.485 $Y=2.245
+ $X2=0 $Y2=0
cc_352 N_A_27_74#_c_306_n N_A_409_81#_c_2083_n 0.0187713f $X=2.365 $Y=2.135
+ $X2=0 $Y2=0
cc_353 N_A_27_74#_c_308_n N_A_409_81#_c_2083_n 0.0133567f $X=2.5 $Y=1.995 $X2=0
+ $Y2=0
cc_354 N_A_27_74#_M1008_g N_VGND_c_2283_n 0.00126524f $X=1.485 $Y=0.615 $X2=0
+ $Y2=0
cc_355 N_A_27_74#_c_299_n N_VGND_c_2283_n 0.0179429f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_356 N_A_27_74#_c_301_n N_VGND_c_2283_n 0.0288081f $X=1.23 $Y=1.145 $X2=0
+ $Y2=0
cc_357 N_A_27_74#_c_299_n N_VGND_c_2291_n 0.011066f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_358 N_A_27_74#_M1008_g N_VGND_c_2292_n 9.15902e-19 $X=1.485 $Y=0.615 $X2=0
+ $Y2=0
cc_359 N_A_27_74#_c_299_n N_VGND_c_2297_n 0.00915947f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_c_301_n N_noxref_25_c_2421_n 0.0201381f $X=1.23 $Y=1.145 $X2=0
+ $Y2=0
cc_361 N_A_27_74#_c_302_n N_noxref_25_c_2421_n 0.00573089f $X=1.23 $Y=1.145
+ $X2=0 $Y2=0
cc_362 N_A_27_74#_M1008_g N_noxref_25_c_2422_n 0.0158911f $X=1.485 $Y=0.615
+ $X2=0 $Y2=0
cc_363 N_SCE_c_377_n N_D_M1012_g 0.00880032f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_364 N_SCE_c_378_n N_D_M1012_g 0.00164308f $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_365 N_SCE_c_379_n N_D_c_473_n 0.0147903f $X=2.395 $Y=1.575 $X2=0 $Y2=0
cc_366 N_SCE_c_380_n N_D_c_473_n 3.10088e-19 $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_367 N_SCE_c_383_n N_D_c_473_n 0.0188435f $X=1.615 $Y=1.715 $X2=0 $Y2=0
cc_368 N_SCE_c_386_n N_D_c_473_n 0.00533998f $X=1.795 $Y=1.685 $X2=0 $Y2=0
cc_369 N_SCE_c_389_n N_D_c_477_n 0.0188435f $X=1.615 $Y=2.155 $X2=0 $Y2=0
cc_370 N_SCE_c_390_n N_D_c_477_n 0.0378156f $X=1.615 $Y=2.245 $X2=0 $Y2=0
cc_371 N_SCE_c_378_n N_D_c_474_n 0.00850567f $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_372 N_SCE_c_380_n N_D_c_474_n 0.00124809f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_373 N_SCE_c_381_n N_D_c_474_n 0.0202526f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_374 N_SCE_c_386_n N_D_c_474_n 0.00410294f $X=1.795 $Y=1.685 $X2=0 $Y2=0
cc_375 N_SCE_c_378_n N_D_c_475_n 2.90043e-19 $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_376 N_SCE_c_380_n N_D_c_475_n 0.0024647f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_377 N_SCE_c_383_n N_D_c_475_n 9.21412e-19 $X=1.615 $Y=1.715 $X2=0 $Y2=0
cc_378 N_SCE_c_384_n N_D_c_475_n 9.26106e-19 $X=2.51 $Y=1.26 $X2=0 $Y2=0
cc_379 N_SCE_c_385_n N_D_c_475_n 0.0411265f $X=1.6 $Y=1.685 $X2=0 $Y2=0
cc_380 N_SCE_c_377_n N_SCD_M1016_g 0.0408623f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_381 N_SCE_c_380_n N_SCD_M1016_g 0.00391172f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_382 N_SCE_c_384_n N_SCD_M1016_g 0.0171335f $X=2.51 $Y=1.26 $X2=0 $Y2=0
cc_383 N_SCE_c_380_n SCD 0.0148325f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_384 N_SCE_c_380_n N_SCD_c_521_n 0.00257809f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_385 N_SCE_c_381_n N_SCD_c_521_n 0.00936322f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_386 N_SCE_c_388_n N_VPWR_c_1882_n 0.00645742f $X=1.115 $Y=2.245 $X2=0 $Y2=0
cc_387 N_SCE_c_390_n N_VPWR_c_1882_n 0.013944f $X=1.615 $Y=2.245 $X2=0 $Y2=0
cc_388 N_SCE_c_388_n N_VPWR_c_1890_n 0.0044455f $X=1.115 $Y=2.245 $X2=0 $Y2=0
cc_389 N_SCE_c_390_n N_VPWR_c_1897_n 0.00413917f $X=1.615 $Y=2.245 $X2=0 $Y2=0
cc_390 N_SCE_c_388_n N_VPWR_c_1881_n 0.00858576f $X=1.115 $Y=2.245 $X2=0 $Y2=0
cc_391 N_SCE_c_390_n N_VPWR_c_1881_n 0.00817532f $X=1.615 $Y=2.245 $X2=0 $Y2=0
cc_392 N_SCE_c_378_n N_A_409_81#_c_2067_n 0.00703377f $X=2.625 $Y=1.05 $X2=0
+ $Y2=0
cc_393 N_SCE_c_380_n N_A_409_81#_c_2067_n 0.00943064f $X=2.51 $Y=1.425 $X2=0
+ $Y2=0
cc_394 N_SCE_c_384_n N_A_409_81#_c_2067_n 0.00186435f $X=2.51 $Y=1.26 $X2=0
+ $Y2=0
cc_395 N_SCE_c_390_n N_A_409_81#_c_2083_n 0.00169852f $X=1.615 $Y=2.245 $X2=0
+ $Y2=0
cc_396 N_SCE_c_377_n N_A_409_81#_c_2074_n 0.00655329f $X=2.625 $Y=0.9 $X2=0
+ $Y2=0
cc_397 N_SCE_c_378_n N_A_409_81#_c_2074_n 0.00469207f $X=2.625 $Y=1.05 $X2=0
+ $Y2=0
cc_398 N_SCE_c_379_n N_A_409_81#_c_2074_n 0.00543911f $X=2.395 $Y=1.575 $X2=0
+ $Y2=0
cc_399 N_SCE_c_380_n N_A_409_81#_c_2074_n 0.0166692f $X=2.51 $Y=1.425 $X2=0
+ $Y2=0
cc_400 N_SCE_c_381_n N_A_409_81#_c_2074_n 0.0023445f $X=2.51 $Y=1.425 $X2=0
+ $Y2=0
cc_401 N_SCE_c_384_n N_A_409_81#_c_2074_n 0.001913f $X=2.51 $Y=1.26 $X2=0 $Y2=0
cc_402 N_SCE_M1032_g N_VGND_c_2283_n 0.0141679f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_403 N_SCE_M1032_g N_VGND_c_2291_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_404 N_SCE_c_377_n N_VGND_c_2292_n 9.15902e-19 $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_405 N_SCE_M1032_g N_VGND_c_2297_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_406 N_SCE_M1032_g N_noxref_25_c_2421_n 7.01965e-19 $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_407 N_SCE_c_377_n N_noxref_25_c_2422_n 0.0118647f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_408 N_SCE_M1032_g N_noxref_25_c_2423_n 6.37214e-19 $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_409 N_SCE_c_377_n N_noxref_25_c_2424_n 0.001431f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_410 N_D_c_477_n N_VPWR_c_1882_n 0.00224533f $X=2.035 $Y=2.245 $X2=0 $Y2=0
cc_411 N_D_c_477_n N_VPWR_c_1897_n 0.00445602f $X=2.035 $Y=2.245 $X2=0 $Y2=0
cc_412 N_D_c_477_n N_VPWR_c_1881_n 0.00858241f $X=2.035 $Y=2.245 $X2=0 $Y2=0
cc_413 N_D_c_477_n N_A_409_81#_c_2083_n 0.0105215f $X=2.035 $Y=2.245 $X2=0 $Y2=0
cc_414 N_D_M1012_g N_A_409_81#_c_2074_n 0.00584318f $X=1.97 $Y=0.615 $X2=0 $Y2=0
cc_415 N_D_c_474_n N_A_409_81#_c_2074_n 9.34668e-19 $X=1.935 $Y=1.145 $X2=0
+ $Y2=0
cc_416 N_D_c_475_n N_A_409_81#_c_2074_n 0.0230366f $X=1.935 $Y=1.145 $X2=0 $Y2=0
cc_417 N_D_M1012_g N_VGND_c_2292_n 9.15902e-19 $X=1.97 $Y=0.615 $X2=0 $Y2=0
cc_418 N_D_M1012_g N_noxref_25_c_2422_n 0.012163f $X=1.97 $Y=0.615 $X2=0 $Y2=0
cc_419 N_D_c_474_n N_noxref_25_c_2422_n 0.00108727f $X=1.935 $Y=1.145 $X2=0
+ $Y2=0
cc_420 N_D_c_475_n N_noxref_25_c_2422_n 0.0130151f $X=1.935 $Y=1.145 $X2=0 $Y2=0
cc_421 N_D_c_475_n noxref_26 0.00349454f $X=1.935 $Y=1.145 $X2=-0.19 $Y2=-0.245
cc_422 N_SCD_M1016_g N_RESET_B_M1036_g 0.0329664f $X=3.04 $Y=0.615 $X2=0 $Y2=0
cc_423 SCD N_RESET_B_M1036_g 0.00426118f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_424 N_SCD_c_521_n N_RESET_B_M1036_g 0.0255354f $X=3.05 $Y=1.605 $X2=0 $Y2=0
cc_425 N_SCD_c_519_n N_RESET_B_c_960_n 0.0255354f $X=3.05 $Y=2.08 $X2=0 $Y2=0
cc_426 N_SCD_c_523_n N_RESET_B_c_963_n 0.01653f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_427 N_SCD_c_523_n N_VPWR_c_1883_n 0.00873254f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_428 N_SCD_c_523_n N_VPWR_c_1897_n 0.00413917f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_429 N_SCD_c_523_n N_VPWR_c_1881_n 0.00399549f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_430 N_SCD_M1016_g N_A_409_81#_c_2067_n 0.0123829f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_431 SCD N_A_409_81#_c_2067_n 0.0149154f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_432 N_SCD_c_521_n N_A_409_81#_c_2067_n 0.00251861f $X=3.05 $Y=1.605 $X2=0
+ $Y2=0
cc_433 N_SCD_c_523_n N_A_409_81#_c_2107_n 0.0159295f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_434 SCD N_A_409_81#_c_2107_n 0.0173868f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_435 N_SCD_M1016_g N_A_409_81#_c_2068_n 0.00207067f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_436 N_SCD_c_523_n N_A_409_81#_c_2068_n 0.00216808f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_437 SCD N_A_409_81#_c_2068_n 0.0513304f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_438 N_SCD_c_521_n N_A_409_81#_c_2068_n 7.83502e-19 $X=3.05 $Y=1.605 $X2=0
+ $Y2=0
cc_439 N_SCD_c_523_n N_A_409_81#_c_2077_n 0.00152026f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_440 N_SCD_c_523_n N_A_409_81#_c_2083_n 0.00179166f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_441 N_SCD_M1016_g N_A_409_81#_c_2074_n 0.00135432f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_442 N_SCD_c_523_n N_A_409_81#_c_2116_n 0.00219891f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_443 N_SCD_M1016_g N_VGND_c_2292_n 9.09315e-19 $X=3.04 $Y=0.615 $X2=0 $Y2=0
cc_444 N_SCD_M1016_g N_noxref_25_c_2422_n 0.00698763f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_445 N_SCD_M1016_g N_noxref_25_c_2424_n 0.01038f $X=3.04 $Y=0.615 $X2=0 $Y2=0
cc_446 N_CLK_c_569_n N_A_1034_392#_c_646_n 2.73677e-19 $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_447 N_CLK_c_562_n N_A_1034_392#_c_626_n 9.65742e-19 $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_448 N_CLK_c_565_n N_RESET_B_M1036_g 0.0424626f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_449 N_CLK_c_566_n N_RESET_B_M1036_g 0.00104889f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_450 N_CLK_c_562_n N_RESET_B_c_950_n 0.0100028f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_451 N_CLK_c_565_n N_RESET_B_c_950_n 0.0043433f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_452 N_CLK_c_566_n N_RESET_B_c_950_n 0.00333603f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_453 N_CLK_c_561_n N_RESET_B_c_959_n 0.021335f $X=4.115 $Y=1.515 $X2=0 $Y2=0
cc_454 N_CLK_c_569_n N_RESET_B_c_959_n 0.00545707f $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_455 N_CLK_c_566_n N_RESET_B_c_959_n 0.00108293f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_456 CLK N_RESET_B_c_966_n 0.00639226f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_457 N_CLK_c_566_n N_RESET_B_c_967_n 8.53947e-19 $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_458 CLK N_RESET_B_c_967_n 0.0034901f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_459 N_CLK_c_561_n N_RESET_B_c_971_n 7.9265e-19 $X=4.115 $Y=1.515 $X2=0 $Y2=0
cc_460 N_CLK_c_569_n N_RESET_B_c_971_n 4.10028e-19 $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_461 N_CLK_c_566_n N_RESET_B_c_971_n 0.0195969f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_462 CLK N_RESET_B_c_971_n 0.00715169f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_463 CLK N_A_835_98#_M1025_s 0.00276012f $X=4.08 $Y=1.295 $X2=-0.19 $Y2=-0.245
cc_464 N_CLK_c_569_n N_A_835_98#_c_1346_n 0.0374488f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_465 N_CLK_c_562_n N_A_835_98#_c_1336_n 0.0211093f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_466 N_CLK_c_562_n N_A_835_98#_c_1363_n 0.00842292f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_467 CLK N_A_835_98#_c_1363_n 0.00802204f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_468 N_CLK_c_562_n N_A_835_98#_c_1342_n 0.00571974f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_469 N_CLK_c_564_n N_A_835_98#_c_1342_n 3.29111e-19 $X=4.62 $Y=1.515 $X2=0
+ $Y2=0
cc_470 CLK N_A_835_98#_c_1342_n 0.0218249f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_471 N_CLK_c_560_n N_A_835_98#_c_1343_n 0.00102376f $X=4.52 $Y=1.515 $X2=0
+ $Y2=0
cc_472 N_CLK_c_562_n N_A_835_98#_c_1343_n 0.0156817f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_473 N_CLK_c_565_n N_A_835_98#_c_1343_n 5.73272e-19 $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_474 N_CLK_c_566_n N_A_835_98#_c_1343_n 0.00745903f $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_475 CLK N_A_835_98#_c_1343_n 0.0251408f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_476 N_CLK_c_560_n N_A_835_98#_c_1344_n 0.00136113f $X=4.52 $Y=1.515 $X2=0
+ $Y2=0
cc_477 N_CLK_c_564_n N_A_835_98#_c_1344_n 0.0058844f $X=4.62 $Y=1.515 $X2=0
+ $Y2=0
cc_478 N_CLK_c_569_n N_A_835_98#_c_1344_n 0.0205213f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_479 CLK N_A_835_98#_c_1344_n 0.0392481f $X=4.08 $Y=1.295 $X2=0 $Y2=0
cc_480 N_CLK_c_564_n N_A_835_98#_c_1345_n 0.0262256f $X=4.62 $Y=1.515 $X2=0
+ $Y2=0
cc_481 N_CLK_c_569_n N_VPWR_c_1884_n 0.0164315f $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_482 N_CLK_c_569_n N_VPWR_c_1892_n 0.00302783f $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_483 N_CLK_c_569_n N_VPWR_c_1881_n 0.00396658f $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_484 N_CLK_c_565_n N_A_409_81#_c_2067_n 8.58559e-19 $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_485 N_CLK_c_566_n N_A_409_81#_c_2067_n 0.0142806f $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_486 N_CLK_c_565_n N_A_409_81#_c_2068_n 0.0029155f $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_487 N_CLK_c_566_n N_A_409_81#_c_2068_n 0.0399925f $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_488 N_CLK_c_569_n N_A_409_81#_c_2076_n 0.0102356f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_489 N_CLK_c_569_n N_A_409_81#_c_2077_n 5.41016e-19 $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_490 N_CLK_c_569_n N_A_409_81#_c_2078_n 0.00644616f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_491 N_CLK_c_569_n N_A_409_81#_c_2084_n 0.00874826f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_492 N_CLK_c_562_n N_VGND_c_2284_n 0.00163608f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_493 N_CLK_c_565_n N_VGND_c_2284_n 4.3252e-19 $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_494 N_CLK_c_566_n N_VGND_c_2284_n 0.00861101f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_495 N_CLK_c_562_n N_VGND_c_2285_n 0.00235542f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_496 N_CLK_c_562_n N_VGND_c_2297_n 9.39239e-19 $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_497 N_A_1034_392#_c_633_n N_A_1367_93#_M1030_d 0.00187547f $X=8.825 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_498 N_A_1034_392#_M1000_g N_A_1367_93#_M1021_g 0.0333609f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_499 N_A_1034_392#_c_628_n N_A_1367_93#_M1021_g 0.00344795f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_500 N_A_1034_392#_c_631_n N_A_1367_93#_M1021_g 0.00262964f $X=7.135 $Y=0.58
+ $X2=0 $Y2=0
cc_501 N_A_1034_392#_c_657_p N_A_1367_93#_M1021_g 0.0026982f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_502 N_A_1034_392#_c_642_n N_A_1367_93#_M1034_g 0.00334209f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_503 N_A_1034_392#_c_641_n N_A_1367_93#_M1034_g 7.41525e-19 $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_504 N_A_1034_392#_c_621_n N_A_1367_93#_c_840_n 0.0333609f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_505 N_A_1034_392#_c_641_n N_A_1367_93#_c_840_n 0.00108114f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_506 N_A_1034_392#_c_628_n N_A_1367_93#_c_841_n 5.94333e-19 $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_507 N_A_1034_392#_c_632_n N_A_1367_93#_c_841_n 0.00304701f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_508 N_A_1034_392#_c_657_p N_A_1367_93#_c_841_n 0.0103944f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_509 N_A_1034_392#_c_625_n N_A_1367_93#_c_842_n 0.00579988f $X=8.735 $Y=1.16
+ $X2=0 $Y2=0
cc_510 N_A_1034_392#_c_636_n N_A_1367_93#_c_842_n 0.0051103f $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_511 N_A_1034_392#_c_625_n N_A_1367_93#_c_843_n 0.0102306f $X=8.735 $Y=1.16
+ $X2=0 $Y2=0
cc_512 N_A_1034_392#_c_636_n N_A_1367_93#_c_843_n 0.00847972f $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_513 N_A_1034_392#_c_638_n N_A_1367_93#_c_843_n 0.00827695f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_514 N_A_1034_392#_c_640_n N_A_1367_93#_c_843_n 0.00615816f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_515 N_A_1034_392#_c_649_n N_A_1367_93#_c_844_n 0.00513948f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_516 N_A_1034_392#_c_640_n N_A_1367_93#_c_844_n 0.0132001f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_517 N_A_1034_392#_c_632_n N_A_1367_93#_c_845_n 0.0560854f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_518 N_A_1034_392#_c_633_n N_A_1367_93#_c_845_n 0.00353238f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_519 N_A_1034_392#_c_623_n N_A_1367_93#_c_846_n 0.00883423f $X=8.66 $Y=1.085
+ $X2=0 $Y2=0
cc_520 N_A_1034_392#_c_625_n N_A_1367_93#_c_846_n 2.35907e-19 $X=8.735 $Y=1.16
+ $X2=0 $Y2=0
cc_521 N_A_1034_392#_c_633_n N_A_1367_93#_c_846_n 0.0195702f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_522 N_A_1034_392#_c_635_n N_A_1367_93#_c_846_n 0.0232075f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_523 N_A_1034_392#_c_636_n N_A_1367_93#_c_846_n 4.87277e-19 $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_524 N_A_1034_392#_c_638_n N_A_1367_93#_c_846_n 0.0146226f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_525 N_A_1034_392#_M1000_g N_RESET_B_c_950_n 0.00882199f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_526 N_A_1034_392#_c_628_n N_RESET_B_c_950_n 0.0294278f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_527 N_A_1034_392#_c_629_n N_RESET_B_c_950_n 0.00992957f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_528 N_A_1034_392#_c_628_n N_RESET_B_M1011_g 0.00466687f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_529 N_A_1034_392#_c_631_n N_RESET_B_M1011_g 0.00445709f $X=7.135 $Y=0.58
+ $X2=0 $Y2=0
cc_530 N_A_1034_392#_c_632_n N_RESET_B_M1011_g 0.0128168f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_531 N_A_1034_392#_c_687_p N_RESET_B_M1011_g 0.0035287f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_532 N_A_1034_392#_c_634_n N_RESET_B_M1011_g 6.46496e-19 $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_533 N_A_1034_392#_c_642_n N_RESET_B_c_966_n 0.00315542f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_534 N_A_1034_392#_c_621_n N_RESET_B_c_966_n 0.00325193f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_535 N_A_1034_392#_c_646_n N_RESET_B_c_966_n 0.0144304f $X=5.45 $Y=2.085 $X2=0
+ $Y2=0
cc_536 N_A_1034_392#_c_647_n N_RESET_B_c_966_n 0.017308f $X=5.63 $Y=1.71 $X2=0
+ $Y2=0
cc_537 N_A_1034_392#_c_630_n N_RESET_B_c_966_n 0.0155597f $X=6.085 $Y=1.71 $X2=0
+ $Y2=0
cc_538 N_A_1034_392#_c_641_n N_RESET_B_c_966_n 0.00379596f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_539 N_A_1034_392#_c_645_n N_RESET_B_c_968_n 0.0053373f $X=9.77 $Y=2.37 $X2=0
+ $Y2=0
cc_540 N_A_1034_392#_c_649_n N_RESET_B_c_968_n 0.0136948f $X=9.67 $Y=2.065 $X2=0
+ $Y2=0
cc_541 N_A_1034_392#_c_640_n N_RESET_B_c_968_n 0.0078678f $X=9.63 $Y=1.46 $X2=0
+ $Y2=0
cc_542 N_A_1034_392#_c_623_n N_A_1234_119#_M1030_g 0.0251416f $X=8.66 $Y=1.085
+ $X2=0 $Y2=0
cc_543 N_A_1034_392#_c_633_n N_A_1234_119#_M1030_g 0.0116969f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_544 N_A_1034_392#_c_621_n N_A_1234_119#_c_1207_n 9.01642e-19 $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_545 N_A_1034_392#_M1000_g N_A_1234_119#_c_1199_n 0.0110407f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_546 N_A_1034_392#_c_628_n N_A_1234_119#_c_1199_n 0.0110883f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_547 N_A_1034_392#_M1000_g N_A_1234_119#_c_1200_n 0.0071804f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_548 N_A_1034_392#_c_621_n N_A_1234_119#_c_1204_n 6.46907e-19 $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_549 N_A_1034_392#_M1000_g N_A_1234_119#_c_1204_n 0.00636651f $X=6.525
+ $Y=0.805 $X2=0 $Y2=0
cc_550 N_A_1034_392#_c_628_n N_A_1234_119#_c_1204_n 0.019863f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_551 N_A_1034_392#_c_657_p N_A_1234_119#_c_1204_n 0.00486547f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_552 N_A_1034_392#_c_642_n N_A_1234_119#_c_1212_n 2.99618e-19 $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_553 N_A_1034_392#_c_625_n N_A_1234_119#_c_1205_n 0.00319679f $X=8.735 $Y=1.16
+ $X2=0 $Y2=0
cc_554 N_A_1034_392#_c_646_n N_A_835_98#_c_1346_n 0.00258584f $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_555 N_A_1034_392#_c_647_n N_A_835_98#_c_1346_n 6.39872e-19 $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_556 N_A_1034_392#_c_626_n N_A_835_98#_c_1336_n 0.00991252f $X=5.36 $Y=0.78
+ $X2=0 $Y2=0
cc_557 N_A_1034_392#_c_627_n N_A_835_98#_c_1336_n 8.65367e-19 $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_558 N_A_1034_392#_c_637_n N_A_835_98#_c_1336_n 0.00191547f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_559 N_A_1034_392#_c_642_n N_A_835_98#_c_1347_n 0.0111007f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_560 N_A_1034_392#_c_643_n N_A_835_98#_c_1347_n 0.0130881f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_561 N_A_1034_392#_c_646_n N_A_835_98#_c_1347_n 4.97235e-19 $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_562 N_A_1034_392#_c_647_n N_A_835_98#_c_1347_n 0.0104193f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_563 N_A_1034_392#_c_643_n N_A_835_98#_c_1348_n 0.00899632f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_564 N_A_1034_392#_c_628_n N_A_835_98#_c_1337_n 0.00139627f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_565 N_A_1034_392#_c_630_n N_A_835_98#_c_1337_n 0.00441445f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_566 N_A_1034_392#_c_641_n N_A_835_98#_c_1337_n 0.0160947f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_567 N_A_1034_392#_M1000_g N_A_835_98#_c_1338_n 0.0223151f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_568 N_A_1034_392#_c_626_n N_A_835_98#_c_1338_n 0.00472785f $X=5.36 $Y=0.78
+ $X2=0 $Y2=0
cc_569 N_A_1034_392#_c_628_n N_A_835_98#_c_1338_n 0.00330666f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_570 N_A_1034_392#_c_643_n N_A_835_98#_M1010_g 0.0140799f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_571 N_A_1034_392#_c_621_n N_A_835_98#_M1010_g 0.00296839f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_572 N_A_1034_392#_c_645_n N_A_835_98#_c_1352_n 0.00464206f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_573 N_A_1034_392#_c_645_n N_A_835_98#_M1013_g 0.00689007f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_574 N_A_1034_392#_c_649_n N_A_835_98#_M1013_g 0.00157762f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_575 N_A_1034_392#_c_645_n N_A_835_98#_c_1339_n 0.0191375f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_576 N_A_1034_392#_c_636_n N_A_835_98#_c_1339_n 3.3013e-19 $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_577 N_A_1034_392#_c_649_n N_A_835_98#_c_1339_n 0.00813875f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_578 N_A_1034_392#_c_639_n N_A_835_98#_c_1339_n 0.0125871f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_579 N_A_1034_392#_c_640_n N_A_835_98#_c_1339_n 0.0175647f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_580 N_A_1034_392#_c_624_n N_A_835_98#_c_1340_n 0.0125871f $X=9.105 $Y=1.16
+ $X2=0 $Y2=0
cc_581 N_A_1034_392#_c_633_n N_A_835_98#_M1009_g 0.00370145f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_582 N_A_1034_392#_c_635_n N_A_835_98#_M1009_g 0.00158974f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_583 N_A_1034_392#_c_636_n N_A_835_98#_M1009_g 0.00266955f $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_584 N_A_1034_392#_c_639_n N_A_835_98#_M1009_g 0.0176907f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_585 N_A_1034_392#_c_640_n N_A_835_98#_M1009_g 0.00700032f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_586 N_A_1034_392#_c_627_n N_A_835_98#_c_1342_n 0.00563685f $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_587 N_A_1034_392#_c_646_n N_A_835_98#_c_1344_n 0.0199151f $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_588 N_A_1034_392#_c_627_n N_A_835_98#_c_1344_n 0.0236806f $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_589 N_A_1034_392#_c_647_n N_A_835_98#_c_1344_n 0.00665415f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_590 N_A_1034_392#_c_637_n N_A_835_98#_c_1344_n 0.00267749f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_591 N_A_1034_392#_c_646_n N_A_835_98#_c_1345_n 0.00634613f $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_592 N_A_1034_392#_c_627_n N_A_835_98#_c_1345_n 0.0141907f $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_593 N_A_1034_392#_c_628_n N_A_835_98#_c_1345_n 0.00385788f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_594 N_A_1034_392#_c_647_n N_A_835_98#_c_1345_n 0.0120306f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_595 N_A_1034_392#_c_630_n N_A_835_98#_c_1345_n 0.0116804f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_596 N_A_1034_392#_c_637_n N_A_835_98#_c_1345_n 0.0122529f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_597 N_A_1034_392#_c_641_n N_A_835_98#_c_1345_n 0.021574f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_598 N_A_1034_392#_c_640_n N_A_2008_48#_M1003_g 2.03511e-19 $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_599 N_A_1034_392#_c_645_n N_A_2008_48#_c_1516_n 0.0294704f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_600 N_A_1034_392#_c_649_n N_A_2008_48#_c_1516_n 0.0016211f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_601 N_A_1034_392#_c_645_n N_A_2008_48#_c_1524_n 0.0336986f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_602 N_A_1034_392#_c_633_n N_A_1747_74#_M1020_d 0.00174298f $X=8.825 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_603 N_A_1034_392#_c_635_n N_A_1747_74#_M1020_d 0.0115696f $X=8.91 $Y=0.905
+ $X2=-0.19 $Y2=-0.245
cc_604 N_A_1034_392#_c_638_n N_A_1747_74#_M1020_d 0.0018696f $X=9.27 $Y=1.07
+ $X2=-0.19 $Y2=-0.245
cc_605 N_A_1034_392#_c_645_n N_A_1747_74#_c_1678_n 0.00430249f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_606 N_A_1034_392#_c_649_n N_A_1747_74#_c_1678_n 0.0330459f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_607 N_A_1034_392#_c_640_n N_A_1747_74#_c_1678_n 0.0150349f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_608 N_A_1034_392#_c_623_n N_A_1747_74#_c_1681_n 6.51156e-19 $X=8.66 $Y=1.085
+ $X2=0 $Y2=0
cc_609 N_A_1034_392#_c_633_n N_A_1747_74#_c_1681_n 0.00169938f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_610 N_A_1034_392#_c_635_n N_A_1747_74#_c_1681_n 0.0248816f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_611 N_A_1034_392#_c_638_n N_A_1747_74#_c_1681_n 0.0199783f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_612 N_A_1034_392#_c_639_n N_A_1747_74#_c_1681_n 0.00615122f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_613 N_A_1034_392#_c_640_n N_A_1747_74#_c_1681_n 0.00536065f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_614 N_A_1034_392#_c_645_n N_A_1747_74#_c_1672_n 0.0159422f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_615 N_A_1034_392#_c_649_n N_A_1747_74#_c_1672_n 0.0169381f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_616 N_A_1034_392#_c_635_n N_A_1747_74#_c_1659_n 0.00508102f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_617 N_A_1034_392#_c_638_n N_A_1747_74#_c_1659_n 0.0078055f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_618 N_A_1034_392#_c_639_n N_A_1747_74#_c_1659_n 2.98286e-19 $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_619 N_A_1034_392#_c_645_n N_A_1747_74#_c_1660_n 0.00418565f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_620 N_A_1034_392#_c_649_n N_A_1747_74#_c_1660_n 0.0483469f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_621 N_A_1034_392#_c_640_n N_A_1747_74#_c_1660_n 0.0109876f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_622 N_A_1034_392#_c_636_n N_A_1747_74#_c_1661_n 0.015348f $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_623 N_A_1034_392#_c_638_n N_A_1747_74#_c_1661_n 0.00610378f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_624 N_A_1034_392#_c_639_n N_A_1747_74#_c_1661_n 0.00101813f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_625 N_A_1034_392#_c_640_n N_A_1747_74#_c_1661_n 0.0202102f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_626 N_A_1034_392#_c_645_n N_VPWR_c_1899_n 0.0038628f $X=9.77 $Y=2.37 $X2=0
+ $Y2=0
cc_627 N_A_1034_392#_c_643_n N_VPWR_c_1881_n 9.49986e-19 $X=6.135 $Y=2.21 $X2=0
+ $Y2=0
cc_628 N_A_1034_392#_c_645_n N_VPWR_c_1881_n 0.00515964f $X=9.77 $Y=2.37 $X2=0
+ $Y2=0
cc_629 N_A_1034_392#_M1028_d N_A_409_81#_c_2078_n 0.00695361f $X=5.17 $Y=1.96
+ $X2=0 $Y2=0
cc_630 N_A_1034_392#_c_646_n N_A_409_81#_c_2078_n 0.016647f $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_631 N_A_1034_392#_c_647_n N_A_409_81#_c_2078_n 0.0134529f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_632 N_A_1034_392#_c_630_n N_A_409_81#_c_2078_n 0.0029069f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_633 N_A_1034_392#_c_626_n N_A_409_81#_c_2069_n 0.0311322f $X=5.36 $Y=0.78
+ $X2=0 $Y2=0
cc_634 N_A_1034_392#_c_628_n N_A_409_81#_c_2069_n 0.013349f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_635 N_A_1034_392#_M1000_g N_A_409_81#_c_2070_n 3.66002e-19 $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_636 N_A_1034_392#_c_626_n N_A_409_81#_c_2070_n 0.00571418f $X=5.36 $Y=0.78
+ $X2=0 $Y2=0
cc_637 N_A_1034_392#_c_637_n N_A_409_81#_c_2070_n 0.00980399f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_638 N_A_1034_392#_c_643_n N_A_409_81#_c_2079_n 0.00783906f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_639 N_A_1034_392#_M1000_g N_A_409_81#_c_2071_n 0.00551398f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_640 N_A_1034_392#_c_630_n N_A_409_81#_c_2071_n 0.0142722f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_641 N_A_1034_392#_c_641_n N_A_409_81#_c_2071_n 0.00577594f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_642 N_A_1034_392#_c_630_n N_A_409_81#_c_2072_n 0.0145081f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_643 N_A_1034_392#_c_637_n N_A_409_81#_c_2072_n 0.013579f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_644 N_A_1034_392#_c_641_n N_A_409_81#_c_2072_n 3.38485e-19 $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_645 N_A_1034_392#_c_642_n N_A_409_81#_c_2080_n 0.00390532f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_646 N_A_1034_392#_c_643_n N_A_409_81#_c_2080_n 0.00843492f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_647 N_A_1034_392#_c_621_n N_A_409_81#_c_2080_n 0.00177679f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_648 N_A_1034_392#_c_630_n N_A_409_81#_c_2080_n 0.00615957f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_649 N_A_1034_392#_c_641_n N_A_409_81#_c_2080_n 6.46491e-19 $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_650 N_A_1034_392#_c_642_n N_A_409_81#_c_2081_n 0.00121768f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_651 N_A_1034_392#_c_643_n N_A_409_81#_c_2081_n 0.00154832f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_652 N_A_1034_392#_c_647_n N_A_409_81#_c_2081_n 0.0116706f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_653 N_A_1034_392#_c_630_n N_A_409_81#_c_2081_n 0.016874f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_654 N_A_1034_392#_c_641_n N_A_409_81#_c_2081_n 0.00278662f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_655 N_A_1034_392#_c_642_n N_A_409_81#_c_2073_n 0.00400586f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_656 N_A_1034_392#_c_621_n N_A_409_81#_c_2073_n 0.0122247f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_657 N_A_1034_392#_M1000_g N_A_409_81#_c_2073_n 0.00504469f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_658 N_A_1034_392#_c_630_n N_A_409_81#_c_2073_n 0.0250842f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_659 N_A_1034_392#_c_641_n N_A_409_81#_c_2073_n 0.00171299f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_660 N_A_1034_392#_c_632_n N_VGND_M1011_d 0.0170511f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_661 N_A_1034_392#_c_687_p N_VGND_M1011_d 0.00275919f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_662 N_A_1034_392#_c_634_n N_VGND_M1011_d 7.93589e-19 $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_663 N_A_1034_392#_c_626_n N_VGND_c_2285_n 0.0159443f $X=5.36 $Y=0.78 $X2=0
+ $Y2=0
cc_664 N_A_1034_392#_c_629_n N_VGND_c_2285_n 0.0144411f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_665 N_A_1034_392#_c_628_n N_VGND_c_2293_n 0.103356f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_666 N_A_1034_392#_c_629_n N_VGND_c_2293_n 0.0276098f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_667 N_A_1034_392#_c_632_n N_VGND_c_2293_n 0.00402072f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_668 N_A_1034_392#_c_623_n N_VGND_c_2294_n 0.00278271f $X=8.66 $Y=1.085 $X2=0
+ $Y2=0
cc_669 N_A_1034_392#_c_632_n N_VGND_c_2294_n 0.00335833f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_670 N_A_1034_392#_c_633_n N_VGND_c_2294_n 0.0579173f $X=8.825 $Y=0.34 $X2=0
+ $Y2=0
cc_671 N_A_1034_392#_c_634_n N_VGND_c_2294_n 0.0118998f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_672 N_A_1034_392#_c_623_n N_VGND_c_2297_n 0.00358617f $X=8.66 $Y=1.085 $X2=0
+ $Y2=0
cc_673 N_A_1034_392#_c_628_n N_VGND_c_2297_n 0.0538367f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_674 N_A_1034_392#_c_629_n N_VGND_c_2297_n 0.0138923f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_675 N_A_1034_392#_c_632_n N_VGND_c_2297_n 0.0122484f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_676 N_A_1034_392#_c_633_n N_VGND_c_2297_n 0.0324866f $X=8.825 $Y=0.34 $X2=0
+ $Y2=0
cc_677 N_A_1034_392#_c_634_n N_VGND_c_2297_n 0.00655543f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_678 N_A_1034_392#_c_628_n N_VGND_c_2300_n 0.0118008f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_679 N_A_1034_392#_c_632_n N_VGND_c_2300_n 0.0246154f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_680 N_A_1034_392#_c_634_n N_VGND_c_2300_n 0.0135793f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_681 N_A_1034_392#_c_657_p A_1397_119# 0.00349303f $X=7.22 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_682 N_A_1367_93#_M1021_g N_RESET_B_c_950_n 0.00882199f $X=6.91 $Y=0.805 $X2=0
+ $Y2=0
cc_683 N_A_1367_93#_c_841_n N_RESET_B_c_950_n 2.57602e-19 $X=7.265 $Y=1.005
+ $X2=0 $Y2=0
cc_684 N_A_1367_93#_M1021_g N_RESET_B_M1011_g 0.0398547f $X=6.91 $Y=0.805 $X2=0
+ $Y2=0
cc_685 N_A_1367_93#_c_839_n N_RESET_B_M1011_g 0.00116633f $X=7.145 $Y=1.64 $X2=0
+ $Y2=0
cc_686 N_A_1367_93#_c_841_n N_RESET_B_M1011_g 0.00250892f $X=7.265 $Y=1.005
+ $X2=0 $Y2=0
cc_687 N_A_1367_93#_c_845_n N_RESET_B_M1011_g 0.0104334f $X=8.27 $Y=0.842 $X2=0
+ $Y2=0
cc_688 N_A_1367_93#_M1021_g N_RESET_B_c_953_n 0.00178049f $X=6.91 $Y=0.805 $X2=0
+ $Y2=0
cc_689 N_A_1367_93#_c_839_n N_RESET_B_c_953_n 7.18471e-19 $X=7.145 $Y=1.64 $X2=0
+ $Y2=0
cc_690 N_A_1367_93#_c_840_n N_RESET_B_c_953_n 0.0209381f $X=7.145 $Y=1.64 $X2=0
+ $Y2=0
cc_691 N_A_1367_93#_c_839_n N_RESET_B_c_955_n 0.00822559f $X=7.145 $Y=1.64 $X2=0
+ $Y2=0
cc_692 N_A_1367_93#_c_840_n N_RESET_B_c_955_n 0.0059618f $X=7.145 $Y=1.64 $X2=0
+ $Y2=0
cc_693 N_A_1367_93#_c_845_n N_RESET_B_c_955_n 0.00903119f $X=8.27 $Y=0.842 $X2=0
+ $Y2=0
cc_694 N_A_1367_93#_M1034_g N_RESET_B_c_966_n 0.0065779f $X=6.945 $Y=2.495 $X2=0
+ $Y2=0
cc_695 N_A_1367_93#_c_839_n N_RESET_B_c_966_n 0.00621585f $X=7.145 $Y=1.64 $X2=0
+ $Y2=0
cc_696 N_A_1367_93#_c_840_n N_RESET_B_c_966_n 0.00171088f $X=7.145 $Y=1.64 $X2=0
+ $Y2=0
cc_697 N_A_1367_93#_M1040_d N_RESET_B_c_968_n 0.00328043f $X=8.62 $Y=1.735 $X2=0
+ $Y2=0
cc_698 N_A_1367_93#_c_843_n N_RESET_B_c_968_n 0.00640786f $X=8.81 $Y=1.415 $X2=0
+ $Y2=0
cc_699 N_A_1367_93#_c_844_n N_RESET_B_c_968_n 0.0247803f $X=8.77 $Y=1.88 $X2=0
+ $Y2=0
cc_700 N_A_1367_93#_M1034_g N_RESET_B_c_972_n 0.0207015f $X=6.945 $Y=2.495 $X2=0
+ $Y2=0
cc_701 N_A_1367_93#_c_842_n N_A_1234_119#_M1030_g 0.00325974f $X=8.57 $Y=1.245
+ $X2=0 $Y2=0
cc_702 N_A_1367_93#_c_845_n N_A_1234_119#_M1030_g 0.01076f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_703 N_A_1367_93#_c_846_n N_A_1234_119#_M1030_g 0.0114971f $X=8.57 $Y=0.842
+ $X2=0 $Y2=0
cc_704 N_A_1367_93#_c_844_n N_A_1234_119#_c_1206_n 0.00507431f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_705 N_A_1367_93#_M1034_g N_A_1234_119#_c_1207_n 0.00128347f $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_706 N_A_1367_93#_M1021_g N_A_1234_119#_c_1199_n 0.00419324f $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_707 N_A_1367_93#_c_841_n N_A_1234_119#_c_1199_n 0.00492865f $X=7.265 $Y=1.005
+ $X2=0 $Y2=0
cc_708 N_A_1367_93#_M1021_g N_A_1234_119#_c_1200_n 0.00722399f $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_709 N_A_1367_93#_M1034_g N_A_1234_119#_c_1200_n 0.00308621f $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_710 N_A_1367_93#_c_839_n N_A_1234_119#_c_1200_n 0.0512142f $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_711 N_A_1367_93#_c_840_n N_A_1234_119#_c_1200_n 0.00805995f $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_712 N_A_1367_93#_c_841_n N_A_1234_119#_c_1200_n 0.00480618f $X=7.265 $Y=1.005
+ $X2=0 $Y2=0
cc_713 N_A_1367_93#_M1034_g N_A_1234_119#_c_1209_n 0.00178971f $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_714 N_A_1367_93#_M1034_g N_A_1234_119#_c_1210_n 0.0175598f $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_715 N_A_1367_93#_c_839_n N_A_1234_119#_c_1210_n 0.0155534f $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_716 N_A_1367_93#_c_840_n N_A_1234_119#_c_1210_n 0.00383298f $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_717 N_A_1367_93#_M1034_g N_A_1234_119#_c_1201_n 0.00183154f $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_718 N_A_1367_93#_c_839_n N_A_1234_119#_c_1201_n 0.0190372f $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_719 N_A_1367_93#_c_840_n N_A_1234_119#_c_1201_n 0.00157419f $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_720 N_A_1367_93#_c_839_n N_A_1234_119#_c_1202_n 0.0243296f $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_721 N_A_1367_93#_c_840_n N_A_1234_119#_c_1202_n 4.90401e-19 $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_722 N_A_1367_93#_c_845_n N_A_1234_119#_c_1202_n 0.0135838f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_723 N_A_1367_93#_c_843_n N_A_1234_119#_c_1203_n 0.0132094f $X=8.81 $Y=1.415
+ $X2=0 $Y2=0
cc_724 N_A_1367_93#_c_844_n N_A_1234_119#_c_1203_n 0.00590456f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_725 N_A_1367_93#_c_845_n N_A_1234_119#_c_1203_n 0.0536947f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_726 N_A_1367_93#_M1021_g N_A_1234_119#_c_1204_n 0.00107025f $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_727 N_A_1367_93#_M1034_g N_A_1234_119#_c_1214_n 6.64763e-19 $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_728 N_A_1367_93#_c_843_n N_A_1234_119#_c_1205_n 0.00786811f $X=8.81 $Y=1.415
+ $X2=0 $Y2=0
cc_729 N_A_1367_93#_c_844_n N_A_1234_119#_c_1205_n 0.00580388f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_730 N_A_1367_93#_c_845_n N_A_1234_119#_c_1205_n 0.00365093f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_731 N_A_1367_93#_c_846_n N_A_1234_119#_c_1205_n 0.00401195f $X=8.57 $Y=0.842
+ $X2=0 $Y2=0
cc_732 N_A_1367_93#_M1034_g N_A_835_98#_M1010_g 0.0385033f $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_733 N_A_1367_93#_M1034_g N_A_835_98#_c_1351_n 0.00907339f $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_734 N_A_1367_93#_c_844_n N_A_835_98#_c_1351_n 0.00262042f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_735 N_A_1367_93#_c_844_n N_A_835_98#_c_1352_n 5.08057e-19 $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_736 N_A_1367_93#_c_844_n N_A_835_98#_M1013_g 0.0124176f $X=8.77 $Y=1.88 $X2=0
+ $Y2=0
cc_737 N_A_1367_93#_c_844_n N_A_835_98#_c_1340_n 0.00543498f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_738 N_A_1367_93#_c_844_n N_A_1747_74#_c_1678_n 0.0261048f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_739 N_A_1367_93#_c_844_n N_A_1747_74#_c_1673_n 0.0128087f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_740 N_A_1367_93#_M1034_g N_VPWR_c_1885_n 0.0033811f $X=6.945 $Y=2.495 $X2=0
+ $Y2=0
cc_741 N_A_1367_93#_c_844_n N_VPWR_c_1886_n 0.0670793f $X=8.77 $Y=1.88 $X2=0
+ $Y2=0
cc_742 N_A_1367_93#_c_846_n N_VPWR_c_1886_n 0.00607188f $X=8.57 $Y=0.842 $X2=0
+ $Y2=0
cc_743 N_A_1367_93#_c_844_n N_VPWR_c_1899_n 0.00567879f $X=8.77 $Y=1.88 $X2=0
+ $Y2=0
cc_744 N_A_1367_93#_M1034_g N_VPWR_c_1881_n 9.49986e-19 $X=6.945 $Y=2.495 $X2=0
+ $Y2=0
cc_745 N_A_1367_93#_c_844_n N_VPWR_c_1881_n 0.00684413f $X=8.77 $Y=1.88 $X2=0
+ $Y2=0
cc_746 N_A_1367_93#_M1034_g N_A_409_81#_c_2080_n 3.2345e-19 $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_747 N_A_1367_93#_M1021_g N_A_409_81#_c_2073_n 3.00253e-19 $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_748 N_A_1367_93#_M1034_g N_A_409_81#_c_2073_n 3.97102e-19 $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_749 N_A_1367_93#_c_840_n N_A_409_81#_c_2073_n 2.16488e-19 $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_750 N_A_1367_93#_c_845_n N_VGND_M1011_d 0.00911951f $X=8.27 $Y=0.842 $X2=0
+ $Y2=0
cc_751 N_A_1367_93#_c_841_n A_1397_119# 0.00138862f $X=7.265 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_752 N_RESET_B_c_955_n N_A_1234_119#_M1030_g 0.00443283f $X=7.595 $Y=1.19
+ $X2=0 $Y2=0
cc_753 N_RESET_B_c_968_n N_A_1234_119#_c_1206_n 0.00726918f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_754 N_RESET_B_c_966_n N_A_1234_119#_c_1207_n 0.00849024f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_755 N_RESET_B_M1011_g N_A_1234_119#_c_1199_n 3.7607e-19 $X=7.3 $Y=0.805 $X2=0
+ $Y2=0
cc_756 N_RESET_B_c_966_n N_A_1234_119#_c_1200_n 0.00946491f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_966_n N_A_1234_119#_c_1210_n 0.0312549f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_758 N_RESET_B_c_972_n N_A_1234_119#_c_1210_n 0.0100553f $X=7.595 $Y=2.002
+ $X2=0 $Y2=0
cc_759 N_RESET_B_c_953_n N_A_1234_119#_c_1201_n 0.0095642f $X=7.595 $Y=1.795
+ $X2=0 $Y2=0
cc_760 N_RESET_B_c_966_n N_A_1234_119#_c_1201_n 0.0099676f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_761 N_RESET_B_c_969_n N_A_1234_119#_c_1201_n 0.00109185f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_762 N_RESET_B_c_972_n N_A_1234_119#_c_1201_n 0.00515561f $X=7.595 $Y=2.002
+ $X2=0 $Y2=0
cc_763 N_RESET_B_c_973_n N_A_1234_119#_c_1201_n 0.0127277f $X=7.86 $Y=1.96 $X2=0
+ $Y2=0
cc_764 N_RESET_B_c_953_n N_A_1234_119#_c_1202_n 0.00374691f $X=7.595 $Y=1.795
+ $X2=0 $Y2=0
cc_765 N_RESET_B_c_955_n N_A_1234_119#_c_1202_n 0.00371515f $X=7.595 $Y=1.19
+ $X2=0 $Y2=0
cc_766 N_RESET_B_c_953_n N_A_1234_119#_c_1203_n 0.00661563f $X=7.595 $Y=1.795
+ $X2=0 $Y2=0
cc_767 N_RESET_B_c_955_n N_A_1234_119#_c_1203_n 5.9918e-19 $X=7.595 $Y=1.19
+ $X2=0 $Y2=0
cc_768 N_RESET_B_c_966_n N_A_1234_119#_c_1203_n 0.00552418f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_769 N_RESET_B_c_968_n N_A_1234_119#_c_1203_n 0.00610904f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_770 N_RESET_B_c_969_n N_A_1234_119#_c_1203_n 0.00265438f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_771 N_RESET_B_c_972_n N_A_1234_119#_c_1203_n 0.00540006f $X=7.595 $Y=2.002
+ $X2=0 $Y2=0
cc_772 N_RESET_B_c_973_n N_A_1234_119#_c_1203_n 0.0133891f $X=7.86 $Y=1.96 $X2=0
+ $Y2=0
cc_773 N_RESET_B_c_966_n N_A_1234_119#_c_1212_n 0.0126021f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_774 N_RESET_B_c_966_n N_A_1234_119#_c_1281_n 0.0125017f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_775 N_RESET_B_c_969_n N_A_1234_119#_c_1281_n 0.00115111f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_776 N_RESET_B_c_972_n N_A_1234_119#_c_1281_n 0.00650869f $X=7.595 $Y=2.002
+ $X2=0 $Y2=0
cc_777 N_RESET_B_c_973_n N_A_1234_119#_c_1281_n 0.0109284f $X=7.86 $Y=1.96 $X2=0
+ $Y2=0
cc_778 N_RESET_B_c_961_n N_A_1234_119#_c_1213_n 0.00633065f $X=7.395 $Y=2.21
+ $X2=0 $Y2=0
cc_779 N_RESET_B_c_966_n N_A_1234_119#_c_1213_n 0.00702421f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_780 N_RESET_B_c_972_n N_A_1234_119#_c_1213_n 0.00724773f $X=7.595 $Y=2.002
+ $X2=0 $Y2=0
cc_781 N_RESET_B_c_961_n N_A_1234_119#_c_1214_n 0.00390298f $X=7.395 $Y=2.21
+ $X2=0 $Y2=0
cc_782 N_RESET_B_c_972_n N_A_1234_119#_c_1214_n 0.00528559f $X=7.595 $Y=2.002
+ $X2=0 $Y2=0
cc_783 N_RESET_B_c_953_n N_A_1234_119#_c_1205_n 5.38903e-19 $X=7.595 $Y=1.795
+ $X2=0 $Y2=0
cc_784 N_RESET_B_c_955_n N_A_1234_119#_c_1205_n 0.0132285f $X=7.595 $Y=1.19
+ $X2=0 $Y2=0
cc_785 N_RESET_B_c_968_n N_A_1234_119#_c_1205_n 0.00423661f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_786 N_RESET_B_c_969_n N_A_1234_119#_c_1205_n 7.23568e-19 $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_787 N_RESET_B_c_972_n N_A_1234_119#_c_1205_n 0.0023769f $X=7.595 $Y=2.002
+ $X2=0 $Y2=0
cc_788 N_RESET_B_c_973_n N_A_1234_119#_c_1205_n 3.48298e-19 $X=7.86 $Y=1.96
+ $X2=0 $Y2=0
cc_789 N_RESET_B_c_966_n N_A_835_98#_M1024_s 0.00114217f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_790 N_RESET_B_c_966_n N_A_835_98#_c_1346_n 0.00350083f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_791 N_RESET_B_c_950_n N_A_835_98#_c_1336_n 0.0103973f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_792 N_RESET_B_c_966_n N_A_835_98#_c_1347_n 0.00218847f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_793 N_RESET_B_c_950_n N_A_835_98#_c_1338_n 0.00882199f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_794 N_RESET_B_c_966_n N_A_835_98#_M1010_g 0.00325607f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_795 N_RESET_B_c_961_n N_A_835_98#_c_1351_n 0.00889176f $X=7.395 $Y=2.21 $X2=0
+ $Y2=0
cc_796 N_RESET_B_c_968_n N_A_835_98#_M1013_g 0.0105606f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_797 N_RESET_B_c_968_n N_A_835_98#_c_1339_n 0.00463969f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_798 N_RESET_B_c_950_n N_A_835_98#_c_1363_n 0.00146684f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_799 N_RESET_B_M1036_g N_A_835_98#_c_1343_n 0.00389848f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_800 N_RESET_B_c_950_n N_A_835_98#_c_1343_n 0.00806854f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_801 N_RESET_B_c_959_n N_A_835_98#_c_1344_n 0.0011403f $X=3.93 $Y=1.995 $X2=0
+ $Y2=0
cc_802 N_RESET_B_c_960_n N_A_835_98#_c_1344_n 0.00130059f $X=3.695 $Y=1.995
+ $X2=0 $Y2=0
cc_803 N_RESET_B_c_966_n N_A_835_98#_c_1344_n 0.0468629f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_804 N_RESET_B_c_967_n N_A_835_98#_c_1344_n 0.00284227f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_805 N_RESET_B_c_971_n N_A_835_98#_c_1344_n 0.0281559f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_806 N_RESET_B_c_966_n N_A_835_98#_c_1345_n 0.00151487f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_807 N_RESET_B_M1005_g N_A_2008_48#_M1003_g 0.0358144f $X=10.545 $Y=0.58 $X2=0
+ $Y2=0
cc_808 N_RESET_B_c_957_n N_A_2008_48#_M1003_g 0.00188557f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_809 N_RESET_B_c_956_n N_A_2008_48#_c_1516_n 0.0030428f $X=10.81 $Y=1.335
+ $X2=0 $Y2=0
cc_810 N_RESET_B_c_968_n N_A_2008_48#_c_1516_n 0.00247648f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_811 RESET_B N_A_2008_48#_c_1516_n 7.14482e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_812 N_RESET_B_c_975_n N_A_2008_48#_c_1516_n 0.00169359f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_813 N_RESET_B_c_957_n N_A_2008_48#_c_1516_n 0.0249721f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_814 N_RESET_B_c_964_n N_A_2008_48#_c_1523_n 0.00373821f $X=10.81 $Y=2.22
+ $X2=0 $Y2=0
cc_815 N_RESET_B_c_965_n N_A_2008_48#_c_1523_n 0.00276573f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_816 N_RESET_B_c_968_n N_A_2008_48#_c_1523_n 0.00755701f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_817 N_RESET_B_c_974_n N_A_2008_48#_c_1523_n 6.88508e-19 $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_818 N_RESET_B_c_965_n N_A_2008_48#_c_1524_n 0.0107901f $X=10.81 $Y=2.37 $X2=0
+ $Y2=0
cc_819 N_RESET_B_c_964_n N_A_2008_48#_c_1517_n 0.00199769f $X=10.81 $Y=2.22
+ $X2=0 $Y2=0
cc_820 N_RESET_B_c_965_n N_A_2008_48#_c_1517_n 0.00241136f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_821 N_RESET_B_c_968_n N_A_2008_48#_c_1517_n 0.0174665f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_822 RESET_B N_A_2008_48#_c_1517_n 0.00269473f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_823 N_RESET_B_c_974_n N_A_2008_48#_c_1517_n 4.38169e-19 $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_824 N_RESET_B_c_975_n N_A_2008_48#_c_1517_n 0.0344591f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_825 N_RESET_B_c_957_n N_A_2008_48#_c_1517_n 2.34208e-19 $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_826 N_RESET_B_c_965_n N_A_2008_48#_c_1526_n 0.00976826f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_827 N_RESET_B_c_968_n N_A_2008_48#_c_1526_n 0.00560031f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_828 RESET_B N_A_2008_48#_c_1526_n 0.00309934f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_829 N_RESET_B_c_975_n N_A_2008_48#_c_1526_n 0.00989058f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_830 N_RESET_B_c_965_n N_A_2008_48#_c_1528_n 0.00646344f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_831 N_RESET_B_c_964_n N_A_2008_48#_c_1529_n 0.0015825f $X=10.81 $Y=2.22 $X2=0
+ $Y2=0
cc_832 N_RESET_B_c_965_n N_A_2008_48#_c_1529_n 5.62382e-19 $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_833 RESET_B N_A_2008_48#_c_1529_n 0.00125949f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_834 N_RESET_B_c_974_n N_A_2008_48#_c_1529_n 0.00110518f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_835 N_RESET_B_c_975_n N_A_2008_48#_c_1529_n 0.0258608f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_836 N_RESET_B_c_974_n N_A_2008_48#_c_1519_n 8.24141e-19 $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_837 N_RESET_B_c_975_n N_A_2008_48#_c_1519_n 0.00968802f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_838 N_RESET_B_c_957_n N_A_2008_48#_c_1519_n 0.00111902f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_839 N_RESET_B_c_965_n N_A_2008_48#_c_1532_n 0.00389165f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_840 RESET_B N_A_2008_48#_c_1532_n 7.29139e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_841 N_RESET_B_c_974_n N_A_2008_48#_c_1532_n 8.21335e-19 $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_842 N_RESET_B_c_975_n N_A_2008_48#_c_1532_n 0.0169044f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_843 N_RESET_B_M1005_g N_A_2008_48#_c_1521_n 0.00108873f $X=10.545 $Y=0.58
+ $X2=0 $Y2=0
cc_844 N_RESET_B_c_968_n N_A_1747_74#_M1013_d 0.00220193f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_845 N_RESET_B_M1005_g N_A_1747_74#_c_1651_n 0.0481778f $X=10.545 $Y=0.58
+ $X2=0 $Y2=0
cc_846 N_RESET_B_c_956_n N_A_1747_74#_c_1652_n 0.00304958f $X=10.81 $Y=1.335
+ $X2=0 $Y2=0
cc_847 N_RESET_B_c_974_n N_A_1747_74#_c_1652_n 0.00202705f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_848 N_RESET_B_M1005_g N_A_1747_74#_c_1653_n 0.00503338f $X=10.545 $Y=0.58
+ $X2=0 $Y2=0
cc_849 N_RESET_B_c_965_n N_A_1747_74#_c_1663_n 0.00937718f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_850 N_RESET_B_c_964_n N_A_1747_74#_c_1664_n 0.00655145f $X=10.81 $Y=2.22
+ $X2=0 $Y2=0
cc_851 N_RESET_B_c_975_n N_A_1747_74#_c_1664_n 8.64724e-19 $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_852 N_RESET_B_c_956_n N_A_1747_74#_c_1656_n 0.0113835f $X=10.81 $Y=1.335
+ $X2=0 $Y2=0
cc_853 N_RESET_B_c_974_n N_A_1747_74#_c_1656_n 0.0205072f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_854 N_RESET_B_c_957_n N_A_1747_74#_c_1656_n 0.00965718f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_855 N_RESET_B_c_965_n N_A_1747_74#_c_1670_n 0.00814266f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_856 N_RESET_B_c_968_n N_A_1747_74#_c_1678_n 0.0211312f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_857 N_RESET_B_c_965_n N_A_1747_74#_c_1672_n 7.86001e-19 $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_858 N_RESET_B_c_968_n N_A_1747_74#_c_1672_n 0.0154438f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_859 N_RESET_B_c_968_n N_A_1747_74#_c_1660_n 0.0224891f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_860 N_RESET_B_c_957_n N_A_1747_74#_c_1660_n 9.47605e-19 $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_861 N_RESET_B_M1005_g N_A_1747_74#_c_1662_n 0.0173454f $X=10.545 $Y=0.58
+ $X2=0 $Y2=0
cc_862 N_RESET_B_c_956_n N_A_1747_74#_c_1662_n 0.0168092f $X=10.81 $Y=1.335
+ $X2=0 $Y2=0
cc_863 N_RESET_B_c_968_n N_A_1747_74#_c_1662_n 0.0108974f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_864 RESET_B N_A_1747_74#_c_1662_n 0.00277891f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_865 N_RESET_B_c_974_n N_A_1747_74#_c_1662_n 0.00194273f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_866 N_RESET_B_c_975_n N_A_1747_74#_c_1662_n 0.0211796f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_867 N_RESET_B_c_957_n N_A_1747_74#_c_1662_n 0.00355179f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_868 N_RESET_B_c_966_n N_VPWR_M1024_d 5.797e-19 $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_869 N_RESET_B_c_968_n N_VPWR_M1040_s 0.00248619f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_870 N_RESET_B_c_963_n N_VPWR_c_1883_n 0.00529153f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_871 N_RESET_B_c_961_n N_VPWR_c_1885_n 0.00279283f $X=7.395 $Y=2.21 $X2=0
+ $Y2=0
cc_872 N_RESET_B_c_966_n N_VPWR_c_1885_n 0.00177009f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_873 N_RESET_B_c_953_n N_VPWR_c_1886_n 0.00118732f $X=7.595 $Y=1.795 $X2=0
+ $Y2=0
cc_874 N_RESET_B_c_968_n N_VPWR_c_1886_n 0.0257367f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_875 N_RESET_B_c_969_n N_VPWR_c_1886_n 0.00264233f $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_876 N_RESET_B_c_972_n N_VPWR_c_1886_n 0.00234646f $X=7.595 $Y=2.002 $X2=0
+ $Y2=0
cc_877 N_RESET_B_c_973_n N_VPWR_c_1886_n 0.0221742f $X=7.86 $Y=1.96 $X2=0 $Y2=0
cc_878 N_RESET_B_c_965_n N_VPWR_c_1887_n 0.00552432f $X=10.81 $Y=2.37 $X2=0
+ $Y2=0
cc_879 N_RESET_B_c_968_n N_VPWR_c_1887_n 0.00114209f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_880 N_RESET_B_c_963_n N_VPWR_c_1892_n 0.00445602f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_881 N_RESET_B_c_965_n N_VPWR_c_1900_n 0.00497687f $X=10.81 $Y=2.37 $X2=0
+ $Y2=0
cc_882 N_RESET_B_c_961_n N_VPWR_c_1881_n 9.49986e-19 $X=7.395 $Y=2.21 $X2=0
+ $Y2=0
cc_883 N_RESET_B_c_963_n N_VPWR_c_1881_n 0.00443364f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_884 N_RESET_B_c_965_n N_VPWR_c_1881_n 0.00515964f $X=10.81 $Y=2.37 $X2=0
+ $Y2=0
cc_885 N_RESET_B_M1036_g N_A_409_81#_c_2067_n 0.0137342f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_886 N_RESET_B_c_960_n N_A_409_81#_c_2107_n 8.35086e-19 $X=3.695 $Y=1.995
+ $X2=0 $Y2=0
cc_887 N_RESET_B_M1036_g N_A_409_81#_c_2068_n 0.018686f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_888 N_RESET_B_c_960_n N_A_409_81#_c_2068_n 0.0188904f $X=3.695 $Y=1.995 $X2=0
+ $Y2=0
cc_889 N_RESET_B_c_963_n N_A_409_81#_c_2068_n 0.00445911f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_890 N_RESET_B_c_967_n N_A_409_81#_c_2068_n 0.00108729f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_891 N_RESET_B_c_971_n N_A_409_81#_c_2068_n 0.0243953f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_892 N_RESET_B_c_966_n N_A_409_81#_c_2076_n 0.00515092f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_893 N_RESET_B_c_959_n N_A_409_81#_c_2077_n 0.00525707f $X=3.93 $Y=1.995 $X2=0
+ $Y2=0
cc_894 N_RESET_B_c_963_n N_A_409_81#_c_2077_n 0.0137138f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_895 N_RESET_B_c_966_n N_A_409_81#_c_2077_n 0.00101627f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_896 N_RESET_B_c_967_n N_A_409_81#_c_2077_n 0.00440623f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_897 N_RESET_B_c_971_n N_A_409_81#_c_2077_n 0.0258218f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_898 N_RESET_B_c_966_n N_A_409_81#_c_2078_n 0.0137461f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_899 N_RESET_B_c_966_n N_A_409_81#_c_2071_n 0.00348472f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_900 N_RESET_B_c_966_n N_A_409_81#_c_2080_n 0.0172886f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_901 N_RESET_B_c_966_n N_A_409_81#_c_2081_n 0.0167671f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_902 N_RESET_B_c_966_n N_A_409_81#_c_2073_n 0.00940891f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_903 N_RESET_B_c_963_n N_A_409_81#_c_2084_n 0.00549198f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_904 N_RESET_B_M1036_g N_VGND_c_2284_n 0.00141396f $X=3.5 $Y=0.615 $X2=0 $Y2=0
cc_905 N_RESET_B_c_950_n N_VGND_c_2284_n 0.0208132f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_906 N_RESET_B_c_950_n N_VGND_c_2285_n 0.0253641f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_907 N_RESET_B_M1005_g N_VGND_c_2286_n 0.0110663f $X=10.545 $Y=0.58 $X2=0
+ $Y2=0
cc_908 N_RESET_B_c_950_n N_VGND_c_2289_n 0.0242408f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_909 N_RESET_B_c_951_n N_VGND_c_2292_n 0.0064002f $X=3.575 $Y=0.18 $X2=0 $Y2=0
cc_910 N_RESET_B_c_950_n N_VGND_c_2293_n 0.0512939f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_911 N_RESET_B_M1005_g N_VGND_c_2295_n 0.00383152f $X=10.545 $Y=0.58 $X2=0
+ $Y2=0
cc_912 N_RESET_B_c_950_n N_VGND_c_2297_n 0.0887542f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_913 N_RESET_B_c_951_n N_VGND_c_2297_n 0.0113744f $X=3.575 $Y=0.18 $X2=0 $Y2=0
cc_914 N_RESET_B_M1005_g N_VGND_c_2297_n 0.0075694f $X=10.545 $Y=0.58 $X2=0
+ $Y2=0
cc_915 N_RESET_B_c_950_n N_VGND_c_2300_n 0.00939536f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_916 N_RESET_B_M1036_g N_noxref_25_c_2424_n 0.00190559f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_917 N_A_1234_119#_c_1207_n N_A_835_98#_c_1348_n 0.00321336f $X=6.685 $Y=2.555
+ $X2=0 $Y2=0
cc_918 N_A_1234_119#_c_1204_n N_A_835_98#_c_1338_n 0.00566398f $X=6.31 $Y=0.81
+ $X2=0 $Y2=0
cc_919 N_A_1234_119#_c_1207_n N_A_835_98#_M1010_g 0.0121868f $X=6.685 $Y=2.555
+ $X2=0 $Y2=0
cc_920 N_A_1234_119#_c_1209_n N_A_835_98#_M1010_g 0.00150864f $X=6.77 $Y=2.385
+ $X2=0 $Y2=0
cc_921 N_A_1234_119#_c_1206_n N_A_835_98#_c_1351_n 0.0103562f $X=8.545 $Y=1.66
+ $X2=0 $Y2=0
cc_922 N_A_1234_119#_c_1207_n N_A_835_98#_c_1351_n 0.00208418f $X=6.685 $Y=2.555
+ $X2=0 $Y2=0
cc_923 N_A_1234_119#_c_1213_n N_A_835_98#_c_1351_n 0.00592408f $X=7.62 $Y=2.53
+ $X2=0 $Y2=0
cc_924 N_A_1234_119#_c_1206_n N_A_835_98#_c_1352_n 0.00249951f $X=8.545 $Y=1.66
+ $X2=0 $Y2=0
cc_925 N_A_1234_119#_c_1206_n N_A_835_98#_M1013_g 0.00575058f $X=8.545 $Y=1.66
+ $X2=0 $Y2=0
cc_926 N_A_1234_119#_c_1205_n N_A_835_98#_c_1340_n 0.00675058f $X=8.22 $Y=1.452
+ $X2=0 $Y2=0
cc_927 N_A_1234_119#_c_1207_n N_VPWR_c_1885_n 0.00162755f $X=6.685 $Y=2.555
+ $X2=0 $Y2=0
cc_928 N_A_1234_119#_c_1210_n N_VPWR_c_1885_n 0.0152964f $X=7.435 $Y=2.075 $X2=0
+ $Y2=0
cc_929 N_A_1234_119#_c_1213_n N_VPWR_c_1885_n 0.0165552f $X=7.62 $Y=2.53 $X2=0
+ $Y2=0
cc_930 N_A_1234_119#_c_1206_n N_VPWR_c_1886_n 0.0152342f $X=8.545 $Y=1.66 $X2=0
+ $Y2=0
cc_931 N_A_1234_119#_c_1201_n N_VPWR_c_1886_n 0.00208581f $X=7.52 $Y=1.985 $X2=0
+ $Y2=0
cc_932 N_A_1234_119#_c_1203_n N_VPWR_c_1886_n 0.00632637f $X=8.15 $Y=1.41 $X2=0
+ $Y2=0
cc_933 N_A_1234_119#_c_1281_n N_VPWR_c_1886_n 4.28343e-19 $X=7.52 $Y=2.075 $X2=0
+ $Y2=0
cc_934 N_A_1234_119#_c_1213_n N_VPWR_c_1886_n 0.0158369f $X=7.62 $Y=2.53 $X2=0
+ $Y2=0
cc_935 N_A_1234_119#_c_1214_n N_VPWR_c_1886_n 0.00433112f $X=7.6 $Y=2.32 $X2=0
+ $Y2=0
cc_936 N_A_1234_119#_c_1205_n N_VPWR_c_1886_n 0.00664035f $X=8.22 $Y=1.452 $X2=0
+ $Y2=0
cc_937 N_A_1234_119#_c_1207_n N_VPWR_c_1894_n 0.0122106f $X=6.685 $Y=2.555 $X2=0
+ $Y2=0
cc_938 N_A_1234_119#_c_1213_n N_VPWR_c_1898_n 0.00718093f $X=7.62 $Y=2.53 $X2=0
+ $Y2=0
cc_939 N_A_1234_119#_c_1206_n N_VPWR_c_1881_n 8.51577e-19 $X=8.545 $Y=1.66 $X2=0
+ $Y2=0
cc_940 N_A_1234_119#_c_1207_n N_VPWR_c_1881_n 0.0157408f $X=6.685 $Y=2.555 $X2=0
+ $Y2=0
cc_941 N_A_1234_119#_c_1213_n N_VPWR_c_1881_n 0.00888445f $X=7.62 $Y=2.53 $X2=0
+ $Y2=0
cc_942 N_A_1234_119#_c_1204_n N_A_409_81#_c_2070_n 0.0168132f $X=6.31 $Y=0.81
+ $X2=0 $Y2=0
cc_943 N_A_1234_119#_c_1207_n N_A_409_81#_c_2079_n 0.0139433f $X=6.685 $Y=2.555
+ $X2=0 $Y2=0
cc_944 N_A_1234_119#_c_1209_n N_A_409_81#_c_2079_n 0.00314452f $X=6.77 $Y=2.385
+ $X2=0 $Y2=0
cc_945 N_A_1234_119#_c_1199_n N_A_409_81#_c_2071_n 0.00342789f $X=6.685 $Y=0.945
+ $X2=0 $Y2=0
cc_946 N_A_1234_119#_c_1200_n N_A_409_81#_c_2071_n 0.0136392f $X=6.77 $Y=1.985
+ $X2=0 $Y2=0
cc_947 N_A_1234_119#_c_1204_n N_A_409_81#_c_2071_n 0.0270482f $X=6.31 $Y=0.81
+ $X2=0 $Y2=0
cc_948 N_A_1234_119#_c_1207_n N_A_409_81#_c_2080_n 0.0180051f $X=6.685 $Y=2.555
+ $X2=0 $Y2=0
cc_949 N_A_1234_119#_c_1209_n N_A_409_81#_c_2080_n 0.00396213f $X=6.77 $Y=2.385
+ $X2=0 $Y2=0
cc_950 N_A_1234_119#_c_1212_n N_A_409_81#_c_2080_n 0.0100574f $X=6.77 $Y=2.075
+ $X2=0 $Y2=0
cc_951 N_A_1234_119#_c_1200_n N_A_409_81#_c_2073_n 0.0447672f $X=6.77 $Y=1.985
+ $X2=0 $Y2=0
cc_952 N_A_1234_119#_c_1212_n N_A_409_81#_c_2073_n 0.00431721f $X=6.77 $Y=2.075
+ $X2=0 $Y2=0
cc_953 N_A_1234_119#_M1030_g N_VGND_c_2294_n 0.00278271f $X=8.22 $Y=0.69 $X2=0
+ $Y2=0
cc_954 N_A_1234_119#_M1030_g N_VGND_c_2297_n 0.00358617f $X=8.22 $Y=0.69 $X2=0
+ $Y2=0
cc_955 N_A_1234_119#_M1030_g N_VGND_c_2300_n 0.00111149f $X=8.22 $Y=0.69 $X2=0
+ $Y2=0
cc_956 N_A_1234_119#_c_1199_n A_1320_119# 0.00179335f $X=6.685 $Y=0.945
+ $X2=-0.19 $Y2=-0.245
cc_957 N_A_835_98#_M1009_g N_A_2008_48#_M1003_g 0.0422064f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_958 N_A_835_98#_c_1339_n N_A_2008_48#_c_1516_n 0.0427595f $X=9.68 $Y=1.585
+ $X2=0 $Y2=0
cc_959 N_A_835_98#_M1013_g N_A_1747_74#_c_1678_n 2.44304e-19 $X=8.995 $Y=2.235
+ $X2=0 $Y2=0
cc_960 N_A_835_98#_c_1339_n N_A_1747_74#_c_1678_n 0.00473791f $X=9.68 $Y=1.585
+ $X2=0 $Y2=0
cc_961 N_A_835_98#_M1009_g N_A_1747_74#_c_1681_n 0.0150096f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_962 N_A_835_98#_M1013_g N_A_1747_74#_c_1673_n 0.00211239f $X=8.995 $Y=2.235
+ $X2=0 $Y2=0
cc_963 N_A_835_98#_M1009_g N_A_1747_74#_c_1659_n 0.00884302f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_964 N_A_835_98#_M1009_g N_A_1747_74#_c_1660_n 0.0014557f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_965 N_A_835_98#_c_1339_n N_A_1747_74#_c_1661_n 4.03784e-19 $X=9.68 $Y=1.585
+ $X2=0 $Y2=0
cc_966 N_A_835_98#_M1009_g N_A_1747_74#_c_1661_n 0.0141061f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_967 N_A_835_98#_c_1344_n N_VPWR_M1024_d 0.00264465f $X=4.93 $Y=1.852 $X2=0
+ $Y2=0
cc_968 N_A_835_98#_c_1346_n N_VPWR_c_1884_n 0.00850453f $X=5.095 $Y=1.875 $X2=0
+ $Y2=0
cc_969 N_A_835_98#_c_1347_n N_VPWR_c_1884_n 0.00158412f $X=5.615 $Y=3.075 $X2=0
+ $Y2=0
cc_970 N_A_835_98#_c_1349_n N_VPWR_c_1884_n 0.00232909f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_971 N_A_835_98#_M1010_g N_VPWR_c_1885_n 0.00714317f $X=6.585 $Y=2.495 $X2=0
+ $Y2=0
cc_972 N_A_835_98#_c_1351_n N_VPWR_c_1885_n 0.0210626f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_973 N_A_835_98#_c_1351_n N_VPWR_c_1886_n 0.0213056f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_974 N_A_835_98#_c_1352_n N_VPWR_c_1886_n 0.00613773f $X=8.995 $Y=2.9 $X2=0
+ $Y2=0
cc_975 N_A_835_98#_M1013_g N_VPWR_c_1886_n 6.49178e-19 $X=8.995 $Y=2.235 $X2=0
+ $Y2=0
cc_976 N_A_835_98#_c_1346_n N_VPWR_c_1894_n 0.00303678f $X=5.095 $Y=1.875 $X2=0
+ $Y2=0
cc_977 N_A_835_98#_c_1349_n N_VPWR_c_1894_n 0.0423252f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_978 N_A_835_98#_c_1351_n N_VPWR_c_1898_n 0.0305306f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_979 N_A_835_98#_c_1351_n N_VPWR_c_1899_n 0.0193014f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_980 N_A_835_98#_c_1346_n N_VPWR_c_1881_n 0.00394737f $X=5.095 $Y=1.875 $X2=0
+ $Y2=0
cc_981 N_A_835_98#_c_1348_n N_VPWR_c_1881_n 0.0241704f $X=6.51 $Y=3.15 $X2=0
+ $Y2=0
cc_982 N_A_835_98#_c_1349_n N_VPWR_c_1881_n 0.00688721f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_983 N_A_835_98#_c_1351_n N_VPWR_c_1881_n 0.077582f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_984 N_A_835_98#_c_1357_n N_VPWR_c_1881_n 0.00423956f $X=6.585 $Y=3.15 $X2=0
+ $Y2=0
cc_985 N_A_835_98#_M1024_s N_A_409_81#_c_2076_n 0.00851724f $X=4.275 $Y=1.96
+ $X2=0 $Y2=0
cc_986 N_A_835_98#_c_1344_n N_A_409_81#_c_2076_n 0.0175531f $X=4.93 $Y=1.852
+ $X2=0 $Y2=0
cc_987 N_A_835_98#_c_1346_n N_A_409_81#_c_2078_n 0.0151931f $X=5.095 $Y=1.875
+ $X2=0 $Y2=0
cc_988 N_A_835_98#_c_1347_n N_A_409_81#_c_2078_n 0.0148953f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_989 N_A_835_98#_c_1348_n N_A_409_81#_c_2078_n 7.24606e-19 $X=6.51 $Y=3.15
+ $X2=0 $Y2=0
cc_990 N_A_835_98#_c_1344_n N_A_409_81#_c_2078_n 0.0189697f $X=4.93 $Y=1.852
+ $X2=0 $Y2=0
cc_991 N_A_835_98#_c_1345_n N_A_409_81#_c_2078_n 4.98991e-19 $X=5.115 $Y=1.635
+ $X2=0 $Y2=0
cc_992 N_A_835_98#_c_1337_n N_A_409_81#_c_2070_n 0.00777044f $X=6.02 $Y=1.225
+ $X2=0 $Y2=0
cc_993 N_A_835_98#_c_1338_n N_A_409_81#_c_2070_n 0.00423903f $X=6.095 $Y=1.115
+ $X2=0 $Y2=0
cc_994 N_A_835_98#_c_1347_n N_A_409_81#_c_2079_n 0.00760865f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_995 N_A_835_98#_c_1348_n N_A_409_81#_c_2079_n 0.00469098f $X=6.51 $Y=3.15
+ $X2=0 $Y2=0
cc_996 N_A_835_98#_M1010_g N_A_409_81#_c_2079_n 5.52147e-19 $X=6.585 $Y=2.495
+ $X2=0 $Y2=0
cc_997 N_A_835_98#_c_1337_n N_A_409_81#_c_2071_n 0.0119917f $X=6.02 $Y=1.225
+ $X2=0 $Y2=0
cc_998 N_A_835_98#_c_1337_n N_A_409_81#_c_2072_n 0.00600188f $X=6.02 $Y=1.225
+ $X2=0 $Y2=0
cc_999 N_A_835_98#_c_1345_n N_A_409_81#_c_2072_n 7.71188e-19 $X=5.115 $Y=1.635
+ $X2=0 $Y2=0
cc_1000 N_A_835_98#_M1010_g N_A_409_81#_c_2080_n 0.00138335f $X=6.585 $Y=2.495
+ $X2=0 $Y2=0
cc_1001 N_A_835_98#_c_1347_n N_A_409_81#_c_2081_n 0.00126f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_1002 N_A_835_98#_c_1345_n N_A_409_81#_c_2073_n 0.00436361f $X=5.115 $Y=1.635
+ $X2=0 $Y2=0
cc_1003 N_A_835_98#_c_1363_n N_VGND_M1025_d 0.00765303f $X=4.815 $Y=0.925 $X2=0
+ $Y2=0
cc_1004 N_A_835_98#_c_1342_n N_VGND_M1025_d 0.00533363f $X=4.93 $Y=1.455 $X2=0
+ $Y2=0
cc_1005 N_A_835_98#_c_1343_n N_VGND_c_2284_n 0.0158255f $X=4.32 $Y=0.665 $X2=0
+ $Y2=0
cc_1006 N_A_835_98#_c_1336_n N_VGND_c_2285_n 0.00167937f $X=5.145 $Y=1.41 $X2=0
+ $Y2=0
cc_1007 N_A_835_98#_c_1363_n N_VGND_c_2285_n 0.0243898f $X=4.815 $Y=0.925 $X2=0
+ $Y2=0
cc_1008 N_A_835_98#_c_1343_n N_VGND_c_2285_n 0.0105328f $X=4.32 $Y=0.665 $X2=0
+ $Y2=0
cc_1009 N_A_835_98#_M1009_g N_VGND_c_2286_n 0.00177088f $X=9.755 $Y=0.58 $X2=0
+ $Y2=0
cc_1010 N_A_835_98#_c_1343_n N_VGND_c_2289_n 0.0104074f $X=4.32 $Y=0.665 $X2=0
+ $Y2=0
cc_1011 N_A_835_98#_M1009_g N_VGND_c_2294_n 0.00358451f $X=9.755 $Y=0.58 $X2=0
+ $Y2=0
cc_1012 N_A_835_98#_c_1336_n N_VGND_c_2297_n 9.10391e-19 $X=5.145 $Y=1.41 $X2=0
+ $Y2=0
cc_1013 N_A_835_98#_M1009_g N_VGND_c_2297_n 0.00569641f $X=9.755 $Y=0.58 $X2=0
+ $Y2=0
cc_1014 N_A_835_98#_c_1363_n N_VGND_c_2297_n 0.00633041f $X=4.815 $Y=0.925 $X2=0
+ $Y2=0
cc_1015 N_A_835_98#_c_1343_n N_VGND_c_2297_n 0.0115264f $X=4.32 $Y=0.665 $X2=0
+ $Y2=0
cc_1016 N_A_2008_48#_c_1520_n N_A_1747_74#_c_1651_n 0.0023753f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_1017 N_A_2008_48#_c_1521_n N_A_1747_74#_c_1651_n 0.00741302f $X=11.12 $Y=0.55
+ $X2=0 $Y2=0
cc_1018 N_A_2008_48#_c_1518_n N_A_1747_74#_c_1652_n 0.00406259f $X=11.675
+ $Y=0.665 $X2=0 $Y2=0
cc_1019 N_A_2008_48#_c_1520_n N_A_1747_74#_c_1652_n 0.00385495f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_1020 N_A_2008_48#_c_1521_n N_A_1747_74#_c_1652_n 0.00768727f $X=11.12 $Y=0.55
+ $X2=0 $Y2=0
cc_1021 N_A_2008_48#_c_1528_n N_A_1747_74#_c_1663_n 0.00562099f $X=11.02
+ $Y=2.655 $X2=0 $Y2=0
cc_1022 N_A_2008_48#_c_1532_n N_A_1747_74#_c_1663_n 0.00739298f $X=11.13
+ $Y=2.405 $X2=0 $Y2=0
cc_1023 N_A_2008_48#_c_1529_n N_A_1747_74#_c_1664_n 0.0105765f $X=11.32 $Y=2.32
+ $X2=0 $Y2=0
cc_1024 N_A_2008_48#_c_1530_n N_A_1747_74#_c_1664_n 0.00277596f $X=11.675
+ $Y=1.715 $X2=0 $Y2=0
cc_1025 N_A_2008_48#_c_1519_n N_A_1747_74#_c_1664_n 0.00167941f $X=11.405
+ $Y=1.715 $X2=0 $Y2=0
cc_1026 N_A_2008_48#_c_1529_n N_A_1747_74#_c_1665_n 6.41559e-19 $X=11.32 $Y=2.32
+ $X2=0 $Y2=0
cc_1027 N_A_2008_48#_c_1530_n N_A_1747_74#_c_1665_n 3.71546e-19 $X=11.675
+ $Y=1.715 $X2=0 $Y2=0
cc_1028 N_A_2008_48#_c_1520_n N_A_1747_74#_c_1654_n 0.00507794f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_1029 N_A_2008_48#_c_1521_n N_A_1747_74#_c_1654_n 0.00413357f $X=11.12 $Y=0.55
+ $X2=0 $Y2=0
cc_1030 N_A_2008_48#_c_1518_n N_A_1747_74#_c_1656_n 0.00447579f $X=11.675
+ $Y=0.665 $X2=0 $Y2=0
cc_1031 N_A_2008_48#_c_1530_n N_A_1747_74#_c_1656_n 0.0228154f $X=11.675
+ $Y=1.715 $X2=0 $Y2=0
cc_1032 N_A_2008_48#_c_1519_n N_A_1747_74#_c_1656_n 0.00406088f $X=11.405
+ $Y=1.715 $X2=0 $Y2=0
cc_1033 N_A_2008_48#_c_1520_n N_A_1747_74#_c_1656_n 0.0258377f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_1034 N_A_2008_48#_c_1529_n N_A_1747_74#_c_1670_n 0.00434917f $X=11.32 $Y=2.32
+ $X2=0 $Y2=0
cc_1035 N_A_2008_48#_c_1532_n N_A_1747_74#_c_1670_n 0.00686891f $X=11.13
+ $Y=2.405 $X2=0 $Y2=0
cc_1036 N_A_2008_48#_M1003_g N_A_1747_74#_c_1681_n 0.00100303f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_1037 N_A_2008_48#_c_1524_n N_A_1747_74#_c_1672_n 0.00888546f $X=10.16 $Y=2.37
+ $X2=0 $Y2=0
cc_1038 N_A_2008_48#_c_1527_n N_A_1747_74#_c_1672_n 0.00364065f $X=10.525
+ $Y=2.405 $X2=0 $Y2=0
cc_1039 N_A_2008_48#_M1003_g N_A_1747_74#_c_1659_n 0.00151652f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_1040 N_A_2008_48#_M1003_g N_A_1747_74#_c_1660_n 0.00175137f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_1041 N_A_2008_48#_c_1516_n N_A_1747_74#_c_1660_n 0.0146343f $X=10.16 $Y=1.98
+ $X2=0 $Y2=0
cc_1042 N_A_2008_48#_c_1523_n N_A_1747_74#_c_1660_n 0.0045792f $X=10.16 $Y=2.28
+ $X2=0 $Y2=0
cc_1043 N_A_2008_48#_c_1524_n N_A_1747_74#_c_1660_n 0.00266565f $X=10.16 $Y=2.37
+ $X2=0 $Y2=0
cc_1044 N_A_2008_48#_c_1517_n N_A_1747_74#_c_1660_n 0.0472402f $X=10.36 $Y=1.815
+ $X2=0 $Y2=0
cc_1045 N_A_2008_48#_c_1527_n N_A_1747_74#_c_1660_n 0.00840223f $X=10.525
+ $Y=2.405 $X2=0 $Y2=0
cc_1046 N_A_2008_48#_M1003_g N_A_1747_74#_c_1661_n 0.00782885f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_1047 N_A_2008_48#_M1003_g N_A_1747_74#_c_1662_n 0.0151836f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_1048 N_A_2008_48#_c_1516_n N_A_1747_74#_c_1662_n 0.00516648f $X=10.16 $Y=1.98
+ $X2=0 $Y2=0
cc_1049 N_A_2008_48#_c_1517_n N_A_1747_74#_c_1662_n 0.0174506f $X=10.36 $Y=1.815
+ $X2=0 $Y2=0
cc_1050 N_A_2008_48#_c_1518_n N_A_1747_74#_c_1662_n 0.00792529f $X=11.675
+ $Y=0.665 $X2=0 $Y2=0
cc_1051 N_A_2008_48#_c_1530_n N_A_1747_74#_c_1662_n 0.00127707f $X=11.675
+ $Y=1.715 $X2=0 $Y2=0
cc_1052 N_A_2008_48#_c_1519_n N_A_1747_74#_c_1662_n 0.0125719f $X=11.405
+ $Y=1.715 $X2=0 $Y2=0
cc_1053 N_A_2008_48#_c_1520_n N_A_1747_74#_c_1662_n 0.0245935f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_1054 N_A_2008_48#_c_1521_n N_A_1747_74#_c_1662_n 0.017591f $X=11.12 $Y=0.55
+ $X2=0 $Y2=0
cc_1055 N_A_2008_48#_c_1526_n N_VPWR_M1017_d 0.00157126f $X=10.855 $Y=2.405
+ $X2=0 $Y2=0
cc_1056 N_A_2008_48#_c_1527_n N_VPWR_M1017_d 0.00330343f $X=10.525 $Y=2.405
+ $X2=0 $Y2=0
cc_1057 N_A_2008_48#_c_1532_n N_VPWR_M1041_d 7.76434e-19 $X=11.13 $Y=2.405 $X2=0
+ $Y2=0
cc_1058 N_A_2008_48#_c_1516_n N_VPWR_c_1887_n 6.38002e-19 $X=10.16 $Y=1.98 $X2=0
+ $Y2=0
cc_1059 N_A_2008_48#_c_1524_n N_VPWR_c_1887_n 0.0080003f $X=10.16 $Y=2.37 $X2=0
+ $Y2=0
cc_1060 N_A_2008_48#_c_1526_n N_VPWR_c_1887_n 0.00951507f $X=10.855 $Y=2.405
+ $X2=0 $Y2=0
cc_1061 N_A_2008_48#_c_1527_n N_VPWR_c_1887_n 0.0187155f $X=10.525 $Y=2.405
+ $X2=0 $Y2=0
cc_1062 N_A_2008_48#_c_1528_n N_VPWR_c_1887_n 0.0152062f $X=11.02 $Y=2.655 $X2=0
+ $Y2=0
cc_1063 N_A_2008_48#_c_1528_n N_VPWR_c_1998_n 0.00796791f $X=11.02 $Y=2.655
+ $X2=0 $Y2=0
cc_1064 N_A_2008_48#_c_1529_n N_VPWR_c_1998_n 0.0240111f $X=11.32 $Y=2.32 $X2=0
+ $Y2=0
cc_1065 N_A_2008_48#_c_1530_n N_VPWR_c_1998_n 0.019153f $X=11.675 $Y=1.715 $X2=0
+ $Y2=0
cc_1066 N_A_2008_48#_c_1532_n N_VPWR_c_1998_n 0.0135229f $X=11.13 $Y=2.405 $X2=0
+ $Y2=0
cc_1067 N_A_2008_48#_c_1528_n N_VPWR_c_1896_n 0.00744123f $X=11.02 $Y=2.655
+ $X2=0 $Y2=0
cc_1068 N_A_2008_48#_c_1532_n N_VPWR_c_1896_n 0.00211481f $X=11.13 $Y=2.405
+ $X2=0 $Y2=0
cc_1069 N_A_2008_48#_c_1524_n N_VPWR_c_1899_n 0.00502154f $X=10.16 $Y=2.37 $X2=0
+ $Y2=0
cc_1070 N_A_2008_48#_c_1528_n N_VPWR_c_1900_n 0.0103547f $X=11.02 $Y=2.655 $X2=0
+ $Y2=0
cc_1071 N_A_2008_48#_c_1524_n N_VPWR_c_1881_n 0.00515964f $X=10.16 $Y=2.37 $X2=0
+ $Y2=0
cc_1072 N_A_2008_48#_c_1526_n N_VPWR_c_1881_n 0.00704664f $X=10.855 $Y=2.405
+ $X2=0 $Y2=0
cc_1073 N_A_2008_48#_c_1527_n N_VPWR_c_1881_n 0.00241369f $X=10.525 $Y=2.405
+ $X2=0 $Y2=0
cc_1074 N_A_2008_48#_c_1528_n N_VPWR_c_1881_n 0.011288f $X=11.02 $Y=2.655 $X2=0
+ $Y2=0
cc_1075 N_A_2008_48#_c_1532_n N_VPWR_c_1881_n 0.00672753f $X=11.13 $Y=2.405
+ $X2=0 $Y2=0
cc_1076 N_A_2008_48#_c_1529_n Q_N 0.00264229f $X=11.32 $Y=2.32 $X2=0 $Y2=0
cc_1077 N_A_2008_48#_c_1530_n Q_N 0.0140768f $X=11.675 $Y=1.715 $X2=0 $Y2=0
cc_1078 N_A_2008_48#_c_1520_n Q_N 0.0510002f $X=11.76 $Y=1.63 $X2=0 $Y2=0
cc_1079 N_A_2008_48#_c_1518_n N_VGND_M1006_s 0.00795702f $X=11.675 $Y=0.665
+ $X2=0 $Y2=0
cc_1080 N_A_2008_48#_c_1520_n N_VGND_M1006_s 0.00751007f $X=11.76 $Y=1.63 $X2=0
+ $Y2=0
cc_1081 N_A_2008_48#_M1003_g N_VGND_c_2286_n 0.0106684f $X=10.115 $Y=0.58 $X2=0
+ $Y2=0
cc_1082 N_A_2008_48#_c_1521_n N_VGND_c_2286_n 0.0133829f $X=11.12 $Y=0.55 $X2=0
+ $Y2=0
cc_1083 N_A_2008_48#_M1003_g N_VGND_c_2294_n 0.00383152f $X=10.115 $Y=0.58 $X2=0
+ $Y2=0
cc_1084 N_A_2008_48#_c_1518_n N_VGND_c_2295_n 0.00463151f $X=11.675 $Y=0.665
+ $X2=0 $Y2=0
cc_1085 N_A_2008_48#_c_1521_n N_VGND_c_2295_n 0.0140232f $X=11.12 $Y=0.55 $X2=0
+ $Y2=0
cc_1086 N_A_2008_48#_M1003_g N_VGND_c_2297_n 0.0075694f $X=10.115 $Y=0.58 $X2=0
+ $Y2=0
cc_1087 N_A_2008_48#_c_1518_n N_VGND_c_2297_n 0.00869887f $X=11.675 $Y=0.665
+ $X2=0 $Y2=0
cc_1088 N_A_2008_48#_c_1521_n N_VGND_c_2297_n 0.0117897f $X=11.12 $Y=0.55 $X2=0
+ $Y2=0
cc_1089 N_A_2008_48#_c_1518_n N_VGND_c_2302_n 0.0253659f $X=11.675 $Y=0.665
+ $X2=0 $Y2=0
cc_1090 N_A_2008_48#_c_1521_n N_VGND_c_2302_n 0.00410713f $X=11.12 $Y=0.55 $X2=0
+ $Y2=0
cc_1091 N_A_1747_74#_M1001_g N_A_2513_424#_M1031_g 0.0206457f $X=12.93 $Y=0.645
+ $X2=0 $Y2=0
cc_1092 N_A_1747_74#_c_1668_n N_A_2513_424#_c_1832_n 0.00504987f $X=12.915
+ $Y=1.955 $X2=0 $Y2=0
cc_1093 N_A_1747_74#_c_1669_n N_A_2513_424#_c_1832_n 0.00577491f $X=12.915
+ $Y=2.045 $X2=0 $Y2=0
cc_1094 N_A_1747_74#_M1001_g N_A_2513_424#_c_1832_n 0.0214527f $X=12.93 $Y=0.645
+ $X2=0 $Y2=0
cc_1095 N_A_1747_74#_c_1658_n N_A_2513_424#_c_1832_n 0.00491452f $X=12.915
+ $Y=1.52 $X2=0 $Y2=0
cc_1096 N_A_1747_74#_c_1654_n N_A_2513_424#_c_1833_n 0.00194375f $X=11.965
+ $Y=1.235 $X2=0 $Y2=0
cc_1097 N_A_1747_74#_M1001_g N_A_2513_424#_c_1833_n 0.0144342f $X=12.93 $Y=0.645
+ $X2=0 $Y2=0
cc_1098 N_A_1747_74#_c_1655_n N_A_2513_424#_c_1837_n 0.00842101f $X=12.825
+ $Y=1.52 $X2=0 $Y2=0
cc_1099 N_A_1747_74#_c_1668_n N_A_2513_424#_c_1837_n 0.00946828f $X=12.915
+ $Y=1.955 $X2=0 $Y2=0
cc_1100 N_A_1747_74#_c_1669_n N_A_2513_424#_c_1837_n 0.0176712f $X=12.915
+ $Y=2.045 $X2=0 $Y2=0
cc_1101 N_A_1747_74#_c_1658_n N_A_2513_424#_c_1837_n 0.00107618f $X=12.915
+ $Y=1.52 $X2=0 $Y2=0
cc_1102 N_A_1747_74#_M1001_g N_A_2513_424#_c_1834_n 0.00833371f $X=12.93
+ $Y=0.645 $X2=0 $Y2=0
cc_1103 N_A_1747_74#_c_1658_n N_A_2513_424#_c_1834_n 0.0134227f $X=12.915
+ $Y=1.52 $X2=0 $Y2=0
cc_1104 N_A_1747_74#_c_1655_n N_A_2513_424#_c_1835_n 0.0160046f $X=12.825
+ $Y=1.52 $X2=0 $Y2=0
cc_1105 N_A_1747_74#_c_1656_n N_A_2513_424#_c_1835_n 2.29508e-19 $X=12.04
+ $Y=1.52 $X2=0 $Y2=0
cc_1106 N_A_1747_74#_M1001_g N_A_2513_424#_c_1835_n 0.00105416f $X=12.93
+ $Y=0.645 $X2=0 $Y2=0
cc_1107 N_A_1747_74#_c_1658_n N_A_2513_424#_c_1835_n 7.76856e-19 $X=12.915
+ $Y=1.52 $X2=0 $Y2=0
cc_1108 N_A_1747_74#_c_1672_n N_VPWR_c_1887_n 0.00666746f $X=9.925 $Y=2.59 $X2=0
+ $Y2=0
cc_1109 N_A_1747_74#_c_1665_n N_VPWR_c_1888_n 0.007084f $X=11.925 $Y=1.765 $X2=0
+ $Y2=0
cc_1110 N_A_1747_74#_c_1663_n N_VPWR_c_1998_n 0.00224083f $X=11.245 $Y=2.37
+ $X2=0 $Y2=0
cc_1111 N_A_1747_74#_c_1664_n N_VPWR_c_1998_n 0.00306886f $X=11.35 $Y=2.22 $X2=0
+ $Y2=0
cc_1112 N_A_1747_74#_c_1656_n N_VPWR_c_1998_n 0.00131549f $X=12.04 $Y=1.52 $X2=0
+ $Y2=0
cc_1113 N_A_1747_74#_c_1668_n N_VPWR_c_1889_n 0.00204598f $X=12.915 $Y=1.955
+ $X2=0 $Y2=0
cc_1114 N_A_1747_74#_c_1669_n N_VPWR_c_1889_n 0.00440242f $X=12.915 $Y=2.045
+ $X2=0 $Y2=0
cc_1115 N_A_1747_74#_c_1663_n N_VPWR_c_1896_n 0.00493443f $X=11.245 $Y=2.37
+ $X2=0 $Y2=0
cc_1116 N_A_1747_74#_c_1670_n N_VPWR_c_1896_n 0.00100251f $X=11.35 $Y=2.295
+ $X2=0 $Y2=0
cc_1117 N_A_1747_74#_c_1672_n N_VPWR_c_1899_n 0.0144557f $X=9.925 $Y=2.59 $X2=0
+ $Y2=0
cc_1118 N_A_1747_74#_c_1673_n N_VPWR_c_1899_n 0.00507318f $X=9.325 $Y=2.59 $X2=0
+ $Y2=0
cc_1119 N_A_1747_74#_c_1663_n N_VPWR_c_1900_n 0.00497687f $X=11.245 $Y=2.37
+ $X2=0 $Y2=0
cc_1120 N_A_1747_74#_c_1665_n N_VPWR_c_1901_n 0.00461464f $X=11.925 $Y=1.765
+ $X2=0 $Y2=0
cc_1121 N_A_1747_74#_c_1669_n N_VPWR_c_1901_n 0.00445602f $X=12.915 $Y=2.045
+ $X2=0 $Y2=0
cc_1122 N_A_1747_74#_c_1663_n N_VPWR_c_1881_n 0.00515964f $X=11.245 $Y=2.37
+ $X2=0 $Y2=0
cc_1123 N_A_1747_74#_c_1665_n N_VPWR_c_1881_n 0.00917882f $X=11.925 $Y=1.765
+ $X2=0 $Y2=0
cc_1124 N_A_1747_74#_c_1669_n N_VPWR_c_1881_n 0.00862843f $X=12.915 $Y=2.045
+ $X2=0 $Y2=0
cc_1125 N_A_1747_74#_c_1672_n N_VPWR_c_1881_n 0.023611f $X=9.925 $Y=2.59 $X2=0
+ $Y2=0
cc_1126 N_A_1747_74#_c_1673_n N_VPWR_c_1881_n 0.00697584f $X=9.325 $Y=2.59 $X2=0
+ $Y2=0
cc_1127 N_A_1747_74#_c_1672_n A_1969_489# 0.0021089f $X=9.925 $Y=2.59 $X2=-0.19
+ $Y2=-0.245
cc_1128 N_A_1747_74#_c_1665_n Q_N 0.00308691f $X=11.925 $Y=1.765 $X2=0 $Y2=0
cc_1129 N_A_1747_74#_c_1654_n Q_N 0.0192064f $X=11.965 $Y=1.235 $X2=0 $Y2=0
cc_1130 N_A_1747_74#_c_1655_n Q_N 0.0275523f $X=12.825 $Y=1.52 $X2=0 $Y2=0
cc_1131 N_A_1747_74#_c_1656_n Q_N 0.0123682f $X=12.04 $Y=1.52 $X2=0 $Y2=0
cc_1132 N_A_1747_74#_c_1668_n Q_N 0.00153041f $X=12.915 $Y=1.955 $X2=0 $Y2=0
cc_1133 N_A_1747_74#_c_1669_n Q_N 0.00229735f $X=12.915 $Y=2.045 $X2=0 $Y2=0
cc_1134 N_A_1747_74#_M1001_g Q_N 0.00438444f $X=12.93 $Y=0.645 $X2=0 $Y2=0
cc_1135 N_A_1747_74#_c_1651_n N_VGND_c_2286_n 0.00170773f $X=10.905 $Y=0.87
+ $X2=0 $Y2=0
cc_1136 N_A_1747_74#_c_1681_n N_VGND_c_2286_n 0.0133484f $X=9.605 $Y=0.57 $X2=0
+ $Y2=0
cc_1137 N_A_1747_74#_c_1659_n N_VGND_c_2286_n 8.97539e-19 $X=9.69 $Y=1.005 $X2=0
+ $Y2=0
cc_1138 N_A_1747_74#_c_1662_n N_VGND_c_2286_n 0.0179642f $X=11.26 $Y=1.27 $X2=0
+ $Y2=0
cc_1139 N_A_1747_74#_c_1654_n N_VGND_c_2287_n 0.00434272f $X=11.965 $Y=1.235
+ $X2=0 $Y2=0
cc_1140 N_A_1747_74#_M1001_g N_VGND_c_2287_n 0.00461464f $X=12.93 $Y=0.645 $X2=0
+ $Y2=0
cc_1141 N_A_1747_74#_M1001_g N_VGND_c_2288_n 0.0103391f $X=12.93 $Y=0.645 $X2=0
+ $Y2=0
cc_1142 N_A_1747_74#_c_1681_n N_VGND_c_2294_n 0.0196922f $X=9.605 $Y=0.57 $X2=0
+ $Y2=0
cc_1143 N_A_1747_74#_c_1651_n N_VGND_c_2295_n 0.00434272f $X=10.905 $Y=0.87
+ $X2=0 $Y2=0
cc_1144 N_A_1747_74#_c_1651_n N_VGND_c_2297_n 0.00825669f $X=10.905 $Y=0.87
+ $X2=0 $Y2=0
cc_1145 N_A_1747_74#_c_1654_n N_VGND_c_2297_n 0.0083017f $X=11.965 $Y=1.235
+ $X2=0 $Y2=0
cc_1146 N_A_1747_74#_M1001_g N_VGND_c_2297_n 0.00914946f $X=12.93 $Y=0.645 $X2=0
+ $Y2=0
cc_1147 N_A_1747_74#_c_1681_n N_VGND_c_2297_n 0.0208801f $X=9.605 $Y=0.57 $X2=0
+ $Y2=0
cc_1148 N_A_1747_74#_c_1651_n N_VGND_c_2302_n 0.00289541f $X=10.905 $Y=0.87
+ $X2=0 $Y2=0
cc_1149 N_A_1747_74#_c_1654_n N_VGND_c_2302_n 0.00583402f $X=11.965 $Y=1.235
+ $X2=0 $Y2=0
cc_1150 N_A_2513_424#_c_1832_n N_VPWR_c_1889_n 0.00624321f $X=13.435 $Y=1.765
+ $X2=0 $Y2=0
cc_1151 N_A_2513_424#_c_1837_n N_VPWR_c_1889_n 0.0507962f $X=12.69 $Y=2.265
+ $X2=0 $Y2=0
cc_1152 N_A_2513_424#_c_1834_n N_VPWR_c_1889_n 0.0222736f $X=13.38 $Y=1.465
+ $X2=0 $Y2=0
cc_1153 N_A_2513_424#_c_1837_n N_VPWR_c_1901_n 0.0125859f $X=12.69 $Y=2.265
+ $X2=0 $Y2=0
cc_1154 N_A_2513_424#_c_1832_n N_VPWR_c_1902_n 0.00461464f $X=13.435 $Y=1.765
+ $X2=0 $Y2=0
cc_1155 N_A_2513_424#_c_1832_n N_VPWR_c_1881_n 0.0091238f $X=13.435 $Y=1.765
+ $X2=0 $Y2=0
cc_1156 N_A_2513_424#_c_1837_n N_VPWR_c_1881_n 0.0103846f $X=12.69 $Y=2.265
+ $X2=0 $Y2=0
cc_1157 N_A_2513_424#_c_1833_n Q_N 0.0571733f $X=12.715 $Y=0.645 $X2=0 $Y2=0
cc_1158 N_A_2513_424#_c_1837_n Q_N 0.0895806f $X=12.69 $Y=2.265 $X2=0 $Y2=0
cc_1159 N_A_2513_424#_c_1835_n Q_N 0.0215198f $X=12.712 $Y=1.465 $X2=0 $Y2=0
cc_1160 N_A_2513_424#_M1031_g Q 0.00811057f $X=13.42 $Y=0.74 $X2=0 $Y2=0
cc_1161 N_A_2513_424#_M1031_g Q 0.00301691f $X=13.42 $Y=0.74 $X2=0 $Y2=0
cc_1162 N_A_2513_424#_c_1832_n Q 0.00230594f $X=13.435 $Y=1.765 $X2=0 $Y2=0
cc_1163 N_A_2513_424#_c_1834_n Q 0.00111755f $X=13.38 $Y=1.465 $X2=0 $Y2=0
cc_1164 N_A_2513_424#_c_1832_n Q 0.00190204f $X=13.435 $Y=1.765 $X2=0 $Y2=0
cc_1165 N_A_2513_424#_M1031_g N_Q_c_2265_n 0.0040915f $X=13.42 $Y=0.74 $X2=0
+ $Y2=0
cc_1166 N_A_2513_424#_c_1832_n N_Q_c_2265_n 0.0129497f $X=13.435 $Y=1.765 $X2=0
+ $Y2=0
cc_1167 N_A_2513_424#_c_1834_n N_Q_c_2265_n 0.0250949f $X=13.38 $Y=1.465 $X2=0
+ $Y2=0
cc_1168 N_A_2513_424#_c_1833_n N_VGND_c_2287_n 0.00778672f $X=12.715 $Y=0.645
+ $X2=0 $Y2=0
cc_1169 N_A_2513_424#_M1031_g N_VGND_c_2288_n 0.00330159f $X=13.42 $Y=0.74 $X2=0
+ $Y2=0
cc_1170 N_A_2513_424#_c_1832_n N_VGND_c_2288_n 0.00172388f $X=13.435 $Y=1.765
+ $X2=0 $Y2=0
cc_1171 N_A_2513_424#_c_1833_n N_VGND_c_2288_n 0.035427f $X=12.715 $Y=0.645
+ $X2=0 $Y2=0
cc_1172 N_A_2513_424#_c_1834_n N_VGND_c_2288_n 0.0145561f $X=13.38 $Y=1.465
+ $X2=0 $Y2=0
cc_1173 N_A_2513_424#_M1031_g N_VGND_c_2296_n 0.00434272f $X=13.42 $Y=0.74 $X2=0
+ $Y2=0
cc_1174 N_A_2513_424#_M1031_g N_VGND_c_2297_n 0.00824587f $X=13.42 $Y=0.74 $X2=0
+ $Y2=0
cc_1175 N_A_2513_424#_c_1833_n N_VGND_c_2297_n 0.00976756f $X=12.715 $Y=0.645
+ $X2=0 $Y2=0
cc_1176 N_VPWR_c_1897_n N_A_409_81#_c_2085_n 0.00497007f $X=3.095 $Y=3.33 $X2=0
+ $Y2=0
cc_1177 N_VPWR_c_1881_n N_A_409_81#_c_2085_n 0.0104121f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1178 N_VPWR_M1023_d N_A_409_81#_c_2107_n 0.0109237f $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1179 N_VPWR_c_1883_n N_A_409_81#_c_2107_n 0.0213202f $X=3.26 $Y=2.815 $X2=0
+ $Y2=0
cc_1180 N_VPWR_c_1881_n N_A_409_81#_c_2107_n 0.00646454f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1181 N_VPWR_c_1892_n N_A_409_81#_c_2076_n 0.00543175f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1182 N_VPWR_c_1881_n N_A_409_81#_c_2076_n 0.0102994f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1183 N_VPWR_M1023_d N_A_409_81#_c_2077_n 0.0014741f $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1184 N_VPWR_c_1892_n N_A_409_81#_c_2077_n 0.00409815f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1185 N_VPWR_c_1881_n N_A_409_81#_c_2077_n 0.0149416f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1186 N_VPWR_M1024_d N_A_409_81#_c_2078_n 0.00387164f $X=4.72 $Y=1.96 $X2=0
+ $Y2=0
cc_1187 N_VPWR_c_1884_n N_A_409_81#_c_2078_n 0.0167709f $X=4.87 $Y=2.835 $X2=0
+ $Y2=0
cc_1188 N_VPWR_c_1892_n N_A_409_81#_c_2078_n 7.54393e-19 $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1189 N_VPWR_c_1894_n N_A_409_81#_c_2078_n 0.0103722f $X=7.025 $Y=3.33 $X2=0
+ $Y2=0
cc_1190 N_VPWR_c_1881_n N_A_409_81#_c_2078_n 0.0213354f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1191 N_VPWR_c_1894_n N_A_409_81#_c_2079_n 0.00535093f $X=7.025 $Y=3.33 $X2=0
+ $Y2=0
cc_1192 N_VPWR_c_1881_n N_A_409_81#_c_2079_n 0.00675054f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1193 N_VPWR_c_1882_n N_A_409_81#_c_2083_n 0.0176046f $X=1.39 $Y=2.475 $X2=0
+ $Y2=0
cc_1194 N_VPWR_c_1883_n N_A_409_81#_c_2083_n 0.00746073f $X=3.26 $Y=2.815 $X2=0
+ $Y2=0
cc_1195 N_VPWR_c_1897_n N_A_409_81#_c_2083_n 0.0197634f $X=3.095 $Y=3.33 $X2=0
+ $Y2=0
cc_1196 N_VPWR_c_1881_n N_A_409_81#_c_2083_n 0.016073f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1197 N_VPWR_c_1883_n N_A_409_81#_c_2084_n 0.014926f $X=3.26 $Y=2.815 $X2=0
+ $Y2=0
cc_1198 N_VPWR_c_1892_n N_A_409_81#_c_2084_n 0.0144865f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1199 N_VPWR_c_1881_n N_A_409_81#_c_2084_n 0.012005f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1200 N_VPWR_c_1888_n Q_N 0.00144265f $X=11.592 $Y=3.245 $X2=0 $Y2=0
cc_1201 N_VPWR_c_1901_n Q_N 0.0146357f $X=13.045 $Y=3.33 $X2=0 $Y2=0
cc_1202 N_VPWR_c_1881_n Q_N 0.0121141f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1203 N_VPWR_c_1889_n Q 0.00249543f $X=13.21 $Y=1.985 $X2=0 $Y2=0
cc_1204 N_VPWR_c_1902_n Q 0.0124046f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1205 N_VPWR_c_1881_n Q 0.0102675f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1206 N_A_409_81#_c_2085_n A_512_464# 0.0111613f $X=2.84 $Y=2.495 $X2=-0.19
+ $Y2=-0.245
cc_1207 N_A_409_81#_c_2116_n A_512_464# 0.00319536f $X=2.945 $Y=2.495 $X2=-0.19
+ $Y2=-0.245
cc_1208 N_A_409_81#_M1012_d N_noxref_25_c_2422_n 0.00874665f $X=2.045 $Y=0.405
+ $X2=0 $Y2=0
cc_1209 N_A_409_81#_c_2067_n N_noxref_25_c_2422_n 0.0126305f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1210 N_A_409_81#_c_2074_n N_noxref_25_c_2422_n 0.019982f $X=2.435 $Y=0.68
+ $X2=0 $Y2=0
cc_1211 N_A_409_81#_c_2067_n N_noxref_25_c_2424_n 0.0234737f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1212 N_A_409_81#_c_2074_n N_noxref_25_c_2424_n 0.00520956f $X=2.435 $Y=0.68
+ $X2=0 $Y2=0
cc_1213 Q_N N_VGND_c_2287_n 0.0145639f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1214 Q_N N_VGND_c_2297_n 0.0119984f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1215 Q_N N_VGND_c_2302_n 0.00297405f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1216 Q N_VGND_c_2288_n 0.0297276f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1217 Q N_VGND_c_2296_n 0.0161257f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1218 Q N_VGND_c_2297_n 0.013291f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1219 N_VGND_c_2283_n N_noxref_25_c_2421_n 0.0253895f $X=0.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1220 N_VGND_c_2292_n N_noxref_25_c_2422_n 0.109804f $X=3.59 $Y=0 $X2=0 $Y2=0
cc_1221 N_VGND_c_2297_n N_noxref_25_c_2422_n 0.0641003f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1222 N_VGND_c_2283_n N_noxref_25_c_2423_n 0.0121617f $X=0.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1223 N_VGND_c_2292_n N_noxref_25_c_2423_n 0.0176516f $X=3.59 $Y=0 $X2=0 $Y2=0
cc_1224 N_VGND_c_2297_n N_noxref_25_c_2423_n 0.00966868f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1225 N_VGND_c_2284_n N_noxref_25_c_2424_n 0.0118481f $X=3.715 $Y=0.565 $X2=0
+ $Y2=0
cc_1226 N_VGND_c_2292_n N_noxref_25_c_2424_n 0.0243596f $X=3.59 $Y=0 $X2=0 $Y2=0
cc_1227 N_VGND_c_2297_n N_noxref_25_c_2424_n 0.0134194f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1228 N_noxref_25_c_2422_n noxref_26 0.00334264f $X=3.06 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1229 N_noxref_25_c_2422_n noxref_27 0.00226367f $X=3.06 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
