* File: sky130_fd_sc_ls__nor4bb_4.pex.spice
* Created: Fri Aug 28 13:41:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NOR4BB_4%B 1 3 6 10 12 14 15 17 20 22 24 27 29 34 36
+ 41 48 57
c120 29 0 1.77894e-19 $X=1.085 $Y=1.485
c121 12 0 1.12408e-19 $X=3 $Y=1.67
r122 57 58 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=3.95 $Y=1.462
+ $X2=3.965 $Y2=1.462
r123 54 55 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=3.45 $Y=1.462
+ $X2=3.465 $Y2=1.462
r124 51 52 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=2.985 $Y=1.462
+ $X2=3 $Y2=1.462
r125 48 63 6.51381 $w=2.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.795
r126 42 57 25.4027 $w=3.7e-07 $l=1.95e-07 $layer=POLY_cond $X=3.755 $Y=1.462
+ $X2=3.95 $Y2=1.462
r127 42 55 37.7784 $w=3.7e-07 $l=2.9e-07 $layer=POLY_cond $X=3.755 $Y=1.462
+ $X2=3.465 $Y2=1.462
r128 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.755
+ $Y=1.42 $X2=3.755 $Y2=1.42
r129 39 54 48.8514 $w=3.7e-07 $l=3.75e-07 $layer=POLY_cond $X=3.075 $Y=1.462
+ $X2=3.45 $Y2=1.462
r130 39 52 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.075 $Y=1.462
+ $X2=3 $Y2=1.462
r131 38 41 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.075 $Y=1.42
+ $X2=3.755 $Y2=1.42
r132 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.075
+ $Y=1.42 $X2=3.075 $Y2=1.42
r133 36 46 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.805 $Y=1.42
+ $X2=2.805 $Y2=1.795
r134 36 38 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.89 $Y=1.42
+ $X2=3.075 $Y2=1.42
r135 35 63 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.315 $Y=1.795
+ $X2=1.2 $Y2=1.795
r136 34 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.72 $Y=1.795
+ $X2=2.805 $Y2=1.795
r137 34 35 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=2.72 $Y=1.795
+ $X2=1.315 $Y2=1.795
r138 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.43
+ $Y=1.485 $X2=0.43 $Y2=1.485
r139 29 48 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.2 $Y=1.485
+ $X2=1.2 $Y2=1.665
r140 29 31 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=1.085 $Y=1.485
+ $X2=0.43 $Y2=1.485
r141 25 58 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.965 $Y=1.255
+ $X2=3.965 $Y2=1.462
r142 25 27 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=3.965 $Y=1.255
+ $X2=3.965 $Y2=0.74
r143 22 57 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.95 $Y=1.67
+ $X2=3.95 $Y2=1.462
r144 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.95 $Y=1.67
+ $X2=3.95 $Y2=2.305
r145 18 55 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.465 $Y=1.255
+ $X2=3.465 $Y2=1.462
r146 18 20 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=3.465 $Y=1.255
+ $X2=3.465 $Y2=0.74
r147 15 54 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.45 $Y=1.67
+ $X2=3.45 $Y2=1.462
r148 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.45 $Y=1.67
+ $X2=3.45 $Y2=2.305
r149 12 52 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3 $Y=1.67 $X2=3
+ $Y2=1.462
r150 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3 $Y=1.67 $X2=3
+ $Y2=2.305
r151 8 51 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.985 $Y=1.255
+ $X2=2.985 $Y2=1.462
r152 8 10 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=2.985 $Y=1.255
+ $X2=2.985 $Y2=0.74
r153 4 32 38.535 $w=3.06e-07 $l=2.14173e-07 $layer=POLY_cond $X=0.565 $Y=1.32
+ $X2=0.452 $Y2=1.485
r154 4 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.565 $Y=1.32
+ $X2=0.565 $Y2=0.74
r155 1 32 56.6494 $w=3.06e-07 $l=3.05352e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.452 $Y2=1.485
r156 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 26 27 28 31 34
c94 31 0 3.21438e-20 $X=2.07 $Y=1.385
c95 7 0 1.77894e-19 $X=1.505 $Y=1.765
c96 4 0 1.44527e-19 $X=1.005 $Y=1.765
r97 41 43 0.561772 $w=4.29e-07 $l=5e-09 $layer=POLY_cond $X=1.99 $Y=1.492
+ $X2=1.995 $Y2=1.492
r98 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.99
+ $Y=1.385 $X2=1.99 $Y2=1.385
r99 39 41 3.9324 $w=4.29e-07 $l=3.5e-08 $layer=POLY_cond $X=1.955 $Y=1.492
+ $X2=1.99 $Y2=1.492
r100 38 39 48.8741 $w=4.29e-07 $l=4.35e-07 $layer=POLY_cond $X=1.52 $Y=1.492
+ $X2=1.955 $Y2=1.492
r101 37 38 1.68531 $w=4.29e-07 $l=1.5e-08 $layer=POLY_cond $X=1.505 $Y=1.492
+ $X2=1.52 $Y2=1.492
r102 36 37 56.1772 $w=4.29e-07 $l=5e-07 $layer=POLY_cond $X=1.005 $Y=1.492
+ $X2=1.505 $Y2=1.492
r103 35 36 1.12354 $w=4.29e-07 $l=1e-08 $layer=POLY_cond $X=0.995 $Y=1.492
+ $X2=1.005 $Y2=1.492
r104 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.33
+ $Y=1.385 $X2=2.33 $Y2=1.385
r105 31 43 11.1166 $w=4.29e-07 $l=1.39549e-07 $layer=POLY_cond $X=2.07 $Y=1.385
+ $X2=1.995 $Y2=1.492
r106 31 33 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=2.07 $Y=1.385
+ $X2=2.33 $Y2=1.385
r107 28 34 5.44209 $w=3.58e-07 $l=1.7e-07 $layer=LI1_cond $X=2.16 $Y=1.36
+ $X2=2.33 $Y2=1.36
r108 28 42 5.44209 $w=3.58e-07 $l=1.7e-07 $layer=LI1_cond $X=2.16 $Y=1.36
+ $X2=1.99 $Y2=1.36
r109 27 42 9.92381 $w=3.58e-07 $l=3.1e-07 $layer=LI1_cond $X=1.68 $Y=1.36
+ $X2=1.99 $Y2=1.36
r110 26 33 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.405 $Y=1.385
+ $X2=2.33 $Y2=1.385
r111 22 26 43.4747 $w=1.95e-07 $l=1.78452e-07 $layer=POLY_cond $X=2.535 $Y=1.22
+ $X2=2.507 $Y2=1.385
r112 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.535 $Y=1.22
+ $X2=2.535 $Y2=0.74
r113 19 26 96.6183 $w=1.95e-07 $l=3.85953e-07 $layer=POLY_cond $X=2.495 $Y=1.765
+ $X2=2.507 $Y2=1.385
r114 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.495 $Y=1.765
+ $X2=2.495 $Y2=2.4
r115 16 43 27.5819 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.995 $Y=1.22
+ $X2=1.995 $Y2=1.492
r116 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.995 $Y=1.22
+ $X2=1.995 $Y2=0.74
r117 13 39 27.5819 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.955 $Y2=1.492
r118 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.955 $Y2=2.4
r119 10 38 27.5819 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.52 $Y=1.22
+ $X2=1.52 $Y2=1.492
r120 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.52 $Y=1.22
+ $X2=1.52 $Y2=0.74
r121 7 37 27.5819 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=1.492
r122 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=2.4
r123 4 36 27.5819 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=1.492
r124 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r125 1 35 27.5819 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.995 $Y=1.22
+ $X2=0.995 $Y2=1.492
r126 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.995 $Y=1.22
+ $X2=0.995 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_4%A_864_48# 1 2 9 11 13 14 16 19 23 25 27 28
+ 30 31 33 37 38 39 44 45 46 47 49 50 51 55 56 57 58 59 63 67 72 74 82
c181 56 0 1.90324e-19 $X=8.71 $Y=1.385
c182 44 0 7.33604e-20 $X=5.27 $Y=1.585
c183 31 0 1.65916e-19 $X=8.11 $Y=1.22
c184 11 0 6.57076e-20 $X=4.41 $Y=1.67
r185 79 80 4.4748 $w=3.77e-07 $l=3.5e-08 $layer=POLY_cond $X=4.86 $Y=1.462
+ $X2=4.895 $Y2=1.462
r186 76 77 1.91777 $w=3.77e-07 $l=1.5e-08 $layer=POLY_cond $X=4.395 $Y=1.462
+ $X2=4.41 $Y2=1.462
r187 74 80 10.4633 $w=3.77e-07 $l=9.3675e-08 $layer=POLY_cond $X=4.97 $Y=1.42
+ $X2=4.895 $Y2=1.462
r188 72 73 16.3921 $w=2.27e-07 $l=3.05e-07 $layer=LI1_cond $X=8.71 $Y=1.81
+ $X2=8.71 $Y2=2.115
r189 71 74 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=5.19 $Y=1.42
+ $X2=4.97 $Y2=1.42
r190 70 71 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.19
+ $Y=1.42 $X2=5.19 $Y2=1.42
r191 65 67 2.72396 $w=2.73e-07 $l=6.5e-08 $layer=LI1_cond $X=9.437 $Y=2.2
+ $X2=9.437 $Y2=2.265
r192 61 63 12.5882 $w=3.23e-07 $l=3.55e-07 $layer=LI1_cond $X=9.422 $Y=1.19
+ $X2=9.422 $Y2=0.835
r193 60 73 2.43258 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.875 $Y=2.115
+ $X2=8.71 $Y2=2.115
r194 59 65 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=9.3 $Y=2.115
+ $X2=9.437 $Y2=2.2
r195 59 60 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.3 $Y=2.115
+ $X2=8.875 $Y2=2.115
r196 57 61 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=9.26 $Y=1.275
+ $X2=9.422 $Y2=1.19
r197 57 58 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.26 $Y=1.275
+ $X2=8.875 $Y2=1.275
r198 56 82 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.71 $Y=1.385
+ $X2=8.545 $Y2=1.385
r199 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.71
+ $Y=1.385 $X2=8.71 $Y2=1.385
r200 53 72 4.34093 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.71 $Y=1.725
+ $X2=8.71 $Y2=1.81
r201 53 55 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.71 $Y=1.725
+ $X2=8.71 $Y2=1.385
r202 52 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.71 $Y=1.36
+ $X2=8.875 $Y2=1.275
r203 52 55 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=8.71 $Y=1.36
+ $X2=8.71 $Y2=1.385
r204 50 72 2.43258 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.545 $Y=1.81
+ $X2=8.71 $Y2=1.81
r205 50 51 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=8.545 $Y=1.81
+ $X2=7.57 $Y2=1.81
r206 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.485 $Y=1.895
+ $X2=7.57 $Y2=1.81
r207 48 49 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.485 $Y=1.895
+ $X2=7.485 $Y2=2.225
r208 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.4 $Y=2.31
+ $X2=7.485 $Y2=2.225
r209 46 47 133.417 $w=1.68e-07 $l=2.045e-06 $layer=LI1_cond $X=7.4 $Y=2.31
+ $X2=5.355 $Y2=2.31
r210 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.27 $Y=2.225
+ $X2=5.355 $Y2=2.31
r211 44 70 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.27 $Y=1.585
+ $X2=5.27 $Y2=1.42
r212 44 45 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.27 $Y=1.585
+ $X2=5.27 $Y2=2.225
r213 42 79 44.748 $w=3.77e-07 $l=3.5e-07 $layer=POLY_cond $X=4.51 $Y=1.462
+ $X2=4.86 $Y2=1.462
r214 42 77 12.7851 $w=3.77e-07 $l=1e-07 $layer=POLY_cond $X=4.51 $Y=1.462
+ $X2=4.41 $Y2=1.462
r215 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.51
+ $Y=1.42 $X2=4.51 $Y2=1.42
r216 39 70 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.185 $Y=1.42
+ $X2=5.27 $Y2=1.42
r217 39 41 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.185 $Y=1.42
+ $X2=4.51 $Y2=1.42
r218 37 71 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=5.32 $Y=1.42
+ $X2=5.19 $Y2=1.42
r219 35 38 4.4846 $w=3.15e-07 $l=1.19248e-07 $layer=POLY_cond $X=8.185 $Y=1.377
+ $X2=8.095 $Y2=1.445
r220 35 82 65.9477 $w=3.15e-07 $l=3.6e-07 $layer=POLY_cond $X=8.185 $Y=1.377
+ $X2=8.545 $Y2=1.377
r221 31 38 35.9208 $w=1.5e-07 $l=2.32379e-07 $layer=POLY_cond $X=8.11 $Y=1.22
+ $X2=8.095 $Y2=1.445
r222 31 33 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.11 $Y=1.22
+ $X2=8.11 $Y2=0.74
r223 28 38 35.9208 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=8.095 $Y=1.67
+ $X2=8.095 $Y2=1.445
r224 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.095 $Y=1.67
+ $X2=8.095 $Y2=2.305
r225 25 37 57.5603 $w=2.35e-07 $l=2.66927e-07 $layer=POLY_cond $X=5.48 $Y=1.67
+ $X2=5.445 $Y2=1.42
r226 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.48 $Y=1.67
+ $X2=5.48 $Y2=2.305
r227 21 37 40.1263 $w=2.35e-07 $l=1.88348e-07 $layer=POLY_cond $X=5.395 $Y=1.255
+ $X2=5.445 $Y2=1.42
r228 21 23 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=5.395 $Y=1.255
+ $X2=5.395 $Y2=0.74
r229 17 80 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.895 $Y=1.255
+ $X2=4.895 $Y2=1.462
r230 17 19 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=4.895 $Y=1.255
+ $X2=4.895 $Y2=0.74
r231 14 79 24.4204 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.86 $Y=1.67
+ $X2=4.86 $Y2=1.462
r232 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.86 $Y=1.67
+ $X2=4.86 $Y2=2.305
r233 11 77 24.4204 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.41 $Y=1.67
+ $X2=4.41 $Y2=1.462
r234 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.41 $Y=1.67
+ $X2=4.41 $Y2=2.305
r235 7 76 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.395 $Y=1.255
+ $X2=4.395 $Y2=1.462
r236 7 9 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=4.395 $Y=1.255
+ $X2=4.395 $Y2=0.74
r237 2 67 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=9.26
+ $Y=2.12 $X2=9.41 $Y2=2.265
r238 1 63 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=9.28
+ $Y=0.37 $X2=9.42 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_4%A_1162_48# 1 2 9 12 13 15 16 19 20 22 25 27
+ 29 31 32 34 35 37 38 40 41 42 43 50 52 53 54 56 57 58 60 61 62 65 67 68 71 74
+ 75
c192 68 0 1.64824e-19 $X=10.395 $Y=2.035
c193 43 0 1.20663e-19 $X=8.205 $Y=1.39
c194 41 0 7.33604e-20 $X=5.915 $Y=1.33
c195 9 0 1.59971e-19 $X=5.885 $Y=0.74
r196 76 77 1.95935 $w=3.69e-07 $l=1.5e-08 $layer=POLY_cond $X=6.825 $Y=1.447
+ $X2=6.84 $Y2=1.447
r197 73 75 4.23118 $w=2.15e-07 $l=1.05119e-07 $layer=LI1_cond $X=10.84 $Y=1.28
+ $X2=10.795 $Y2=1.195
r198 73 74 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.84 $Y=1.28
+ $X2=10.84 $Y2=1.95
r199 69 75 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=10.795 $Y=1.11
+ $X2=10.795 $Y2=1.195
r200 69 71 26.3732 $w=2.58e-07 $l=5.95e-07 $layer=LI1_cond $X=10.795 $Y=1.11
+ $X2=10.795 $Y2=0.515
r201 67 74 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.755 $Y=2.035
+ $X2=10.84 $Y2=1.95
r202 67 68 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=10.755 $Y=2.035
+ $X2=10.395 $Y2=2.035
r203 63 68 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.27 $Y=2.12
+ $X2=10.395 $Y2=2.035
r204 63 65 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=10.27 $Y=2.12
+ $X2=10.27 $Y2=2.265
r205 61 75 2.20034 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.665 $Y=1.195
+ $X2=10.795 $Y2=1.195
r206 61 62 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=10.665 $Y=1.195
+ $X2=9.925 $Y2=1.195
r207 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.84 $Y=1.11
+ $X2=9.925 $Y2=1.195
r208 59 60 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=9.84 $Y=0.425
+ $X2=9.84 $Y2=1.11
r209 57 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.755 $Y=0.34
+ $X2=9.84 $Y2=0.425
r210 57 58 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=9.755 $Y=0.34
+ $X2=9.09 $Y2=0.34
r211 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.005 $Y=0.425
+ $X2=9.09 $Y2=0.34
r212 55 56 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.005 $Y=0.425
+ $X2=9.005 $Y2=0.85
r213 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.92 $Y=0.935
+ $X2=9.005 $Y2=0.85
r214 53 54 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=8.92 $Y=0.935
+ $X2=8.375 $Y2=0.935
r215 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.29 $Y=1.02
+ $X2=8.375 $Y2=0.935
r216 51 52 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.29 $Y=1.02
+ $X2=8.29 $Y2=1.225
r217 50 81 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=7.63 $Y=1.447
+ $X2=7.655 $Y2=1.447
r218 50 79 44.4119 $w=3.69e-07 $l=3.4e-07 $layer=POLY_cond $X=7.63 $Y=1.447
+ $X2=7.29 $Y2=1.447
r219 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.63
+ $Y=1.39 $X2=7.63 $Y2=1.39
r220 46 79 44.4119 $w=3.69e-07 $l=3.4e-07 $layer=POLY_cond $X=6.95 $Y=1.447
+ $X2=7.29 $Y2=1.447
r221 46 77 14.3686 $w=3.69e-07 $l=1.1e-07 $layer=POLY_cond $X=6.95 $Y=1.447
+ $X2=6.84 $Y2=1.447
r222 45 49 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.95 $Y=1.39
+ $X2=7.63 $Y2=1.39
r223 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.95
+ $Y=1.39 $X2=6.95 $Y2=1.39
r224 43 52 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.205 $Y=1.39
+ $X2=8.29 $Y2=1.225
r225 43 49 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=8.205 $Y=1.39
+ $X2=7.63 $Y2=1.39
r226 38 81 23.9013 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=7.655 $Y=1.225
+ $X2=7.655 $Y2=1.447
r227 38 40 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=7.655 $Y=1.225
+ $X2=7.655 $Y2=0.74
r228 35 79 23.9013 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.29 $Y=1.67
+ $X2=7.29 $Y2=1.447
r229 35 37 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.29 $Y=1.67
+ $X2=7.29 $Y2=2.305
r230 32 77 23.9013 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.84 $Y=1.67
+ $X2=6.84 $Y2=1.447
r231 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.84 $Y=1.67
+ $X2=6.84 $Y2=2.305
r232 29 76 23.9013 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.825 $Y=1.225
+ $X2=6.825 $Y2=1.447
r233 29 31 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.825 $Y=1.225
+ $X2=6.825 $Y2=0.74
r234 28 42 13.2179 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.47 $Y=1.33 $X2=6.38
+ $Y2=1.33
r235 27 76 27.2843 $w=3.69e-07 $l=1.4988e-07 $layer=POLY_cond $X=6.75 $Y=1.33
+ $X2=6.825 $Y2=1.447
r236 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.75 $Y=1.33
+ $X2=6.47 $Y2=1.33
r237 23 42 10.9219 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=6.395 $Y=1.255
+ $X2=6.38 $Y2=1.33
r238 23 25 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=6.395 $Y=1.255
+ $X2=6.395 $Y2=0.74
r239 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.38 $Y=1.67
+ $X2=6.38 $Y2=2.305
r240 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.38 $Y=1.58 $X2=6.38
+ $Y2=1.67
r241 18 42 10.9219 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.38 $Y=1.405
+ $X2=6.38 $Y2=1.33
r242 18 19 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=6.38 $Y=1.405
+ $X2=6.38 $Y2=1.58
r243 17 41 6.66866 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=6.02 $Y=1.33
+ $X2=5.915 $Y2=1.33
r244 16 42 13.2179 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.29 $Y=1.33 $X2=6.38
+ $Y2=1.33
r245 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=6.29 $Y=1.33
+ $X2=6.02 $Y2=1.33
r246 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.93 $Y=1.67
+ $X2=5.93 $Y2=2.305
r247 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.93 $Y=1.58 $X2=5.93
+ $Y2=1.67
r248 11 41 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=5.93 $Y=1.405
+ $X2=5.915 $Y2=1.33
r249 11 12 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=5.93 $Y=1.405
+ $X2=5.93 $Y2=1.58
r250 7 41 18.8402 $w=1.65e-07 $l=8.87412e-08 $layer=POLY_cond $X=5.885 $Y=1.255
+ $X2=5.915 $Y2=1.33
r251 7 9 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=5.885 $Y=1.255
+ $X2=5.885 $Y2=0.74
r252 2 65 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=10.16
+ $Y=2.12 $X2=10.31 $Y2=2.265
r253 1 71 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.62
+ $Y=0.37 $X2=10.76 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_4%C_N 1 3 6 8 10 11 12 18
c48 18 0 5.00264e-20 $X=9.26 $Y=1.695
c49 12 0 6.96612e-20 $X=9.84 $Y=1.665
c50 8 0 1.64824e-19 $X=9.635 $Y=2.045
r51 18 20 51.6429 $w=3.5e-07 $l=3.75e-07 $layer=POLY_cond $X=9.26 $Y=1.787
+ $X2=9.635 $Y2=1.787
r52 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.26
+ $Y=1.695 $X2=9.26 $Y2=1.695
r53 16 18 7.57429 $w=3.5e-07 $l=5.5e-08 $layer=POLY_cond $X=9.205 $Y=1.787
+ $X2=9.26 $Y2=1.787
r54 15 16 2.75429 $w=3.5e-07 $l=2e-08 $layer=POLY_cond $X=9.185 $Y=1.787
+ $X2=9.205 $Y2=1.787
r55 11 12 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=1.695
+ $X2=9.84 $Y2=1.695
r56 11 19 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=9.36 $Y=1.695 $X2=9.26
+ $Y2=1.695
r57 8 20 22.6286 $w=1.5e-07 $l=2.58e-07 $layer=POLY_cond $X=9.635 $Y=2.045
+ $X2=9.635 $Y2=1.787
r58 8 10 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.635 $Y=2.045
+ $X2=9.635 $Y2=2.54
r59 4 16 22.6286 $w=1.5e-07 $l=2.57e-07 $layer=POLY_cond $X=9.205 $Y=1.53
+ $X2=9.205 $Y2=1.787
r60 4 6 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=9.205 $Y=1.53
+ $X2=9.205 $Y2=0.74
r61 1 15 22.6286 $w=1.5e-07 $l=2.58e-07 $layer=POLY_cond $X=9.185 $Y=2.045
+ $X2=9.185 $Y2=1.787
r62 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.185 $Y=2.045
+ $X2=9.185 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_4%D_N 2 3 5 7 8 10 13 15 21
c43 15 0 5.00264e-20 $X=10.32 $Y=1.665
r44 21 22 1.46951 $w=3.28e-07 $l=1e-08 $layer=POLY_cond $X=10.535 $Y=1.615
+ $X2=10.545 $Y2=1.615
r45 19 21 36.003 $w=3.28e-07 $l=2.45e-07 $layer=POLY_cond $X=10.29 $Y=1.615
+ $X2=10.535 $Y2=1.615
r46 17 19 30.125 $w=3.28e-07 $l=2.05e-07 $layer=POLY_cond $X=10.085 $Y=1.615
+ $X2=10.29 $Y2=1.615
r47 15 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.29
+ $Y=1.615 $X2=10.29 $Y2=1.615
r48 11 22 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.545 $Y=1.45
+ $X2=10.545 $Y2=1.615
r49 11 13 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=10.545 $Y=1.45
+ $X2=10.545 $Y2=0.74
r50 8 10 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.535 $Y=2.045
+ $X2=10.535 $Y2=2.54
r51 7 8 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.535 $Y=1.955
+ $X2=10.535 $Y2=2.045
r52 6 21 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.535 $Y=1.78
+ $X2=10.535 $Y2=1.615
r53 6 7 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=10.535 $Y=1.78
+ $X2=10.535 $Y2=1.955
r54 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.085 $Y=2.045
+ $X2=10.085 $Y2=2.54
r55 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.085 $Y=1.955
+ $X2=10.085 $Y2=2.045
r56 1 17 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.085 $Y=1.78
+ $X2=10.085 $Y2=1.615
r57 1 2 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=10.085 $Y=1.78
+ $X2=10.085 $Y2=1.955
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_4%A_27_368# 1 2 3 4 5 18 20 24 26 28 31 32 33
+ 38 41 44
c86 18 0 1.44527e-19 $X=0.28 $Y=2.815
r87 47 48 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.225 $Y=1.89
+ $X2=3.225 $Y2=2.135
r88 44 47 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=3.225 $Y=1.84
+ $X2=3.225 $Y2=1.89
r89 41 43 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.135
r90 36 38 27.2947 $w=2.83e-07 $l=6.75e-07 $layer=LI1_cond $X=8.347 $Y=2.905
+ $X2=8.347 $Y2=2.23
r91 33 35 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=4.26 $Y=2.99 $X2=5.17
+ $Y2=2.99
r92 32 36 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=8.205 $Y=2.99
+ $X2=8.347 $Y2=2.905
r93 32 35 198.005 $w=1.68e-07 $l=3.035e-06 $layer=LI1_cond $X=8.205 $Y=2.99
+ $X2=5.17 $Y2=2.99
r94 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.175 $Y=2.905
+ $X2=4.26 $Y2=2.99
r95 29 31 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.175 $Y=2.905
+ $X2=4.175 $Y2=2.72
r96 28 50 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.175 $Y=1.925
+ $X2=4.175 $Y2=1.84
r97 28 31 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=4.175 $Y=1.925
+ $X2=4.175 $Y2=2.72
r98 27 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.39 $Y=1.84
+ $X2=3.225 $Y2=1.84
r99 26 50 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=1.84
+ $X2=4.175 $Y2=1.84
r100 26 27 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.09 $Y=1.84 $X2=3.39
+ $Y2=1.84
r101 22 48 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.225 $Y=2.22
+ $X2=3.225 $Y2=2.135
r102 22 24 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=3.225 $Y=2.22
+ $X2=3.225 $Y2=2.57
r103 21 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.135
+ $X2=0.28 $Y2=2.135
r104 20 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.06 $Y=2.135
+ $X2=3.225 $Y2=2.135
r105 20 21 170.604 $w=1.68e-07 $l=2.615e-06 $layer=LI1_cond $X=3.06 $Y=2.135
+ $X2=0.445 $Y2=2.135
r106 16 43 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.22
+ $X2=0.28 $Y2=2.135
r107 16 18 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=0.28 $Y=2.22
+ $X2=0.28 $Y2=2.815
r108 5 38 300 $w=1.7e-07 $l=5.57136e-07 $layer=licon1_PDIFF $count=2 $X=8.17
+ $Y=1.745 $X2=8.325 $Y2=2.23
r109 4 35 600 $w=1.7e-07 $l=1.35742e-06 $layer=licon1_PDIFF $count=1 $X=4.935
+ $Y=1.745 $X2=5.17 $Y2=2.99
r110 3 50 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=4.025
+ $Y=1.745 $X2=4.175 $Y2=1.92
r111 3 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.025
+ $Y=1.745 $X2=4.175 $Y2=2.72
r112 2 47 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.075
+ $Y=1.745 $X2=3.225 $Y2=1.89
r113 2 24 400 $w=1.7e-07 $l=8.9687e-07 $layer=licon1_PDIFF $count=1 $X=3.075
+ $Y=1.745 $X2=3.225 $Y2=2.57
r114 1 41 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r115 1 18 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_4%A_116_368# 1 2 3 4 15 19 21 23 24 25 26 29
+ 32 34
c61 25 0 6.57076e-20 $X=3.56 $Y=2.99
r62 27 29 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=3.725 $Y=2.905
+ $X2=3.725 $Y2=2.26
r63 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.56 $Y=2.99
+ $X2=3.725 $Y2=2.905
r64 25 26 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.56 $Y=2.99
+ $X2=2.885 $Y2=2.99
r65 24 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.76 $Y=2.905
+ $X2=2.885 $Y2=2.99
r66 23 36 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=2.56 $X2=2.76
+ $Y2=2.475
r67 23 24 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=2.76 $Y=2.56
+ $X2=2.76 $Y2=2.905
r68 22 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.895 $Y=2.475
+ $X2=1.77 $Y2=2.475
r69 21 36 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.635 $Y=2.475
+ $X2=2.76 $Y2=2.475
r70 21 22 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.635 $Y=2.475
+ $X2=1.895 $Y2=2.475
r71 17 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.77 $Y=2.56
+ $X2=1.77 $Y2=2.475
r72 17 19 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.77 $Y=2.56
+ $X2=1.77 $Y2=2.815
r73 16 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=2.475
+ $X2=0.78 $Y2=2.475
r74 15 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.645 $Y=2.475
+ $X2=1.77 $Y2=2.475
r75 15 16 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.645 $Y=2.475
+ $X2=0.945 $Y2=2.475
r76 4 29 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=3.525
+ $Y=1.745 $X2=3.725 $Y2=2.26
r77 3 36 600 $w=1.7e-07 $l=7.86432e-07 $layer=licon1_PDIFF $count=1 $X=2.57
+ $Y=1.84 $X2=2.72 $Y2=2.555
r78 2 34 600 $w=1.7e-07 $l=7.06028e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.73 $Y2=2.475
r79 2 19 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.73 $Y2=2.815
r80 1 32 300 $w=1.7e-07 $l=7.28166e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_4%VPWR 1 2 3 4 5 18 22 26 28 32 34 36 38 40
+ 45 50 58 64 67 70 73 77
c109 22 0 1.12408e-19 $X=2.25 $Y=2.815
r110 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r111 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r112 71 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r113 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r114 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r115 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r116 62 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r117 62 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r118 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r119 59 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.945 $Y=3.33
+ $X2=9.86 $Y2=3.33
r120 59 61 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=9.945 $Y=3.33
+ $X2=10.32 $Y2=3.33
r121 58 76 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=10.595 $Y=3.33
+ $X2=10.817 $Y2=3.33
r122 58 61 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.595 $Y=3.33
+ $X2=10.32 $Y2=3.33
r123 57 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r124 56 57 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r125 54 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r126 53 56 375.786 $w=1.68e-07 $l=5.76e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=8.4 $Y2=3.33
r127 53 54 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r128 51 67 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.435 $Y=3.33
+ $X2=2.25 $Y2=3.33
r129 51 53 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.435 $Y=3.33
+ $X2=2.64 $Y2=3.33
r130 50 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.79 $Y=3.33
+ $X2=8.955 $Y2=3.33
r131 50 56 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.79 $Y=3.33
+ $X2=8.4 $Y2=3.33
r132 49 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r133 49 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r134 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r135 46 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.28 $Y2=3.33
r136 46 48 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.68 $Y2=3.33
r137 45 67 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=2.25 $Y2=3.33
r138 45 48 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=1.68 $Y2=3.33
r139 43 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r140 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r141 40 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.28 $Y2=3.33
r142 40 42 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=0.72 $Y2=3.33
r143 38 57 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=8.4 $Y2=3.33
r144 38 54 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=2.64 $Y2=3.33
r145 34 76 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.76 $Y=3.245
+ $X2=10.817 $Y2=3.33
r146 34 36 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=10.76 $Y=3.245
+ $X2=10.76 $Y2=2.395
r147 30 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.86 $Y=3.245
+ $X2=9.86 $Y2=3.33
r148 30 32 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=9.86 $Y=3.245
+ $X2=9.86 $Y2=2.265
r149 29 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.12 $Y=3.33
+ $X2=8.955 $Y2=3.33
r150 28 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=3.33
+ $X2=9.86 $Y2=3.33
r151 28 29 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=9.775 $Y=3.33
+ $X2=9.12 $Y2=3.33
r152 24 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.955 $Y=3.245
+ $X2=8.955 $Y2=3.33
r153 24 26 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=8.955 $Y=3.245
+ $X2=8.955 $Y2=2.455
r154 20 67 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.25 $Y=3.245
+ $X2=2.25 $Y2=3.33
r155 20 22 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.25 $Y=3.245
+ $X2=2.25 $Y2=2.815
r156 16 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=3.245
+ $X2=1.28 $Y2=3.33
r157 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.28 $Y=3.245
+ $X2=1.28 $Y2=2.815
r158 5 36 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=10.61
+ $Y=2.12 $X2=10.76 $Y2=2.395
r159 4 32 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=9.71
+ $Y=2.12 $X2=9.86 $Y2=2.265
r160 3 26 300 $w=1.7e-07 $l=4.19375e-07 $layer=licon1_PDIFF $count=2 $X=8.765
+ $Y=2.12 $X2=8.955 $Y2=2.455
r161 2 22 600 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.84 $X2=2.25 $Y2=2.815
r162 1 18 600 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.84 $X2=1.28 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_4%A_897_349# 1 2 3 4 13 15 17 25 27
r40 25 32 2.80348 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=7.897 $Y=2.565
+ $X2=7.897 $Y2=2.65
r41 25 27 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=7.897 $Y=2.565
+ $X2=7.897 $Y2=2.23
r42 22 24 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=6.61 $Y=2.65
+ $X2=7.515 $Y2=2.65
r43 20 22 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=5.705 $Y=2.65
+ $X2=6.61 $Y2=2.65
r44 18 30 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.8 $Y=2.65
+ $X2=4.635 $Y2=2.65
r45 18 20 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=4.8 $Y=2.65
+ $X2=5.705 $Y2=2.65
r46 17 32 4.51856 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=7.76 $Y=2.65
+ $X2=7.897 $Y2=2.65
r47 17 24 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.76 $Y=2.65
+ $X2=7.515 $Y2=2.65
r48 13 30 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.635 $Y=2.565
+ $X2=4.635 $Y2=2.65
r49 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.635 $Y=2.565
+ $X2=4.635 $Y2=1.89
r50 4 32 600 $w=1.7e-07 $l=1.12962e-06 $layer=licon1_PDIFF $count=1 $X=7.365
+ $Y=1.745 $X2=7.87 $Y2=2.65
r51 4 27 600 $w=1.7e-07 $l=7.07071e-07 $layer=licon1_PDIFF $count=1 $X=7.365
+ $Y=1.745 $X2=7.87 $Y2=2.23
r52 4 24 600 $w=1.7e-07 $l=9.77126e-07 $layer=licon1_PDIFF $count=1 $X=7.365
+ $Y=1.745 $X2=7.515 $Y2=2.65
r53 3 22 600 $w=1.7e-07 $l=9.79439e-07 $layer=licon1_PDIFF $count=1 $X=6.455
+ $Y=1.745 $X2=6.61 $Y2=2.65
r54 2 20 600 $w=1.7e-07 $l=9.77126e-07 $layer=licon1_PDIFF $count=1 $X=5.555
+ $Y=1.745 $X2=5.705 $Y2=2.65
r55 1 30 400 $w=1.7e-07 $l=8.9687e-07 $layer=licon1_PDIFF $count=1 $X=4.485
+ $Y=1.745 $X2=4.635 $Y2=2.57
r56 1 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.485
+ $Y=1.745 $X2=4.635 $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_4%Y 1 2 3 4 5 6 7 8 9 10 33 35 36 39 41 45 47
+ 51 53 57 59 63 66 67 68 70 73 77 80 81 84 85 86 87 90 94 95 96 100
c183 95 0 1.65916e-19 $X=7.92 $Y=0.555
c184 77 0 1.59971e-19 $X=6.61 $Y=0.515
c185 36 0 3.21438e-20 $X=0.945 $Y=0.925
r186 96 100 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.87 $Y=0.97
+ $X2=7.87 $Y2=0.885
r187 96 100 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=7.87 $Y=0.862
+ $X2=7.87 $Y2=0.885
r188 95 96 12.1181 $w=3.28e-07 $l=3.47e-07 $layer=LI1_cond $X=7.87 $Y=0.515
+ $X2=7.87 $Y2=0.862
r189 82 94 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.775 $Y=0.97
+ $X2=6.61 $Y2=0.97
r190 81 96 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.705 $Y=0.97
+ $X2=7.87 $Y2=0.97
r191 81 82 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=7.705 $Y=0.97
+ $X2=6.775 $Y2=0.97
r192 80 90 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.53 $Y=1.3
+ $X2=6.53 $Y2=1.385
r193 79 94 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=6.53 $Y=1.055
+ $X2=6.61 $Y2=0.97
r194 79 80 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.53 $Y=1.055
+ $X2=6.53 $Y2=1.3
r195 75 94 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.61 $Y=0.885
+ $X2=6.61 $Y2=0.97
r196 75 77 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.61 $Y=0.885
+ $X2=6.61 $Y2=0.515
r197 71 93 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.32 $Y=1.89
+ $X2=6.155 $Y2=1.89
r198 71 73 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=6.32 $Y=1.89
+ $X2=7.065 $Y2=1.89
r199 70 93 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.155 $Y=1.725
+ $X2=6.155 $Y2=1.89
r200 69 90 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.155 $Y=1.385
+ $X2=6.53 $Y2=1.385
r201 69 70 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.155 $Y=1.47
+ $X2=6.155 $Y2=1.725
r202 67 69 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.99 $Y=1.385
+ $X2=6.155 $Y2=1.385
r203 67 68 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.99 $Y=1.385
+ $X2=5.775 $Y2=1.385
r204 66 68 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.65 $Y=1.3
+ $X2=5.775 $Y2=1.385
r205 65 88 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.65 $Y=1.085
+ $X2=5.65 $Y2=1
r206 65 66 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=5.65 $Y=1.085
+ $X2=5.65 $Y2=1.3
r207 61 88 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.65 $Y=0.915
+ $X2=5.65 $Y2=1
r208 61 63 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=5.65 $Y=0.915
+ $X2=5.65 $Y2=0.515
r209 60 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.845 $Y=1 $X2=4.68
+ $Y2=1
r210 59 88 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.525 $Y=1 $X2=5.65
+ $Y2=1
r211 59 60 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.525 $Y=1
+ $X2=4.845 $Y2=1
r212 55 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.68 $Y=0.915
+ $X2=4.68 $Y2=1
r213 55 57 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=4.68 $Y=0.915 $X2=4.68
+ $Y2=0.515
r214 54 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.845 $Y=1 $X2=3.72
+ $Y2=1
r215 53 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.515 $Y=1 $X2=4.68
+ $Y2=1
r216 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.515 $Y=1
+ $X2=3.845 $Y2=1
r217 49 86 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.915
+ $X2=3.72 $Y2=1
r218 49 51 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=3.72 $Y=0.915
+ $X2=3.72 $Y2=0.515
r219 48 85 7.02821 $w=1.7e-07 $l=1.42741e-07 $layer=LI1_cond $X=2.915 $Y=1
+ $X2=2.79 $Y2=0.962
r220 47 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.595 $Y=1 $X2=3.72
+ $Y2=1
r221 47 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.595 $Y=1
+ $X2=2.915 $Y2=1
r222 43 85 0.00168595 $w=2.5e-07 $l=1.22e-07 $layer=LI1_cond $X=2.79 $Y=0.84
+ $X2=2.79 $Y2=0.962
r223 43 45 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=2.79 $Y=0.84
+ $X2=2.79 $Y2=0.515
r224 42 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0.925
+ $X2=1.78 $Y2=0.925
r225 41 85 7.02821 $w=1.7e-07 $l=1.42302e-07 $layer=LI1_cond $X=2.665 $Y=0.925
+ $X2=2.79 $Y2=0.962
r226 41 42 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.665 $Y=0.925
+ $X2=1.945 $Y2=0.925
r227 37 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=0.84
+ $X2=1.78 $Y2=0.925
r228 37 39 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.78 $Y=0.84
+ $X2=1.78 $Y2=0.515
r229 35 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=0.925
+ $X2=1.78 $Y2=0.925
r230 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=0.925
+ $X2=0.945 $Y2=0.925
r231 31 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=0.84
+ $X2=0.945 $Y2=0.925
r232 31 33 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.78 $Y=0.84
+ $X2=0.78 $Y2=0.515
r233 10 73 600 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_PDIFF $count=1 $X=6.915
+ $Y=1.745 $X2=7.065 $Y2=1.93
r234 9 93 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.005
+ $Y=1.745 $X2=6.155 $Y2=1.89
r235 8 95 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.73
+ $Y=0.37 $X2=7.87 $Y2=0.515
r236 7 77 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.47
+ $Y=0.37 $X2=6.61 $Y2=0.515
r237 6 63 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.47
+ $Y=0.37 $X2=5.61 $Y2=0.515
r238 5 57 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=4.47
+ $Y=0.37 $X2=4.68 $Y2=0.515
r239 4 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.54
+ $Y=0.37 $X2=3.68 $Y2=0.515
r240 3 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.61
+ $Y=0.37 $X2=2.75 $Y2=0.515
r241 2 84 182 $w=1.7e-07 $l=6.40859e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.37 $X2=1.78 $Y2=0.925
r242 2 39 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.37 $X2=1.78 $Y2=0.515
r243 1 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NOR4BB_4%VGND 1 2 3 4 5 6 7 8 9 10 31 33 37 39 43 45
+ 49 51 55 57 61 63 67 69 73 77 81 83 85 90 95 105 106 112 115 118 121 124 127
+ 130 135 138
r165 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r166 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r167 131 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r168 130 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r169 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r170 128 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r171 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r172 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r173 122 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.04 $Y2=0
r174 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r175 119 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=4.08 $Y2=0
r176 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r177 116 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=3.12 $Y2=0
r178 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r179 113 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=2.16 $Y2=0
r180 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r181 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r182 106 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r183 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r184 103 138 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=10.495 $Y=0
+ $X2=10.295 $Y2=0
r185 103 105 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.495 $Y=0
+ $X2=10.8 $Y2=0
r186 102 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r187 101 102 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r188 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.84 $Y2=0
r189 99 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r190 98 101 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r191 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r192 96 135 11.8853 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=8.75 $Y=0
+ $X2=8.477 $Y2=0
r193 96 98 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=8.75 $Y=0 $X2=8.88
+ $Y2=0
r194 95 138 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=10.095 $Y=0
+ $X2=10.295 $Y2=0
r195 95 101 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.095 $Y=0
+ $X2=9.84 $Y2=0
r196 94 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r197 94 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r198 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r199 91 130 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=7.535 $Y=0
+ $X2=7.24 $Y2=0
r200 91 93 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.535 $Y=0
+ $X2=7.92 $Y2=0
r201 90 135 11.8853 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=8.205 $Y=0
+ $X2=8.477 $Y2=0
r202 90 93 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.205 $Y=0
+ $X2=7.92 $Y2=0
r203 89 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r204 89 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r205 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r206 86 109 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r207 86 88 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r208 85 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=1.28 $Y2=0
r209 85 88 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=0.72 $Y2=0
r210 83 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r211 83 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r212 79 138 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=10.295 $Y=0.085
+ $X2=10.295 $Y2=0
r213 79 81 12.3888 $w=3.98e-07 $l=4.3e-07 $layer=LI1_cond $X=10.295 $Y=0.085
+ $X2=10.295 $Y2=0.515
r214 75 135 2.29102 $w=5.45e-07 $l=8.5e-08 $layer=LI1_cond $X=8.477 $Y=0.085
+ $X2=8.477 $Y2=0
r215 75 77 9.43695 $w=5.43e-07 $l=4.3e-07 $layer=LI1_cond $X=8.477 $Y=0.085
+ $X2=8.477 $Y2=0.515
r216 71 130 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.24 $Y=0.085
+ $X2=7.24 $Y2=0
r217 71 73 8.71718 $w=5.88e-07 $l=4.3e-07 $layer=LI1_cond $X=7.24 $Y=0.085
+ $X2=7.24 $Y2=0.515
r218 70 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=0
+ $X2=6.11 $Y2=0
r219 69 130 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=6.945 $Y=0
+ $X2=7.24 $Y2=0
r220 69 70 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.945 $Y=0
+ $X2=6.275 $Y2=0
r221 65 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.11 $Y=0.085
+ $X2=6.11 $Y2=0
r222 65 67 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.11 $Y=0.085
+ $X2=6.11 $Y2=0.515
r223 64 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.345 $Y=0
+ $X2=5.18 $Y2=0
r224 63 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.945 $Y=0
+ $X2=6.11 $Y2=0
r225 63 64 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.945 $Y=0 $X2=5.345
+ $Y2=0
r226 59 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.18 $Y=0.085
+ $X2=5.18 $Y2=0
r227 59 61 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.18 $Y=0.085
+ $X2=5.18 $Y2=0.58
r228 58 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.345 $Y=0
+ $X2=4.18 $Y2=0
r229 57 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.015 $Y=0
+ $X2=5.18 $Y2=0
r230 57 58 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.015 $Y=0
+ $X2=4.345 $Y2=0
r231 53 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.18 $Y=0.085
+ $X2=4.18 $Y2=0
r232 53 55 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.18 $Y=0.085
+ $X2=4.18 $Y2=0.58
r233 52 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=0
+ $X2=3.25 $Y2=0
r234 51 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=0
+ $X2=4.18 $Y2=0
r235 51 52 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.015 $Y=0 $X2=3.415
+ $Y2=0
r236 47 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0
r237 47 49 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0.58
r238 46 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0
+ $X2=2.28 $Y2=0
r239 45 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=0
+ $X2=3.25 $Y2=0
r240 45 46 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=2.445
+ $Y2=0
r241 41 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0
r242 41 43 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0.55
r243 40 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0
+ $X2=1.28 $Y2=0
r244 39 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=0
+ $X2=2.28 $Y2=0
r245 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=0
+ $X2=1.445 $Y2=0
r246 35 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0
r247 35 37 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0.55
r248 31 109 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r249 31 33 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.515
r250 10 81 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=10.115
+ $Y=0.37 $X2=10.33 $Y2=0.515
r251 9 77 91 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=2 $X=8.185
+ $Y=0.37 $X2=8.665 $Y2=0.515
r252 8 73 91 $w=1.7e-07 $l=6.08194e-07 $layer=licon1_NDIFF $count=2 $X=6.9
+ $Y=0.37 $X2=7.44 $Y2=0.515
r253 7 67 91 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=2 $X=5.96
+ $Y=0.37 $X2=6.11 $Y2=0.515
r254 6 61 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=4.97
+ $Y=0.37 $X2=5.18 $Y2=0.58
r255 5 55 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.04
+ $Y=0.37 $X2=4.18 $Y2=0.58
r256 4 49 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=3.06
+ $Y=0.37 $X2=3.25 $Y2=0.58
r257 3 43 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.37 $X2=2.28 $Y2=0.55
r258 2 37 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.55
r259 1 33 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

