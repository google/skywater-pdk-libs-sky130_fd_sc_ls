* NGSPICE file created from sky130_fd_sc_ls__dfrbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR CLK a_319_392# VPB phighvt w=1e+06u l=150000u
+  ad=1.9859e+12p pd=1.77e+07u as=2.95e+11p ps=2.59e+06u
M1001 VGND CLK a_319_392# VNB nshort w=740000u l=150000u
+  ad=1.43248e+12p pd=1.25e+07u as=2.109e+11p ps=2.05e+06u
M1002 a_841_401# a_705_463# VGND VNB nshort w=640000u l=150000u
+  ad=3.222e+11p pd=2.44e+06u as=0p ps=0u
M1003 VPWR a_1224_74# a_2026_424# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1004 a_1224_74# a_500_392# a_841_401# VNB nshort w=640000u l=150000u
+  ad=4.33e+11p pd=3.08e+06u as=0p ps=0u
M1005 Q a_2026_424# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 VPWR a_841_401# a_796_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 a_125_78# D a_38_78# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.436e+11p ps=2.84e+06u
M1008 VGND a_1224_74# a_2026_424# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1009 Q_N a_1224_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1010 a_832_119# a_500_392# a_705_463# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.47e+11p ps=1.54e+06u
M1011 Q_N a_1224_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.888e+11p pd=3.47e+06u as=0p ps=0u
M1012 a_1224_74# a_319_392# a_841_401# VPB phighvt w=1e+06u l=150000u
+  ad=3.877e+11p pd=3.2e+06u as=3e+11p ps=2.6e+06u
M1013 a_705_463# a_319_392# a_38_78# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1482_48# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1015 VGND RESET_B a_910_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1016 VPWR a_1482_48# a_1465_471# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1017 a_841_401# a_705_463# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1465_471# a_500_392# a_1224_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_705_463# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.457e+11p pd=2.85e+06u as=0p ps=0u
M1020 VPWR a_1224_74# a_1482_48# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_38_78# D VPWR VPB phighvt w=420000u l=150000u
+  ad=2.478e+11p pd=2.86e+06u as=0p ps=0u
M1022 VPWR RESET_B a_38_78# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_705_463# a_500_392# a_38_78# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_1482_48# a_1434_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 a_796_463# a_319_392# a_705_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1624_74# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1027 a_1482_48# a_1224_74# a_1624_74# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1028 VGND RESET_B a_125_78# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_500_392# a_319_392# VGND VNB nshort w=740000u l=150000u
+  ad=2.0885e+11p pd=2.07e+06u as=0p ps=0u
M1030 a_500_392# a_319_392# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1031 Q a_2026_424# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1032 a_1434_74# a_319_392# a_1224_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_910_119# a_841_401# a_832_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

