* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 VPWR a_2087_410# a_2042_508# VPB phighvt w=420000u l=150000u
+  ad=2.13575e+12p pd=1.79e+07u as=1.092e+11p ps=1.36e+06u
M1001 VGND a_2087_410# a_2073_74# VNB nshort w=420000u l=150000u
+  ad=1.77155e+12p pd=1.431e+07u as=1.05e+11p ps=1.34e+06u
M1002 a_284_464# D a_206_464# VPB phighvt w=640000u l=150000u
+  ad=8.151e+11p pd=6.15e+06u as=1.536e+11p ps=1.76e+06u
M1003 a_538_81# SCE a_284_464# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.549e+11p ps=3.37e+06u
M1004 a_1251_463# a_854_74# a_284_464# VPB phighvt w=420000u l=150000u
+  ad=2.499e+11p pd=2.87e+06u as=0p ps=0u
M1005 a_2087_410# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1006 Q a_2492_424# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1007 a_2265_74# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1008 a_2087_410# a_1827_144# a_2265_74# VNB nshort w=420000u l=150000u
+  ad=2.1e+11p pd=1.84e+06u as=0p ps=0u
M1009 a_1827_144# a_1049_347# a_1402_308# VPB phighvt w=1e+06u l=150000u
+  ad=3.128e+11p pd=2.73e+06u as=7.85e+11p ps=3.57e+06u
M1010 a_1049_347# a_854_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1011 VGND RESET_B a_1489_123# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1012 a_854_74# CLK_N VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1013 a_1251_463# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1411_123# a_854_74# a_1251_463# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.289e+11p ps=1.93e+06u
M1015 Q a_2492_424# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1016 VPWR SCD a_471_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1017 VPWR a_1827_144# a_2087_410# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1341_463# a_1049_347# a_1251_463# VPB phighvt w=420000u l=150000u
+  ad=1.281e+11p pd=1.45e+06u as=0p ps=0u
M1019 a_324_81# a_27_88# a_239_81# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.373e+11p ps=2.81e+06u
M1020 a_1402_308# a_1251_463# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_2042_508# a_854_74# a_1827_144# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_284_464# D a_324_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1251_463# a_1049_347# a_284_464# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR CLK_N a_854_74# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=3.35e+11p ps=2.67e+06u
M1025 VPWR a_1402_308# a_1341_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND RESET_B a_239_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_1827_144# a_2492_424# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1028 a_1049_347# a_854_74# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.122e+11p pd=2.67e+06u as=0p ps=0u
M1029 a_1489_123# a_1402_308# a_1411_123# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR SCE a_27_88# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1031 a_206_464# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_2073_74# a_1049_347# a_1827_144# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=6.2565e+11p ps=4.26e+06u
M1033 VGND a_1827_144# a_2492_424# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1034 a_239_81# SCD a_538_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_471_464# a_27_88# a_284_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1402_308# a_1251_463# VGND VNB nshort w=640000u l=150000u
+  ad=3.584e+11p pd=2.4e+06u as=0p ps=0u
M1037 VGND SCE a_27_88# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1038 a_1827_144# a_854_74# a_1402_308# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_284_464# RESET_B VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
