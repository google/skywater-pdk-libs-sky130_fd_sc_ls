* File: sky130_fd_sc_ls__o21a_1.spice
* Created: Fri Aug 28 13:44:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o21a_1.pex.spice"
.subckt sky130_fd_sc_ls__o21a_1  VNB VPB B1 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_83_244#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_320_74#_M1002_d N_B1_M1002_g N_A_83_244#_M1002_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_320_74#_M1002_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_A_320_74#_M1001_d N_A1_M1001_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_A_83_244#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.382657 AS=0.3304 PD=2.01714 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1003 N_A_83_244#_M1003_d N_B1_M1003_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.155491 AS=0.286993 PD=1.23717 PS=1.51286 NRD=2.3443 NRS=43.3794 M=1 R=5.6
+ SA=75001 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1004 A_376_387# N_A2_M1004_g N_A_83_244#_M1003_d VPB PHIGHVT L=0.15 W=1
+ AD=0.21 AS=0.185109 PD=1.42 PS=1.47283 NRD=30.5153 NRS=12.7853 M=1 R=6.66667
+ SA=75001.3 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g A_376_387# VPB PHIGHVT L=0.15 W=1 AD=0.295
+ AS=0.21 PD=2.59 PS=1.42 NRD=1.9503 NRS=30.5153 M=1 R=6.66667 SA=75001.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ls__o21a_1.pxi.spice"
*
.ends
*
*
