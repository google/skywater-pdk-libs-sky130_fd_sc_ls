* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
X0 a_1273_392# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_1273_392# B a_1060_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_193_277# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 a_193_277# a_27_94# a_791_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_193_277# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 X a_193_277# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 VPWR A a_1273_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_193_277# a_678_368# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 a_791_392# a_678_368# a_1060_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_27_94# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 VPWR a_193_277# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 VGND C_N a_678_368# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_27_94# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_1060_392# a_678_368# a_791_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_1060_392# B a_1273_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_193_277# A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 VGND a_193_277# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 VGND B a_193_277# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 VPWR C_N a_678_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_791_392# a_27_94# a_193_277# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VGND a_27_94# a_193_277# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 VPWR a_193_277# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X22 X a_193_277# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X23 X a_193_277# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
