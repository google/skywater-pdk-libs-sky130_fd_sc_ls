* File: sky130_fd_sc_ls__mux2i_1.pxi.spice
* Created: Wed Sep  2 11:10:32 2020
* 
x_PM_SKY130_FD_SC_LS__MUX2I_1%S N_S_M1007_g N_S_c_76_n N_S_M1006_g N_S_c_69_n
+ N_S_c_70_n N_S_c_78_n N_S_M1002_g N_S_c_71_n N_S_M1009_g N_S_c_72_n N_S_c_79_n
+ N_S_c_73_n S S N_S_c_75_n PM_SKY130_FD_SC_LS__MUX2I_1%S
x_PM_SKY130_FD_SC_LS__MUX2I_1%A_114_74# N_A_114_74#_M1007_d N_A_114_74#_M1006_d
+ N_A_114_74#_c_132_n N_A_114_74#_M1005_g N_A_114_74#_M1000_g
+ N_A_114_74#_c_134_n N_A_114_74#_c_135_n N_A_114_74#_c_136_n
+ N_A_114_74#_c_141_n N_A_114_74#_c_137_n N_A_114_74#_c_138_n
+ N_A_114_74#_c_139_n PM_SKY130_FD_SC_LS__MUX2I_1%A_114_74#
x_PM_SKY130_FD_SC_LS__MUX2I_1%A0 N_A0_M1001_g N_A0_c_206_n N_A0_M1004_g A0
+ N_A0_c_204_n N_A0_c_205_n PM_SKY130_FD_SC_LS__MUX2I_1%A0
x_PM_SKY130_FD_SC_LS__MUX2I_1%A1 N_A1_c_237_n N_A1_M1003_g N_A1_c_238_n
+ N_A1_M1008_g A1 PM_SKY130_FD_SC_LS__MUX2I_1%A1
x_PM_SKY130_FD_SC_LS__MUX2I_1%VPWR N_VPWR_M1006_s N_VPWR_M1002_d N_VPWR_c_258_n
+ N_VPWR_c_259_n N_VPWR_c_260_n VPWR N_VPWR_c_261_n N_VPWR_c_262_n
+ N_VPWR_c_257_n N_VPWR_c_264_n PM_SKY130_FD_SC_LS__MUX2I_1%VPWR
x_PM_SKY130_FD_SC_LS__MUX2I_1%A_223_368# N_A_223_368#_M1002_s
+ N_A_223_368#_M1004_s N_A_223_368#_c_294_n N_A_223_368#_c_295_n
+ N_A_223_368#_c_296_n N_A_223_368#_c_297_n
+ PM_SKY130_FD_SC_LS__MUX2I_1%A_223_368#
x_PM_SKY130_FD_SC_LS__MUX2I_1%A_399_368# N_A_399_368#_M1005_d
+ N_A_399_368#_M1008_d N_A_399_368#_c_324_n N_A_399_368#_c_325_n
+ N_A_399_368#_c_326_n N_A_399_368#_c_327_n
+ PM_SKY130_FD_SC_LS__MUX2I_1%A_399_368#
x_PM_SKY130_FD_SC_LS__MUX2I_1%Y N_Y_M1001_d N_Y_M1004_d N_Y_c_368_p N_Y_c_349_n
+ N_Y_c_351_n Y PM_SKY130_FD_SC_LS__MUX2I_1%Y
x_PM_SKY130_FD_SC_LS__MUX2I_1%VGND N_VGND_M1007_s N_VGND_M1009_d N_VGND_c_370_n
+ N_VGND_c_371_n N_VGND_c_372_n VGND N_VGND_c_373_n N_VGND_c_374_n
+ N_VGND_c_375_n N_VGND_c_376_n PM_SKY130_FD_SC_LS__MUX2I_1%VGND
x_PM_SKY130_FD_SC_LS__MUX2I_1%A_225_74# N_A_225_74#_M1009_s N_A_225_74#_M1003_d
+ N_A_225_74#_c_406_n N_A_225_74#_c_407_n N_A_225_74#_c_408_n
+ N_A_225_74#_c_417_n N_A_225_74#_c_409_n N_A_225_74#_c_410_n
+ N_A_225_74#_c_411_n PM_SKY130_FD_SC_LS__MUX2I_1%A_225_74#
cc_1 VNB N_S_M1007_g 0.0378713f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_2 VNB N_S_c_69_n 0.0500851f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.26
cc_3 VNB N_S_c_70_n 0.020162f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.675
cc_4 VNB N_S_c_71_n 0.0203248f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.185
cc_5 VNB N_S_c_72_n 0.0155613f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.26
cc_6 VNB N_S_c_73_n 0.00664804f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.26
cc_7 VNB S 0.0234095f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_S_c_75_n 0.0290861f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.35
cc_9 VNB N_A_114_74#_c_132_n 0.0269713f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.54
cc_10 VNB N_A_114_74#_M1000_g 0.0251947f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.765
cc_11 VNB N_A_114_74#_c_134_n 0.00541105f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.74
cc_12 VNB N_A_114_74#_c_135_n 0.0201137f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.68
cc_13 VNB N_A_114_74#_c_136_n 0.00490111f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_14 VNB N_A_114_74#_c_137_n 0.00341769f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.35
cc_15 VNB N_A_114_74#_c_138_n 0.00106462f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.295
cc_16 VNB N_A_114_74#_c_139_n 0.00166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A0_M1001_g 0.0286315f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_18 VNB N_A0_c_204_n 0.0456805f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.765
cc_19 VNB N_A0_c_205_n 0.00549587f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.4
cc_20 VNB N_A1_c_237_n 0.0257716f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_21 VNB N_A1_c_238_n 0.0728652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB A1 0.00924341f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.54
cc_23 VNB N_VPWR_c_257_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.35
cc_24 VNB N_Y_c_349_n 0.0122596f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.26
cc_25 VNB N_VGND_c_370_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.54
cc_26 VNB N_VGND_c_371_n 0.0325289f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.26
cc_27 VNB N_VGND_c_372_n 0.00969314f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.4
cc_28 VNB N_VGND_c_373_n 0.034428f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.74
cc_29 VNB N_VGND_c_374_n 0.0504776f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.35
cc_30 VNB N_VGND_c_375_n 0.240757f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.35
cc_31 VNB N_VGND_c_376_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_225_74#_c_406_n 0.00874347f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.26
cc_33 VNB N_A_225_74#_c_407_n 0.0100806f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.675
cc_34 VNB N_A_225_74#_c_408_n 0.00386611f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.765
cc_35 VNB N_A_225_74#_c_409_n 0.0070932f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.185
cc_36 VNB N_A_225_74#_c_410_n 0.00124385f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.74
cc_37 VNB N_A_225_74#_c_411_n 0.0279156f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.68
cc_38 VPB N_S_c_76_n 0.0215428f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.045
cc_39 VPB N_S_c_70_n 9.12936e-19 $X=-0.19 $Y=1.66 $X2=1.47 $Y2=1.675
cc_40 VPB N_S_c_78_n 0.0258098f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=1.765
cc_41 VPB N_S_c_79_n 0.0398526f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.68
cc_42 VPB S 0.0120179f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_43 VPB N_S_c_75_n 0.00170579f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.35
cc_44 VPB N_A_114_74#_c_132_n 0.0300925f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.54
cc_45 VPB N_A_114_74#_c_141_n 0.0165755f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.35
cc_46 VPB N_A_114_74#_c_137_n 0.0100316f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.35
cc_47 VPB N_A_114_74#_c_139_n 0.00163415f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A0_c_206_n 0.0188216f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.045
cc_49 VPB N_A0_c_204_n 0.0158841f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=1.765
cc_50 VPB N_A0_c_205_n 0.00433843f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.4
cc_51 VPB N_A1_c_238_n 0.0289127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_258_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.54
cc_53 VPB N_VPWR_c_259_n 0.0472879f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.26
cc_54 VPB N_VPWR_c_260_n 0.00396467f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.4
cc_55 VPB N_VPWR_c_261_n 0.0326305f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.74
cc_56 VPB N_VPWR_c_262_n 0.0489572f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.35
cc_57 VPB N_VPWR_c_257_n 0.0754942f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.35
cc_58 VPB N_VPWR_c_264_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_223_368#_c_294_n 0.00524382f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.54
cc_60 VPB N_A_223_368#_c_295_n 0.00993695f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.26
cc_61 VPB N_A_223_368#_c_296_n 0.0135882f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=1.675
cc_62 VPB N_A_223_368#_c_297_n 0.00743377f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.335
cc_63 VPB N_A_399_368#_c_324_n 0.0069146f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.26
cc_64 VPB N_A_399_368#_c_325_n 0.0244674f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=1.675
cc_65 VPB N_A_399_368#_c_326_n 0.0036816f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=1.765
cc_66 VPB N_A_399_368#_c_327_n 0.0443277f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=1.185
cc_67 VPB N_Y_c_349_n 0.00400788f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.26
cc_68 N_S_c_70_n N_A_114_74#_c_132_n 0.0183509f $X=1.47 $Y=1.675 $X2=0 $Y2=0
cc_69 N_S_c_78_n N_A_114_74#_c_132_n 0.031233f $X=1.47 $Y=1.765 $X2=0 $Y2=0
cc_70 N_S_c_71_n N_A_114_74#_M1000_g 0.026721f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_71 N_S_M1007_g N_A_114_74#_c_134_n 0.00968387f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_72 N_S_c_69_n N_A_114_74#_c_134_n 0.0189538f $X=1.38 $Y=1.26 $X2=0 $Y2=0
cc_73 N_S_c_70_n N_A_114_74#_c_134_n 3.49755e-19 $X=1.47 $Y=1.675 $X2=0 $Y2=0
cc_74 S N_A_114_74#_c_134_n 0.0123511f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_75 N_S_c_75_n N_A_114_74#_c_134_n 3.2525e-19 $X=0.385 $Y=1.35 $X2=0 $Y2=0
cc_76 N_S_c_69_n N_A_114_74#_c_135_n 0.0129614f $X=1.38 $Y=1.26 $X2=0 $Y2=0
cc_77 N_S_c_70_n N_A_114_74#_c_135_n 0.014938f $X=1.47 $Y=1.675 $X2=0 $Y2=0
cc_78 N_S_M1007_g N_A_114_74#_c_136_n 0.009213f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_79 N_S_c_69_n N_A_114_74#_c_136_n 0.0020895f $X=1.38 $Y=1.26 $X2=0 $Y2=0
cc_80 N_S_c_71_n N_A_114_74#_c_136_n 0.0015289f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_81 N_S_c_76_n N_A_114_74#_c_141_n 0.0143683f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_82 N_S_c_79_n N_A_114_74#_c_141_n 7.14971e-19 $X=0.395 $Y=1.68 $X2=0 $Y2=0
cc_83 N_S_c_76_n N_A_114_74#_c_137_n 0.00188924f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_84 N_S_c_70_n N_A_114_74#_c_137_n 0.00609573f $X=1.47 $Y=1.675 $X2=0 $Y2=0
cc_85 N_S_c_78_n N_A_114_74#_c_137_n 0.00148469f $X=1.47 $Y=1.765 $X2=0 $Y2=0
cc_86 N_S_c_79_n N_A_114_74#_c_137_n 0.00689804f $X=0.395 $Y=1.68 $X2=0 $Y2=0
cc_87 S N_A_114_74#_c_137_n 0.0255963f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_88 N_S_c_75_n N_A_114_74#_c_137_n 0.00775954f $X=0.385 $Y=1.35 $X2=0 $Y2=0
cc_89 S N_A_114_74#_c_138_n 0.0145892f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_90 N_S_c_75_n N_A_114_74#_c_138_n 0.00410432f $X=0.385 $Y=1.35 $X2=0 $Y2=0
cc_91 N_S_c_70_n N_A_114_74#_c_139_n 0.00116727f $X=1.47 $Y=1.675 $X2=0 $Y2=0
cc_92 N_S_c_76_n N_VPWR_c_259_n 0.0112103f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_93 N_S_c_79_n N_VPWR_c_259_n 0.00100521f $X=0.395 $Y=1.68 $X2=0 $Y2=0
cc_94 S N_VPWR_c_259_n 0.0158723f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_95 N_S_c_78_n N_VPWR_c_260_n 0.0140627f $X=1.47 $Y=1.765 $X2=0 $Y2=0
cc_96 N_S_c_76_n N_VPWR_c_261_n 0.00445602f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_97 N_S_c_78_n N_VPWR_c_261_n 0.00413917f $X=1.47 $Y=1.765 $X2=0 $Y2=0
cc_98 N_S_c_76_n N_VPWR_c_257_n 0.00865852f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_99 N_S_c_78_n N_VPWR_c_257_n 0.00822528f $X=1.47 $Y=1.765 $X2=0 $Y2=0
cc_100 N_S_c_78_n N_A_223_368#_c_294_n 0.00314968f $X=1.47 $Y=1.765 $X2=0 $Y2=0
cc_101 N_S_c_76_n N_A_223_368#_c_295_n 0.00163285f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_102 N_S_c_78_n N_A_223_368#_c_295_n 0.00729586f $X=1.47 $Y=1.765 $X2=0 $Y2=0
cc_103 N_S_c_78_n N_A_223_368#_c_296_n 0.0139903f $X=1.47 $Y=1.765 $X2=0 $Y2=0
cc_104 N_S_M1007_g N_VGND_c_371_n 0.00800579f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_105 N_S_c_72_n N_VGND_c_371_n 0.0010506f $X=0.395 $Y=1.26 $X2=0 $Y2=0
cc_106 S N_VGND_c_371_n 0.015437f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_107 N_S_c_71_n N_VGND_c_372_n 0.00622602f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_108 N_S_M1007_g N_VGND_c_373_n 0.0043544f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_109 N_S_c_71_n N_VGND_c_373_n 0.00434272f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_110 N_S_M1007_g N_VGND_c_375_n 0.00830065f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_111 N_S_c_71_n N_VGND_c_375_n 0.00826311f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_112 N_S_M1007_g N_A_225_74#_c_406_n 0.0024493f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_113 N_S_c_71_n N_A_225_74#_c_406_n 0.0103339f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_114 N_S_c_71_n N_A_225_74#_c_407_n 0.0117984f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_115 N_S_c_69_n N_A_225_74#_c_408_n 0.00554277f $X=1.38 $Y=1.26 $X2=0 $Y2=0
cc_116 N_S_c_71_n N_A_225_74#_c_408_n 0.00214722f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_117 N_S_c_71_n N_A_225_74#_c_417_n 5.97863e-19 $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_118 N_A_114_74#_M1000_g N_A0_M1001_g 0.0329672f $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_119 N_A_114_74#_c_132_n N_A0_c_204_n 0.0378784f $X=1.92 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A_114_74#_c_139_n N_A0_c_204_n 8.89634e-19 $X=1.965 $Y=1.435 $X2=0
+ $Y2=0
cc_121 N_A_114_74#_c_132_n N_A0_c_205_n 0.00436678f $X=1.92 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A_114_74#_c_139_n N_A0_c_205_n 0.013347f $X=1.965 $Y=1.435 $X2=0 $Y2=0
cc_123 N_A_114_74#_c_141_n N_VPWR_c_259_n 0.0590978f $X=0.72 $Y=2.265 $X2=0
+ $Y2=0
cc_124 N_A_114_74#_c_132_n N_VPWR_c_260_n 0.0110386f $X=1.92 $Y=1.765 $X2=0
+ $Y2=0
cc_125 N_A_114_74#_c_141_n N_VPWR_c_261_n 0.0148169f $X=0.72 $Y=2.265 $X2=0
+ $Y2=0
cc_126 N_A_114_74#_c_132_n N_VPWR_c_262_n 0.00413917f $X=1.92 $Y=1.765 $X2=0
+ $Y2=0
cc_127 N_A_114_74#_c_132_n N_VPWR_c_257_n 0.00822528f $X=1.92 $Y=1.765 $X2=0
+ $Y2=0
cc_128 N_A_114_74#_c_141_n N_VPWR_c_257_n 0.0122313f $X=0.72 $Y=2.265 $X2=0
+ $Y2=0
cc_129 N_A_114_74#_c_135_n N_A_223_368#_c_294_n 0.0142143f $X=1.8 $Y=1.435 $X2=0
+ $Y2=0
cc_130 N_A_114_74#_c_137_n N_A_223_368#_c_294_n 0.0226777f $X=0.722 $Y=2.1 $X2=0
+ $Y2=0
cc_131 N_A_114_74#_c_141_n N_A_223_368#_c_295_n 0.0648591f $X=0.72 $Y=2.265
+ $X2=0 $Y2=0
cc_132 N_A_114_74#_c_132_n N_A_223_368#_c_296_n 0.0179664f $X=1.92 $Y=1.765
+ $X2=0 $Y2=0
cc_133 N_A_114_74#_c_135_n N_A_223_368#_c_296_n 0.0145543f $X=1.8 $Y=1.435 $X2=0
+ $Y2=0
cc_134 N_A_114_74#_c_139_n N_A_223_368#_c_296_n 0.014055f $X=1.965 $Y=1.435
+ $X2=0 $Y2=0
cc_135 N_A_114_74#_c_132_n N_A_223_368#_c_297_n 0.00473866f $X=1.92 $Y=1.765
+ $X2=0 $Y2=0
cc_136 N_A_114_74#_c_132_n N_A_399_368#_c_326_n 0.00292669f $X=1.92 $Y=1.765
+ $X2=0 $Y2=0
cc_137 N_A_114_74#_M1000_g N_Y_c_351_n 2.75206e-19 $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A_114_74#_M1000_g N_VGND_c_372_n 0.00622568f $X=2.055 $Y=0.74 $X2=0
+ $Y2=0
cc_139 N_A_114_74#_c_136_n N_VGND_c_373_n 0.0111177f $X=0.71 $Y=0.645 $X2=0
+ $Y2=0
cc_140 N_A_114_74#_M1000_g N_VGND_c_374_n 0.00433139f $X=2.055 $Y=0.74 $X2=0
+ $Y2=0
cc_141 N_A_114_74#_M1000_g N_VGND_c_375_n 0.00817354f $X=2.055 $Y=0.74 $X2=0
+ $Y2=0
cc_142 N_A_114_74#_c_136_n N_VGND_c_375_n 0.0120515f $X=0.71 $Y=0.645 $X2=0
+ $Y2=0
cc_143 N_A_114_74#_M1000_g N_A_225_74#_c_406_n 6.28869e-19 $X=2.055 $Y=0.74
+ $X2=0 $Y2=0
cc_144 N_A_114_74#_c_136_n N_A_225_74#_c_406_n 0.0424364f $X=0.71 $Y=0.645 $X2=0
+ $Y2=0
cc_145 N_A_114_74#_c_132_n N_A_225_74#_c_407_n 0.00124873f $X=1.92 $Y=1.765
+ $X2=0 $Y2=0
cc_146 N_A_114_74#_M1000_g N_A_225_74#_c_407_n 0.0136151f $X=2.055 $Y=0.74 $X2=0
+ $Y2=0
cc_147 N_A_114_74#_c_135_n N_A_225_74#_c_407_n 0.0265109f $X=1.8 $Y=1.435 $X2=0
+ $Y2=0
cc_148 N_A_114_74#_c_139_n N_A_225_74#_c_407_n 0.0243844f $X=1.965 $Y=1.435
+ $X2=0 $Y2=0
cc_149 N_A_114_74#_c_134_n N_A_225_74#_c_408_n 0.0121698f $X=0.805 $Y=1.35 $X2=0
+ $Y2=0
cc_150 N_A_114_74#_c_135_n N_A_225_74#_c_408_n 0.0275396f $X=1.8 $Y=1.435 $X2=0
+ $Y2=0
cc_151 N_A_114_74#_M1000_g N_A_225_74#_c_417_n 0.00985062f $X=2.055 $Y=0.74
+ $X2=0 $Y2=0
cc_152 N_A_114_74#_M1000_g N_A_225_74#_c_410_n 0.00375375f $X=2.055 $Y=0.74
+ $X2=0 $Y2=0
cc_153 N_A0_M1001_g N_A1_c_237_n 0.0101019f $X=2.445 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_154 N_A0_c_206_n N_A1_c_238_n 0.0222047f $X=2.895 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A0_c_204_n N_A1_c_238_n 0.0163629f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_156 N_A0_c_206_n N_VPWR_c_262_n 0.00278271f $X=2.895 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A0_c_206_n N_VPWR_c_257_n 0.00358708f $X=2.895 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A0_c_204_n N_A_223_368#_c_296_n 0.00415885f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_159 N_A0_c_206_n N_A_223_368#_c_297_n 0.00967983f $X=2.895 $Y=1.765 $X2=0
+ $Y2=0
cc_160 N_A0_c_204_n N_A_223_368#_c_297_n 0.00231888f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_161 N_A0_c_205_n N_A_223_368#_c_297_n 0.0247498f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_162 N_A0_c_206_n N_A_399_368#_c_324_n 0.00469671f $X=2.895 $Y=1.765 $X2=0
+ $Y2=0
cc_163 N_A0_c_206_n N_A_399_368#_c_325_n 0.0154499f $X=2.895 $Y=1.765 $X2=0
+ $Y2=0
cc_164 N_A0_c_206_n N_A_399_368#_c_327_n 9.91116e-19 $X=2.895 $Y=1.765 $X2=0
+ $Y2=0
cc_165 N_A0_M1001_g N_Y_c_349_n 0.00502765f $X=2.445 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A0_c_204_n N_Y_c_349_n 0.010378f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_167 N_A0_c_205_n N_Y_c_349_n 0.0326257f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_168 N_A0_M1001_g N_Y_c_351_n 0.00510039f $X=2.445 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A0_c_204_n N_Y_c_351_n 0.00594294f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_170 N_A0_c_205_n N_Y_c_351_n 0.015419f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_171 N_A0_M1001_g N_VGND_c_374_n 0.00291649f $X=2.445 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A0_M1001_g N_VGND_c_375_n 0.00361693f $X=2.445 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A0_M1001_g N_A_225_74#_c_407_n 0.00451515f $X=2.445 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A0_M1001_g N_A_225_74#_c_417_n 0.00611057f $X=2.445 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A0_M1001_g N_A_225_74#_c_409_n 0.0149352f $X=2.445 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A1_c_238_n N_VPWR_c_262_n 0.00278257f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A1_c_238_n N_VPWR_c_257_n 0.00357366f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A1_c_238_n N_A_399_368#_c_325_n 0.0134197f $X=3.345 $Y=1.765 $X2=0
+ $Y2=0
cc_179 N_A1_c_238_n N_A_399_368#_c_327_n 0.0161774f $X=3.345 $Y=1.765 $X2=0
+ $Y2=0
cc_180 A1 N_A_399_368#_c_327_n 0.0191396f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_181 N_A1_c_237_n N_Y_c_349_n 0.00708472f $X=3.3 $Y=1.22 $X2=0 $Y2=0
cc_182 N_A1_c_238_n N_Y_c_349_n 0.0079021f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_183 A1 N_Y_c_349_n 0.0282043f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_184 N_A1_c_237_n N_VGND_c_374_n 0.00291649f $X=3.3 $Y=1.22 $X2=0 $Y2=0
cc_185 N_A1_c_237_n N_VGND_c_375_n 0.00365785f $X=3.3 $Y=1.22 $X2=0 $Y2=0
cc_186 N_A1_c_237_n N_A_225_74#_c_409_n 0.0142787f $X=3.3 $Y=1.22 $X2=0 $Y2=0
cc_187 N_A1_c_238_n N_A_225_74#_c_411_n 0.00189227f $X=3.345 $Y=1.765 $X2=0
+ $Y2=0
cc_188 A1 N_A_225_74#_c_411_n 0.0232175f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_189 N_VPWR_c_260_n N_A_223_368#_c_295_n 0.0462948f $X=1.695 $Y=2.455 $X2=0
+ $Y2=0
cc_190 N_VPWR_c_261_n N_A_223_368#_c_295_n 0.011066f $X=1.53 $Y=3.33 $X2=0 $Y2=0
cc_191 N_VPWR_c_257_n N_A_223_368#_c_295_n 0.00915947f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_192 N_VPWR_M1002_d N_A_223_368#_c_296_n 0.00507752f $X=1.545 $Y=1.84 $X2=0
+ $Y2=0
cc_193 N_VPWR_c_260_n N_A_223_368#_c_296_n 0.0171814f $X=1.695 $Y=2.455 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_260_n N_A_399_368#_c_324_n 0.0412023f $X=1.695 $Y=2.455 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_262_n N_A_399_368#_c_325_n 0.0932569f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_196 N_VPWR_c_257_n N_A_399_368#_c_325_n 0.0526262f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_197 N_VPWR_c_260_n N_A_399_368#_c_326_n 0.0125885f $X=1.695 $Y=2.455 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_262_n N_A_399_368#_c_326_n 0.0179217f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_199 N_VPWR_c_257_n N_A_399_368#_c_326_n 0.00971942f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_200 N_A_223_368#_c_296_n N_A_399_368#_M1005_d 0.00963455f $X=2.505 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_201 N_A_223_368#_c_296_n N_A_399_368#_c_324_n 0.0202979f $X=2.505 $Y=2.035
+ $X2=0 $Y2=0
cc_202 N_A_223_368#_c_297_n N_A_399_368#_c_324_n 0.0329564f $X=2.67 $Y=2.115
+ $X2=0 $Y2=0
cc_203 N_A_223_368#_M1004_s N_A_399_368#_c_325_n 0.00266942f $X=2.54 $Y=1.84
+ $X2=0 $Y2=0
cc_204 N_A_223_368#_c_297_n N_A_399_368#_c_325_n 0.0206198f $X=2.67 $Y=2.115
+ $X2=0 $Y2=0
cc_205 N_A_223_368#_c_297_n N_Y_c_349_n 0.0522275f $X=2.67 $Y=2.115 $X2=0 $Y2=0
cc_206 N_A_399_368#_c_325_n N_Y_M1004_d 0.00222494f $X=3.405 $Y=2.99 $X2=0 $Y2=0
cc_207 N_A_399_368#_c_325_n N_Y_c_349_n 0.013472f $X=3.405 $Y=2.99 $X2=0 $Y2=0
cc_208 N_A_399_368#_c_327_n N_Y_c_349_n 0.0334931f $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_209 N_Y_c_351_n N_A_225_74#_c_407_n 0.00171692f $X=3.035 $Y=0.87 $X2=0 $Y2=0
cc_210 N_Y_c_351_n N_A_225_74#_c_417_n 0.0195323f $X=3.035 $Y=0.87 $X2=0 $Y2=0
cc_211 N_Y_M1001_d N_A_225_74#_c_409_n 0.00935673f $X=2.52 $Y=0.37 $X2=0 $Y2=0
cc_212 N_Y_c_368_p N_A_225_74#_c_409_n 0.00960383f $X=3.13 $Y=1.035 $X2=0 $Y2=0
cc_213 N_Y_c_351_n N_A_225_74#_c_409_n 0.032664f $X=3.035 $Y=0.87 $X2=0 $Y2=0
cc_214 N_VGND_c_372_n N_A_225_74#_c_406_n 0.0191765f $X=1.77 $Y=0.675 $X2=0
+ $Y2=0
cc_215 N_VGND_c_373_n N_A_225_74#_c_406_n 0.0145639f $X=1.605 $Y=0 $X2=0 $Y2=0
cc_216 N_VGND_c_375_n N_A_225_74#_c_406_n 0.0119984f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_217 N_VGND_M1009_d N_A_225_74#_c_407_n 0.00358162f $X=1.56 $Y=0.37 $X2=0
+ $Y2=0
cc_218 N_VGND_c_372_n N_A_225_74#_c_407_n 0.0248957f $X=1.77 $Y=0.675 $X2=0
+ $Y2=0
cc_219 N_VGND_c_374_n N_A_225_74#_c_409_n 0.044415f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_220 N_VGND_c_375_n N_A_225_74#_c_409_n 0.0381644f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_221 N_VGND_c_372_n N_A_225_74#_c_410_n 0.00795492f $X=1.77 $Y=0.675 $X2=0
+ $Y2=0
cc_222 N_VGND_c_374_n N_A_225_74#_c_410_n 0.00751083f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_223 N_VGND_c_375_n N_A_225_74#_c_410_n 0.00615808f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_224 N_VGND_c_374_n N_A_225_74#_c_411_n 0.0126895f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_225 N_VGND_c_375_n N_A_225_74#_c_411_n 0.0105154f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_226 N_A_225_74#_c_407_n A_426_74# 0.00122604f $X=2.105 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_227 N_A_225_74#_c_417_n A_426_74# 0.00479875f $X=2.19 $Y=1.01 $X2=-0.19
+ $Y2=-0.245
cc_228 N_A_225_74#_c_409_n A_426_74# 0.00141176f $X=3.395 $Y=0.435 $X2=-0.19
+ $Y2=-0.245
