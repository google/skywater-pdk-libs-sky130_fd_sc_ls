* File: sky130_fd_sc_ls__a311o_4.spice
* Created: Fri Aug 28 12:57:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a311o_4.pex.spice"
.subckt sky130_fd_sc_ls__a311o_4  VNB VPB C1 B1 A3 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* A3	A3
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_C1_M1015_g N_A_154_392#_M1015_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75004 A=0.096 P=1.58 MULT=1
MM1024 N_VGND_M1024_d N_C1_M1024_g N_A_154_392#_M1015_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75003.6 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1024_d N_B1_M1000_g N_A_154_392#_M1000_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001
+ SB=75003.2 A=0.096 P=1.58 MULT=1
MM1023 N_VGND_M1023_d N_B1_M1023_g N_A_154_392#_M1000_s VNB NSHORT L=0.15 W=0.64
+ AD=0.108058 AS=0.0896 PD=0.987826 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75002.7 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1023_d N_A_154_392#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.124942 AS=0.1036 PD=1.14217 PS=1.02 NRD=7.296 NRS=0 M=1 R=4.93333
+ SA=75001.7 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_154_392#_M1009_g N_X_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.121562 AS=0.1036 PD=1.08 PS=1.02 NRD=3.24 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1009_d N_A_154_392#_M1017_g N_X_M1017_s VNB NSHORT L=0.15 W=0.74
+ AD=0.121562 AS=0.1036 PD=1.08 PS=1.02 NRD=4.044 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1021_d N_A_154_392#_M1021_g N_X_M1017_s VNB NSHORT L=0.15 W=0.74
+ AD=0.130894 AS=0.1036 PD=1.15826 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003
+ SB=75001 A=0.111 P=1.78 MULT=1
MM1010 N_A_888_105#_M1010_d N_A3_M1010_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.113206 PD=0.92 PS=1.00174 NRD=0 NRS=11.712 M=1 R=4.26667
+ SA=75003.4 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1014 N_A_888_105#_M1010_d N_A3_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.9
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 N_A_154_392#_M1004_d N_A1_M1004_g N_A_1081_39#_M1004_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.3055 PD=0.92 PS=2.71 NRD=0 NRS=79.188 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1005 N_A_154_392#_M1004_d N_A1_M1005_g N_A_1081_39#_M1005_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1088 PD=0.92 PS=0.98 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1011 N_A_1081_39#_M1005_s N_A2_M1011_g N_A_888_105#_M1011_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1088 AS=0.0896 PD=0.98 PS=0.92 NRD=11.244 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1020 N_A_1081_39#_M1020_d N_A2_M1020_g N_A_888_105#_M1011_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_A_154_392#_M1002_d N_C1_M1002_g N_A_69_392#_M1002_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1008 N_A_154_392#_M1002_d N_C1_M1008_g N_A_69_392#_M1008_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.6 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1012 N_A_69_392#_M1008_s N_B1_M1012_g N_A_334_392#_M1012_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1019 N_A_69_392#_M1019_d N_B1_M1019_g N_A_334_392#_M1012_s VPB PHIGHVT L=0.15
+ W=1 AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.5 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1007 N_X_M1007_d N_A_154_392#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75004 A=0.168 P=2.54 MULT=1
MM1018 N_X_M1007_d N_A_154_392#_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75003.6 A=0.168 P=2.54 MULT=1
MM1022 N_X_M1022_d N_A_154_392#_M1022_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1025 N_X_M1022_d N_A_154_392#_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.210264 PD=1.42 PS=1.56906 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1026 N_A_334_392#_M1026_d N_A3_M1026_g N_VPWR_M1025_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.187736 PD=1.3 PS=1.40094 NRD=1.9503 NRS=14.7553 M=1 R=6.66667
+ SA=75002.1 SB=75002.5 A=0.15 P=2.3 MULT=1
MM1027 N_A_334_392#_M1026_d N_A3_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75002.5
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1006 N_A_334_392#_M1006_d N_A1_M1006_g N_VPWR_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75003
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1016 N_A_334_392#_M1006_d N_A1_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.165 PD=1.3 PS=1.33 NRD=1.9503 NRS=4.9053 M=1 R=6.66667 SA=75003.4
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1003 N_A_334_392#_M1003_d N_A2_M1003_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.165 PD=1.3 PS=1.33 NRD=1.9503 NRS=4.9053 M=1 R=6.66667 SA=75003.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1013 N_A_334_392#_M1003_d N_A2_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75004.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=14.9916 P=19.84
c_71 VNB 0 1.44209e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__a311o_4.pxi.spice"
*
.ends
*
*
