* NGSPICE file created from sky130_fd_sc_ls__nand2_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nand2_1 A B VGND VNB VPB VPWR Y
M1000 Y A a_117_74# VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.776e+11p ps=1.96e+06u
M1001 Y B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=6.384e+11p ps=5.62e+06u
M1002 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_117_74# B VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends

