* File: sky130_fd_sc_ls__clkinv_4.pex.spice
* Created: Fri Aug 28 13:11:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__CLKINV_4%A 1 3 4 8 10 12 13 15 18 20 22 23 25 28 30
+ 32 35 37 39 40 41 42 43 62
r108 62 63 1.97003 $w=3.67e-07 $l=1.5e-08 $layer=POLY_cond $X=2.805 $Y=1.557
+ $X2=2.82 $Y2=1.557
r109 60 62 54.5041 $w=3.67e-07 $l=4.15e-07 $layer=POLY_cond $X=2.39 $Y=1.557
+ $X2=2.805 $Y2=1.557
r110 60 61 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.39
+ $Y=1.515 $X2=2.39 $Y2=1.515
r111 58 60 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=2.365 $Y=1.557
+ $X2=2.39 $Y2=1.557
r112 57 58 1.31335 $w=3.67e-07 $l=1e-08 $layer=POLY_cond $X=2.355 $Y=1.557
+ $X2=2.365 $Y2=1.557
r113 56 57 65.6676 $w=3.67e-07 $l=5e-07 $layer=POLY_cond $X=1.855 $Y=1.557
+ $X2=2.355 $Y2=1.557
r114 55 56 7.88011 $w=3.67e-07 $l=6e-08 $layer=POLY_cond $X=1.795 $Y=1.557
+ $X2=1.855 $Y2=1.557
r115 54 55 51.2207 $w=3.67e-07 $l=3.9e-07 $layer=POLY_cond $X=1.405 $Y=1.557
+ $X2=1.795 $Y2=1.557
r116 52 54 49.2507 $w=3.67e-07 $l=3.75e-07 $layer=POLY_cond $X=1.03 $Y=1.557
+ $X2=1.405 $Y2=1.557
r117 52 53 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.03
+ $Y=1.515 $X2=1.03 $Y2=1.515
r118 50 52 9.85014 $w=3.67e-07 $l=7.5e-08 $layer=POLY_cond $X=0.955 $Y=1.557
+ $X2=1.03 $Y2=1.557
r119 49 50 1.97003 $w=3.67e-07 $l=1.5e-08 $layer=POLY_cond $X=0.94 $Y=1.557
+ $X2=0.955 $Y2=1.557
r120 43 61 6.70025 $w=4.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.39 $Y2=1.565
r121 42 61 6.16423 $w=4.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.39 $Y2=1.565
r122 41 42 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=2.16 $Y2=1.565
r123 40 41 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r124 40 53 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.03 $Y2=1.565
r125 39 53 8.30831 $w=4.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.03 $Y2=1.565
r126 33 63 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=1.35
+ $X2=2.82 $Y2=1.557
r127 33 35 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.82 $Y=1.35
+ $X2=2.82 $Y2=0.61
r128 30 62 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.805 $Y=1.765
+ $X2=2.805 $Y2=1.557
r129 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.805 $Y=1.765
+ $X2=2.805 $Y2=2.4
r130 26 58 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.365 $Y=1.35
+ $X2=2.365 $Y2=1.557
r131 26 28 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.365 $Y=1.35
+ $X2=2.365 $Y2=0.61
r132 23 57 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.355 $Y=1.765
+ $X2=2.355 $Y2=1.557
r133 23 25 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.355 $Y=1.765
+ $X2=2.355 $Y2=2.4
r134 20 56 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.557
r135 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r136 16 55 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.795 $Y=1.35
+ $X2=1.795 $Y2=1.557
r137 16 18 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.795 $Y=1.35
+ $X2=1.795 $Y2=0.61
r138 13 54 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.557
r139 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r140 10 50 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.557
r141 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r142 6 49 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=1.35 $X2=0.94
+ $Y2=1.557
r143 6 8 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.94 $Y=1.35 $X2=0.94
+ $Y2=0.61
r144 5 37 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.595 $Y=1.605
+ $X2=0.505 $Y2=1.605
r145 4 49 27.1901 $w=3.67e-07 $l=9.60469e-08 $layer=POLY_cond $X=0.865 $Y=1.605
+ $X2=0.94 $Y2=1.557
r146 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.865 $Y=1.605
+ $X2=0.595 $Y2=1.605
r147 1 37 64.3434 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.605
r148 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_4%VPWR 1 2 3 4 13 15 19 23 25 27 30 31 32 38
+ 42 51 55
r53 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 46 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 46 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 43 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.12 $Y2=3.33
r60 43 45 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 42 54 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.137 $Y2=3.33
r62 42 45 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 38 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.12 $Y2=3.33
r64 38 40 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 37 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r66 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 34 48 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r68 34 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 32 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r70 32 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 32 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 30 36 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r73 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.18 $Y2=3.33
r74 29 40 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r75 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.18 $Y2=3.33
r76 25 54 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.137 $Y2=3.33
r77 25 27 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=2.455
r78 21 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=3.33
r79 21 23 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=2.455
r80 17 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r81 17 19 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.455
r82 13 48 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r83 13 15 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.455
r84 4 27 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=2.88
+ $Y=1.84 $X2=3.08 $Y2=2.455
r85 3 23 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.455
r86 2 19 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.455
r87 1 15 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_4%Y 1 2 3 4 5 17 19 22 24 25 28 30 32 36 40
+ 42 44 52 53 55 56 58 61
r108 60 61 32.8196 $w=2.28e-07 $l=6.55e-07 $layer=LI1_cond $X=3.12 $Y=1.95
+ $X2=3.12 $Y2=1.295
r109 59 61 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.18
+ $X2=3.12 $Y2=1.295
r110 51 53 10.9648 $w=7.23e-07 $l=1.65e-07 $layer=LI1_cond $X=1.58 $Y=0.817
+ $X2=1.745 $Y2=0.817
r111 51 52 17.9763 $w=7.23e-07 $l=5.9e-07 $layer=LI1_cond $X=1.58 $Y=0.817
+ $X2=0.99 $Y2=0.817
r112 46 49 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.35 $Y=2.035
+ $X2=0.73 $Y2=2.035
r113 45 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=2.035
+ $X2=2.58 $Y2=2.035
r114 44 60 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.005 $Y=2.035
+ $X2=3.12 $Y2=1.95
r115 44 45 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.005 $Y=2.035
+ $X2=2.745 $Y2=2.035
r116 43 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=1.095
+ $X2=2.58 $Y2=1.095
r117 42 59 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.005 $Y=1.095
+ $X2=3.12 $Y2=1.18
r118 42 43 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.005 $Y=1.095
+ $X2=2.745 $Y2=1.095
r119 38 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=2.12
+ $X2=2.58 $Y2=2.035
r120 38 40 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.58 $Y=2.12
+ $X2=2.58 $Y2=2.815
r121 34 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=1.01
+ $X2=2.58 $Y2=1.095
r122 34 36 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=2.58 $Y=1.01 $X2=2.58
+ $Y2=0.61
r123 33 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=2.035
+ $X2=1.63 $Y2=2.035
r124 32 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=2.035
+ $X2=2.58 $Y2=2.035
r125 32 33 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.415 $Y=2.035
+ $X2=1.795 $Y2=2.035
r126 30 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=1.095
+ $X2=2.58 $Y2=1.095
r127 30 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.415 $Y=1.095
+ $X2=1.745 $Y2=1.095
r128 26 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=2.12
+ $X2=1.63 $Y2=2.035
r129 26 28 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.63 $Y=2.12
+ $X2=1.63 $Y2=2.815
r130 25 49 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.035
+ $X2=0.73 $Y2=2.035
r131 24 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=1.63 $Y2=2.035
r132 24 25 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=0.895 $Y2=2.035
r133 22 49 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.73 $Y=2.815
+ $X2=0.73 $Y2=2.12
r134 19 52 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=0.435 $Y=1.095
+ $X2=0.99 $Y2=1.095
r135 17 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.35 $Y=1.95
+ $X2=0.35 $Y2=2.035
r136 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.35 $Y=1.18
+ $X2=0.435 $Y2=1.095
r137 16 17 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.35 $Y=1.18
+ $X2=0.35 $Y2=1.95
r138 5 58 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.84 $X2=2.58 $Y2=2.035
r139 5 40 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.84 $X2=2.58 $Y2=2.815
r140 4 55 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.035
r141 4 28 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.815
r142 3 49 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.035
r143 3 22 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r144 2 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.44
+ $Y=0.4 $X2=2.58 $Y2=0.61
r145 1 51 91 $w=1.7e-07 $l=6.65977e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.4 $X2=1.58 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_4%VGND 1 2 3 12 14 16 18 20 25 31 38 42
r31 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r32 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r33 32 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r34 31 36 9.12071 $w=7.29e-07 $l=5.45e-07 $layer=LI1_cond $X=0.41 $Y=0 $X2=0.41
+ $Y2=0.545
r35 31 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r37 29 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r38 29 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r39 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r40 26 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.08
+ $Y2=0
r41 26 28 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.64
+ $Y2=0
r42 25 41 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.137
+ $Y2=0
r43 25 28 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.64
+ $Y2=0
r44 21 31 9.58964 $w=1.7e-07 $l=4.1e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.41
+ $Y2=0
r45 21 23 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=1.68
+ $Y2=0
r46 20 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.915 $Y=0 $X2=2.08
+ $Y2=0
r47 20 23 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=0 $X2=1.68
+ $Y2=0
r48 18 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r49 18 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r50 18 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 14 41 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.137 $Y2=0
r52 14 16 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.61
r53 10 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0
r54 10 12 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0.61
r55 3 16 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.4 $X2=3.08 $Y2=0.61
r56 2 12 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=1.87
+ $Y=0.4 $X2=2.08 $Y2=0.61
r57 1 36 91 $w=1.7e-07 $l=5.88048e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.4 $X2=0.655 $Y2=0.545
.ends

