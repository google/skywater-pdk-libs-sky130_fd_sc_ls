* File: sky130_fd_sc_ls__nor2_1.pex.spice
* Created: Wed Sep  2 11:13:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NOR2_1%A 1 3 6 8 12
r24 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.465 $X2=0.29 $Y2=1.465
r25 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.29 $Y=1.665 $X2=0.29
+ $Y2=1.465
r26 4 11 39.305 $w=3.85e-07 $l=2.29783e-07 $layer=POLY_cond $X=0.515 $Y=1.3
+ $X2=0.36 $Y2=1.465
r27 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.515 $Y=1.3 $X2=0.515
+ $Y2=0.74
r28 1 11 56.2063 $w=3.85e-07 $l=3.65377e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.36 $Y2=1.465
r29 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2_1%B 1 3 6 8 12
r20 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.465 $X2=1.15 $Y2=1.465
r21 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.15 $Y=1.665 $X2=1.15
+ $Y2=1.465
r22 4 11 39.4323 $w=3.92e-07 $l=2.20624e-07 $layer=POLY_cond $X=0.945 $Y=1.3
+ $X2=1.075 $Y2=1.465
r23 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.945 $Y=1.3 $X2=0.945
+ $Y2=0.74
r24 1 11 56.0318 $w=3.92e-07 $l=3.67423e-07 $layer=POLY_cond $X=0.925 $Y=1.765
+ $X2=1.075 $Y2=1.465
r25 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.925 $Y=1.765
+ $X2=0.925 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2_1%VPWR 1 4 6 10 14 15
r15 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r16 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r17 12 18 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r18 12 14 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r19 10 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r20 10 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r21 6 9 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115 $X2=0.28
+ $Y2=2.815
r22 4 18 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r23 4 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245 $X2=0.28
+ $Y2=2.815
r24 1 9 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r25 1 6 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2_1%Y 1 2 9 12 13 14 15
r26 14 15 7.05312 $w=6.4e-07 $l=3.7e-07 $layer=LI1_cond $X=0.98 $Y=2.405
+ $X2=0.98 $Y2=2.775
r27 14 19 5.52812 $w=6.4e-07 $l=2.9e-07 $layer=LI1_cond $X=0.98 $Y=2.405
+ $X2=0.98 $Y2=2.115
r28 12 19 10.6252 $w=6.4e-07 $l=3.22102e-07 $layer=LI1_cond $X=0.73 $Y=1.95
+ $X2=0.98 $Y2=2.115
r29 12 13 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.73 $Y=1.95
+ $X2=0.73 $Y2=1.13
r30 7 13 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.69 $Y=1.005
+ $X2=0.69 $Y2=1.13
r31 7 9 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=0.69 $Y=1.005 $X2=0.69
+ $Y2=0.515
r32 2 15 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1 $Y=1.84
+ $X2=1.15 $Y2=2.815
r33 2 19 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1 $Y=1.84
+ $X2=1.15 $Y2=2.115
r34 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.59
+ $Y=0.37 $X2=0.73 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NOR2_1%VGND 1 2 7 9 11 13 15 17 27
r21 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r22 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r23 18 23 3.98448 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.192
+ $Y2=0
r24 18 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.72
+ $Y2=0
r25 17 26 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=1.217
+ $Y2=0
r26 17 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=0.72
+ $Y2=0
r27 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r28 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r29 15 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r30 11 26 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=1.16 $Y=0.085
+ $X2=1.217 $Y2=0
r31 11 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.16 $Y=0.085
+ $X2=1.16 $Y2=0.515
r32 7 23 3.15868 $w=2.5e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.192 $Y2=0
r33 7 9 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.26 $Y=0.085 $X2=0.26
+ $Y2=0.515
r34 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.02
+ $Y=0.37 $X2=1.16 $Y2=0.515
r35 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.37 $X2=0.3 $Y2=0.515
.ends

