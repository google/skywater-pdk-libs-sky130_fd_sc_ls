# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__o21ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__o21ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.320000 1.795000 1.650000 ;
        RECT 1.085000 1.650000 1.795000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.350000 5.635000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.180000 3.165000 1.550000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.478400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.280000 0.595000 2.530000 0.840000 ;
        RECT 2.280000 0.840000 3.505000 1.010000 ;
        RECT 2.365000 1.820000 3.715000 1.950000 ;
        RECT 2.365000 1.950000 5.190000 2.120000 ;
        RECT 3.220000 0.595000 3.505000 0.840000 ;
        RECT 3.335000 1.010000 3.505000 1.550000 ;
        RECT 3.335000 1.550000 3.715000 1.820000 ;
        RECT 3.960000 2.120000 4.290000 2.735000 ;
        RECT 4.860000 2.120000 5.190000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 0.980000 ;
      RECT 0.115000  0.980000 2.100000 1.010000 ;
      RECT 0.115000  1.010000 1.225000 1.150000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.545000  0.085000 0.875000 0.810000 ;
      RECT 0.565000  1.820000 0.895000 1.950000 ;
      RECT 0.565000  1.950000 1.795000 2.120000 ;
      RECT 0.565000  2.120000 0.895000 2.980000 ;
      RECT 1.055000  0.350000 1.225000 0.840000 ;
      RECT 1.055000  0.840000 2.100000 0.980000 ;
      RECT 1.095000  2.290000 1.265000 3.245000 ;
      RECT 1.405000  0.085000 1.735000 0.670000 ;
      RECT 1.465000  2.120000 1.795000 2.290000 ;
      RECT 1.465000  2.290000 3.790000 2.460000 ;
      RECT 1.465000  2.460000 1.795000 2.980000 ;
      RECT 1.930000  0.255000 3.845000 0.425000 ;
      RECT 1.930000  0.425000 2.100000 0.840000 ;
      RECT 1.995000  2.630000 2.245000 3.245000 ;
      RECT 2.710000  0.425000 3.040000 0.670000 ;
      RECT 2.900000  2.630000 3.230000 3.245000 ;
      RECT 3.460000  2.460000 3.790000 2.905000 ;
      RECT 3.460000  2.905000 5.640000 3.075000 ;
      RECT 3.675000  0.425000 3.845000 1.010000 ;
      RECT 3.675000  1.010000 5.645000 1.180000 ;
      RECT 4.025000  0.085000 4.355000 0.840000 ;
      RECT 4.490000  2.290000 4.660000 2.905000 ;
      RECT 4.535000  0.350000 4.705000 1.010000 ;
      RECT 4.885000  0.085000 5.215000 0.840000 ;
      RECT 5.390000  1.950000 5.640000 2.905000 ;
      RECT 5.395000  0.350000 5.645000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_ls__o21ai_4
END LIBRARY
