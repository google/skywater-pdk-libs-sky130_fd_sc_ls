* File: sky130_fd_sc_ls__dfrtp_4.pex.spice
* Created: Fri Aug 28 13:14:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DFRTP_4%D 2 4 5 7 10 12 13 14 19 20 23
r36 23 25 35.4289 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.42 $Y=1.845
+ $X2=0.42 $Y2=2.01
r37 23 24 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.845 $X2=0.385 $Y2=1.845
r38 19 21 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.42 $Y=1.165
+ $X2=0.42 $Y2=1
r39 19 20 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.165 $X2=0.385 $Y2=1.165
r40 14 24 5.61447 $w=3.88e-07 $l=1.9e-07 $layer=LI1_cond $X=0.32 $Y=2.035
+ $X2=0.32 $Y2=1.845
r41 13 24 5.31897 $w=3.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.32 $Y=1.665
+ $X2=0.32 $Y2=1.845
r42 12 13 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.32 $Y=1.295
+ $X2=0.32 $Y2=1.665
r43 12 20 3.84148 $w=3.88e-07 $l=1.3e-07 $layer=LI1_cond $X=0.32 $Y=1.295
+ $X2=0.32 $Y2=1.165
r44 10 21 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.545 $Y=0.6 $X2=0.545
+ $Y2=1
r45 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.5 $Y=2.465 $X2=0.5
+ $Y2=2.75
r46 4 5 54.6598 $w=1.94e-07 $l=2.27376e-07 $layer=POLY_cond $X=0.515 $Y=2.245
+ $X2=0.5 $Y2=2.465
r47 4 25 74.2101 $w=2.1e-07 $l=2.35e-07 $layer=POLY_cond $X=0.515 $Y=2.245
+ $X2=0.515 $Y2=2.01
r48 2 23 4.86635 $w=4e-07 $l=3.5e-08 $layer=POLY_cond $X=0.42 $Y=1.81 $X2=0.42
+ $Y2=1.845
r49 1 19 4.86635 $w=4e-07 $l=3.5e-08 $layer=POLY_cond $X=0.42 $Y=1.2 $X2=0.42
+ $Y2=1.165
r50 1 2 84.8135 $w=4e-07 $l=6.1e-07 $layer=POLY_cond $X=0.42 $Y=1.2 $X2=0.42
+ $Y2=1.81
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_4%CLK 3 7 8 11 13
c45 8 0 2.50248e-19 $X=2.16 $Y=1.665
c46 3 0 6.36774e-20 $X=1.945 $Y=2.46
r47 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.93 $Y=1.61
+ $X2=1.93 $Y2=1.775
r48 11 13 52.3316 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.93 $Y=1.61 $X2=1.93
+ $Y2=1.41
r49 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.93
+ $Y=1.61 $X2=1.93 $Y2=1.61
r50 8 12 6.19426 $w=4.53e-07 $l=2.3e-07 $layer=LI1_cond $X=2.16 $Y=1.545
+ $X2=1.93 $Y2=1.545
r51 7 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.965 $Y=0.965
+ $X2=1.965 $Y2=1.41
r52 3 14 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=1.945 $Y=2.46
+ $X2=1.945 $Y2=1.775
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_4%A_494_392# 1 2 7 9 10 13 16 18 20 21 22 23
+ 25 28 30 35 36 38 40 44 48 49 54 58 62 68 71
c189 54 0 1.90924e-19 $X=2.915 $Y=1.9
c190 44 0 9.26151e-20 $X=7.905 $Y=2.14
c191 36 0 2.17651e-19 $X=4.305 $Y=0.415
c192 28 0 4.38676e-20 $X=3.985 $Y=1.46
c193 16 0 1.85309e-19 $X=3.985 $Y=0.9
c194 7 0 4.12227e-19 $X=3.42 $Y=2.24
r195 70 71 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=7.905 $Y=1.18
+ $X2=8.19 $Y2=1.18
r196 68 77 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.71 $Y=1.18 $X2=7.71
+ $Y2=1.27
r197 67 70 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=7.71 $Y=1.18
+ $X2=7.905 $Y2=1.18
r198 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.71
+ $Y=1.18 $X2=7.71 $Y2=1.18
r199 62 64 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.48 $Y=0.34
+ $X2=5.48 $Y2=0.625
r200 58 60 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.39 $Y=0.415
+ $X2=4.39 $Y2=0.625
r201 57 73 13.4387 $w=2.69e-07 $l=7.5e-08 $layer=POLY_cond $X=3.37 $Y=1.85
+ $X2=3.37 $Y2=1.775
r202 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.37
+ $Y=1.85 $X2=3.37 $Y2=1.85
r203 54 56 11.3286 $w=4.9e-07 $l=4.55e-07 $layer=LI1_cond $X=2.915 $Y=1.9
+ $X2=3.37 $Y2=1.9
r204 52 53 6.10029 $w=4.58e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=0.72
+ $X2=2.785 $Y2=0.805
r205 49 52 7.93052 $w=4.58e-07 $l=3.05e-07 $layer=LI1_cond $X=2.785 $Y=0.415
+ $X2=2.785 $Y2=0.72
r206 48 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.19 $Y=1.015
+ $X2=8.19 $Y2=1.18
r207 47 48 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.19 $Y=0.425
+ $X2=8.19 $Y2=1.015
r208 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.905
+ $Y=2.14 $X2=7.905 $Y2=2.14
r209 42 70 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.905 $Y=1.345
+ $X2=7.905 $Y2=1.18
r210 42 44 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=7.905 $Y=1.345
+ $X2=7.905 $Y2=2.14
r211 41 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0.34
+ $X2=5.48 $Y2=0.34
r212 40 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.105 $Y=0.34
+ $X2=8.19 $Y2=0.425
r213 40 41 165.711 $w=1.68e-07 $l=2.54e-06 $layer=LI1_cond $X=8.105 $Y=0.34
+ $X2=5.565 $Y2=0.34
r214 39 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.475 $Y=0.625
+ $X2=4.39 $Y2=0.625
r215 38 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0.625
+ $X2=5.48 $Y2=0.625
r216 38 39 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.395 $Y=0.625
+ $X2=4.475 $Y2=0.625
r217 37 49 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.015 $Y=0.415
+ $X2=2.785 $Y2=0.415
r218 36 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.305 $Y=0.415
+ $X2=4.39 $Y2=0.415
r219 36 37 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=4.305 $Y=0.415
+ $X2=3.015 $Y2=0.415
r220 35 54 6.0248 $w=2e-07 $l=3.4e-07 $layer=LI1_cond $X=2.915 $Y=1.56 $X2=2.915
+ $Y2=1.9
r221 35 53 41.8682 $w=1.98e-07 $l=7.55e-07 $layer=LI1_cond $X=2.915 $Y=1.56
+ $X2=2.915 $Y2=0.805
r222 30 54 5.52759 $w=4.9e-07 $l=2.5437e-07 $layer=LI1_cond $X=2.77 $Y=2.092
+ $X2=2.915 $Y2=1.9
r223 30 32 5.85988 $w=2.93e-07 $l=1.5e-07 $layer=LI1_cond $X=2.77 $Y=2.092
+ $X2=2.62 $Y2=2.092
r224 26 28 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=3.875 $Y=1.46
+ $X2=3.985 $Y2=1.46
r225 23 45 50.2556 $w=3.62e-07 $l=3.02076e-07 $layer=POLY_cond $X=8.06 $Y=2.39
+ $X2=7.945 $Y2=2.14
r226 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.06 $Y=2.39
+ $X2=8.06 $Y2=2.675
r227 21 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.545 $Y=1.27
+ $X2=7.71 $Y2=1.27
r228 21 22 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=7.545 $Y=1.27
+ $X2=7.185 $Y2=1.27
r229 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.11 $Y=1.195
+ $X2=7.185 $Y2=1.27
r230 18 20 146.207 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=7.11 $Y=1.195
+ $X2=7.11 $Y2=0.74
r231 14 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.985 $Y=1.385
+ $X2=3.985 $Y2=1.46
r232 14 16 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.985 $Y=1.385
+ $X2=3.985 $Y2=0.9
r233 12 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.875 $Y=1.535
+ $X2=3.875 $Y2=1.46
r234 12 13 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.875 $Y=1.535
+ $X2=3.875 $Y2=1.685
r235 11 73 12.2038 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.535 $Y=1.775
+ $X2=3.37 $Y2=1.775
r236 10 13 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.8 $Y=1.775
+ $X2=3.875 $Y2=1.685
r237 10 11 103.008 $w=1.8e-07 $l=2.65e-07 $layer=POLY_cond $X=3.8 $Y=1.775
+ $X2=3.535 $Y2=1.775
r238 7 57 79.2394 $w=2.69e-07 $l=4.14246e-07 $layer=POLY_cond $X=3.42 $Y=2.24
+ $X2=3.37 $Y2=1.85
r239 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.42 $Y=2.24 $X2=3.42
+ $Y2=2.525
r240 2 32 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.47
+ $Y=1.96 $X2=2.62 $Y2=2.155
r241 1 52 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=2.57
+ $Y=0.595 $X2=2.72 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_4%A_834_355# 1 2 7 9 12 16 20 22 23 25 29 34
c87 34 0 1.52817e-19 $X=6.45 $Y=2.125
c88 29 0 1.42958e-20 $X=5.735 $Y=0.885
c89 23 0 5.12321e-20 $X=6.325 $Y=0.885
c90 20 0 3.05298e-19 $X=4.57 $Y=0.965
c91 12 0 1.36289e-19 $X=4.375 $Y=0.9
c92 7 0 1.60401e-19 $X=4.26 $Y=2.24
r93 28 30 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=5.9 $Y=0.885
+ $X2=6.24 $Y2=0.885
r94 28 29 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.9 $Y=0.885
+ $X2=5.735 $Y2=0.885
r95 23 30 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.325 $Y=0.885
+ $X2=6.24 $Y2=0.885
r96 23 25 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6.325 $Y=0.885
+ $X2=6.825 $Y2=0.885
r97 22 34 8.20383 $w=2.93e-07 $l=2.1e-07 $layer=LI1_cond $X=6.24 $Y=2.087
+ $X2=6.45 $Y2=2.087
r98 21 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.24 $Y=1.05
+ $X2=6.24 $Y2=0.885
r99 21 22 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=6.24 $Y=1.05
+ $X2=6.24 $Y2=1.94
r100 20 29 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=4.57 $Y=0.965
+ $X2=5.735 $Y2=0.965
r101 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.405
+ $Y=1.94 $X2=4.405 $Y2=1.94
r102 14 20 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=4.437 $Y=1.05
+ $X2=4.57 $Y2=0.965
r103 14 16 38.7047 $w=2.63e-07 $l=8.9e-07 $layer=LI1_cond $X=4.437 $Y=1.05
+ $X2=4.437 $Y2=1.94
r104 10 17 38.6446 $w=3.36e-07 $l=1.67481e-07 $layer=POLY_cond $X=4.375 $Y=1.775
+ $X2=4.37 $Y2=1.94
r105 10 12 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=4.375 $Y=1.775
+ $X2=4.375 $Y2=0.9
r106 7 17 58.0107 $w=3.36e-07 $l=3.50714e-07 $layer=POLY_cond $X=4.26 $Y=2.24
+ $X2=4.37 $Y2=1.94
r107 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.26 $Y=2.24 $X2=4.26
+ $Y2=2.525
r108 2 34 600 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=6.3
+ $Y=1.96 $X2=6.45 $Y2=2.125
r109 1 28 182 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_NDIFF $count=1 $X=5.76
+ $Y=0.37 $X2=5.9 $Y2=0.885
r110 1 25 91 $w=1.7e-07 $l=1.29719e-06 $layer=licon1_NDIFF $count=2 $X=5.76
+ $Y=0.37 $X2=6.825 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_4%RESET_B 4 6 8 9 11 12 13 17 19 20 22 24 25
+ 27 30 34 37 38 39 40 41 44 46 47 49 52 56 57 60
c232 56 0 1.17008e-19 $X=1.155 $Y=1.295
c233 52 0 1.66354e-20 $X=5.25 $Y=1.835
c234 44 0 1.36553e-19 $X=5.52 $Y=2.035
c235 41 0 1.63054e-19 $X=5.665 $Y=2.035
c236 37 0 1.42958e-20 $X=4.87 $Y=1.835
c237 20 0 1.20728e-19 $X=4.87 $Y=2.24
c238 12 0 1.19989e-19 $X=4.69 $Y=0.18
r239 60 62 41.3282 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.975
+ $X2=1.09 $Y2=2.14
r240 60 61 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.975 $X2=1.155 $Y2=1.975
r241 57 61 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.155 $Y=1.295
+ $X2=1.155 $Y2=1.975
r242 56 58 47.2161 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.295
+ $X2=1.09 $Y2=1.13
r243 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.295 $X2=1.155 $Y2=1.295
r244 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.25
+ $Y=1.835 $X2=5.25 $Y2=1.835
r245 49 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r246 47 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.975
+ $Y=2.11 $X2=8.975 $Y2=2.11
r247 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=2.035
+ $X2=8.88 $Y2=2.035
r248 44 53 7.17647 $w=4.48e-07 $l=2.7e-07 $layer=LI1_cond $X=5.52 $Y=1.895
+ $X2=5.25 $Y2=1.895
r249 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r250 41 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r251 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=8.88 $Y2=2.035
r252 40 41 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=5.665 $Y2=2.035
r253 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r254 38 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=5.52 $Y2=2.035
r255 38 39 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=1.345 $Y2=2.035
r256 36 52 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=4.96 $Y=1.835
+ $X2=5.25 $Y2=1.835
r257 36 37 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.96 $Y=1.835
+ $X2=4.87 $Y2=1.835
r258 32 34 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=4.765 $Y=1.26
+ $X2=4.885 $Y2=1.26
r259 28 64 38.6072 $w=2.91e-07 $l=2.03101e-07 $layer=POLY_cond $X=9.06 $Y=1.945
+ $X2=8.975 $Y2=2.11
r260 28 30 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=9.06 $Y=1.945
+ $X2=9.06 $Y2=0.615
r261 25 64 57.6553 $w=2.91e-07 $l=3.01662e-07 $layer=POLY_cond $X=9.02 $Y=2.39
+ $X2=8.975 $Y2=2.11
r262 25 27 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.02 $Y=2.39
+ $X2=9.02 $Y2=2.675
r263 24 37 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=4.885 $Y=1.67
+ $X2=4.87 $Y2=1.835
r264 23 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.885 $Y=1.335
+ $X2=4.885 $Y2=1.26
r265 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=4.885 $Y=1.335
+ $X2=4.885 $Y2=1.67
r266 20 22 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.87 $Y=2.24
+ $X2=4.87 $Y2=2.525
r267 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.87 $Y=2.15 $X2=4.87
+ $Y2=2.24
r268 18 37 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=4.87 $Y=2
+ $X2=4.87 $Y2=1.835
r269 18 19 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=4.87 $Y=2 $X2=4.87
+ $Y2=2.15
r270 15 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.765 $Y=1.185
+ $X2=4.765 $Y2=1.26
r271 15 17 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.765 $Y=1.185
+ $X2=4.765 $Y2=0.9
r272 14 17 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=4.765 $Y=0.255
+ $X2=4.765 $Y2=0.9
r273 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.69 $Y=0.18
+ $X2=4.765 $Y2=0.255
r274 12 13 1886.98 $w=1.5e-07 $l=3.68e-06 $layer=POLY_cond $X=4.69 $Y=0.18
+ $X2=1.01 $Y2=0.18
r275 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.95 $Y=2.465
+ $X2=0.95 $Y2=2.75
r276 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.95 $Y=2.375 $X2=0.95
+ $Y2=2.465
r277 8 62 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.95 $Y=2.375
+ $X2=0.95 $Y2=2.14
r278 6 60 7.8587 $w=4.6e-07 $l=6.5e-08 $layer=POLY_cond $X=1.09 $Y=1.91 $X2=1.09
+ $Y2=1.975
r279 5 56 7.8587 $w=4.6e-07 $l=6.5e-08 $layer=POLY_cond $X=1.09 $Y=1.36 $X2=1.09
+ $Y2=1.295
r280 5 6 66.4967 $w=4.6e-07 $l=5.5e-07 $layer=POLY_cond $X=1.09 $Y=1.36 $X2=1.09
+ $Y2=1.91
r281 4 58 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.935 $Y=0.6
+ $X2=0.935 $Y2=1.13
r282 1 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.935 $Y=0.255
+ $X2=1.01 $Y2=0.18
r283 1 4 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.935 $Y=0.255
+ $X2=0.935 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_4%A_299_392# 1 2 9 11 13 15 17 18 19 20 21 24
+ 26 27 28 30 31 34 35 37 38 42 44 45 48 52 55 56 59 61 63 64 70 71 79
c232 71 0 1.76168e-19 $X=5.56 $Y=2.375
c233 70 0 2.76281e-19 $X=5.56 $Y=2.375
c234 61 0 1.17008e-19 $X=1.71 $Y=1.055
c235 59 0 1.35587e-19 $X=6.87 $Y=2.405
c236 55 0 3.79882e-20 $X=2.54 $Y=1.455
c237 20 0 2.7373e-20 $X=3.41 $Y=1.4
c238 17 0 7.60353e-20 $X=2.905 $Y=3.075
c239 15 0 7.00451e-20 $X=2.912 $Y=2.173
c240 11 0 8.78006e-20 $X=2.495 $Y=1.41
c241 9 0 1.23001e-19 $X=2.395 $Y=2.46
r242 77 90 41.4908 $w=2.73e-07 $l=2.35e-07 $layer=POLY_cond $X=6.66 $Y=1.425
+ $X2=6.66 $Y2=1.66
r243 76 79 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=6.66 $Y=1.425
+ $X2=6.87 $Y2=1.425
r244 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.66
+ $Y=1.425 $X2=6.66 $Y2=1.425
r245 71 85 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=5.56 $Y=2.375
+ $X2=5.385 $Y2=2.375
r246 70 73 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=5.56 $Y=2.375
+ $X2=5.56 $Y2=2.49
r247 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.56
+ $Y=2.375 $X2=5.56 $Y2=2.375
r248 68 84 49.1244 $w=3.65e-07 $l=3.72e-07 $layer=POLY_cond $X=2.54 $Y=1.55
+ $X2=2.912 $Y2=1.55
r249 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.54
+ $Y=1.61 $X2=2.54 $Y2=1.61
r250 63 64 9.9702 $w=3.48e-07 $l=2.1e-07 $layer=LI1_cond $X=1.63 $Y=2.155
+ $X2=1.63 $Y2=1.945
r251 58 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.87 $Y=1.59
+ $X2=6.87 $Y2=1.425
r252 58 59 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=6.87 $Y=1.59
+ $X2=6.87 $Y2=2.405
r253 57 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=2.49
+ $X2=5.56 $Y2=2.49
r254 56 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.785 $Y=2.49
+ $X2=6.87 $Y2=2.405
r255 56 57 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=6.785 $Y=2.49
+ $X2=5.725 $Y2=2.49
r256 55 67 9.95263 $w=1.9e-07 $l=1.55e-07 $layer=LI1_cond $X=2.54 $Y=1.455
+ $X2=2.54 $Y2=1.61
r257 54 55 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=2.54 $Y=1.14
+ $X2=2.54 $Y2=1.455
r258 53 61 3.3845 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.875 $Y=1.055
+ $X2=1.665 $Y2=1.055
r259 52 54 7.79998 $w=1.57e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=2.54 $Y2=1.14
r260 52 53 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=1.875 $Y2=1.055
r261 50 61 3.19717 $w=2.95e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.54 $Y=1.14
+ $X2=1.665 $Y2=1.055
r262 50 64 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.54 $Y=1.14
+ $X2=1.54 $Y2=1.945
r263 46 61 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.97
+ $X2=1.665 $Y2=1.055
r264 46 48 6.99698 $w=4.18e-07 $l=2.55e-07 $layer=LI1_cond $X=1.665 $Y=0.97
+ $X2=1.665 $Y2=0.715
r265 40 42 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=8.16 $Y=1.585
+ $X2=8.16 $Y2=0.615
r266 39 90 16.7618 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.825 $Y=1.66
+ $X2=6.66 $Y2=1.66
r267 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.085 $Y=1.66
+ $X2=8.16 $Y2=1.585
r268 38 39 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=8.085 $Y=1.66
+ $X2=6.825 $Y2=1.66
r269 35 90 49.4375 $w=2.73e-07 $l=2.32379e-07 $layer=POLY_cond $X=6.675 $Y=1.885
+ $X2=6.66 $Y2=1.66
r270 35 37 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.675 $Y=1.885
+ $X2=6.675 $Y2=2.46
r271 33 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=2.54
+ $X2=5.385 $Y2=2.375
r272 33 34 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=5.385 $Y=2.54
+ $X2=5.385 $Y2=3.075
r273 32 45 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.96 $Y=3.15 $X2=3.87
+ $Y2=3.15
r274 31 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.31 $Y=3.15
+ $X2=5.385 $Y2=3.075
r275 31 32 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=5.31 $Y=3.15
+ $X2=3.96 $Y2=3.15
r276 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.87 $Y=2.81
+ $X2=3.87 $Y2=2.525
r277 27 45 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.87 $Y=3.075
+ $X2=3.87 $Y2=3.15
r278 26 28 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.87 $Y=2.9 $X2=3.87
+ $Y2=2.81
r279 26 27 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.87 $Y=2.9
+ $X2=3.87 $Y2=3.075
r280 22 24 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=3.485 $Y=1.325
+ $X2=3.485 $Y2=0.9
r281 21 84 35.4153 $w=3.65e-07 $l=2.07846e-07 $layer=POLY_cond $X=3.05 $Y=1.4
+ $X2=2.912 $Y2=1.55
r282 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.41 $Y=1.4
+ $X2=3.485 $Y2=1.325
r283 20 21 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.41 $Y=1.4
+ $X2=3.05 $Y2=1.4
r284 18 45 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.78 $Y=3.15 $X2=3.87
+ $Y2=3.15
r285 18 19 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.78 $Y=3.15 $X2=2.98
+ $Y2=3.15
r286 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.905 $Y=3.075
+ $X2=2.98 $Y2=3.15
r287 17 44 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.905 $Y=3.075
+ $X2=2.905 $Y2=2.255
r288 15 44 36.4579 $w=1.65e-07 $l=8.2e-08 $layer=POLY_cond $X=2.912 $Y=2.173
+ $X2=2.912 $Y2=2.255
r289 14 84 21.4198 $w=1.65e-07 $l=2.25e-07 $layer=POLY_cond $X=2.912 $Y=1.775
+ $X2=2.912 $Y2=1.55
r290 14 15 173.376 $w=1.65e-07 $l=3.98e-07 $layer=POLY_cond $X=2.912 $Y=1.775
+ $X2=2.912 $Y2=2.173
r291 11 68 5.94247 $w=3.65e-07 $l=4.5e-08 $layer=POLY_cond $X=2.495 $Y=1.55
+ $X2=2.54 $Y2=1.55
r292 11 81 13.2055 $w=3.65e-07 $l=1e-07 $layer=POLY_cond $X=2.495 $Y=1.55
+ $X2=2.395 $Y2=1.55
r293 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.495 $Y=1.41
+ $X2=2.495 $Y2=0.965
r294 7 81 23.6381 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.395 $Y=1.775
+ $X2=2.395 $Y2=1.55
r295 7 9 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=2.395 $Y=1.775
+ $X2=2.395 $Y2=2.46
r296 2 63 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.96 $X2=1.64 $Y2=2.155
r297 1 61 182 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_NDIFF $count=1 $X=1.565
+ $Y=0.59 $X2=1.71 $Y2=1.055
r298 1 48 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.565
+ $Y=0.59 $X2=1.71 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_4%A_699_463# 1 2 3 10 12 15 17 18 19 20 21 27
+ 30 31 33 37 39 40 43
c138 40 0 2.07252e-19 $X=4.097 $Y=2.4
c139 39 0 3.12839e-20 $X=4.097 $Y=2.485
c140 30 0 1.38917e-19 $X=4.83 $Y=2.295
c141 27 0 1.50343e-19 $X=4.745 $Y=2.485
c142 21 0 2.36436e-19 $X=3.965 $Y=2.64
c143 20 0 1.30745e-19 $X=6.225 $Y=1.73
c144 18 0 2.99607e-19 $X=5.76 $Y=1.385
c145 15 0 5.6074e-20 $X=6.225 $Y=1.885
r146 43 45 8.354 $w=3.87e-07 $l=2.65e-07 $layer=LI1_cond $X=4.83 $Y=2.525
+ $X2=5.095 $Y2=2.525
r147 39 40 5.17317 $w=2.63e-07 $l=8.5e-08 $layer=LI1_cond $X=4.097 $Y=2.485
+ $X2=4.097 $Y2=2.4
r148 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.82
+ $Y=1.385 $X2=5.82 $Y2=1.385
r149 31 33 37.2486 $w=2.78e-07 $l=9.05e-07 $layer=LI1_cond $X=4.915 $Y=1.36
+ $X2=5.82 $Y2=1.36
r150 30 43 5.57805 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=4.83 $Y=2.295
+ $X2=4.83 $Y2=2.525
r151 29 31 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.83 $Y=1.5
+ $X2=4.915 $Y2=1.36
r152 29 30 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=4.83 $Y=1.5
+ $X2=4.83 $Y2=2.295
r153 28 39 3.33486 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.23 $Y=2.485
+ $X2=4.097 $Y2=2.485
r154 27 43 6.57826 $w=3.87e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.745 $Y=2.485
+ $X2=4.83 $Y2=2.525
r155 27 28 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.745 $Y=2.485
+ $X2=4.23 $Y2=2.485
r156 25 37 11.3867 $w=3e-07 $l=3.62767e-07 $layer=LI1_cond $X=4.05 $Y=1.05
+ $X2=3.77 $Y2=0.86
r157 25 40 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=4.05 $Y=1.05
+ $X2=4.05 $Y2=2.4
r158 21 39 6.7407 $w=2.63e-07 $l=1.55e-07 $layer=LI1_cond $X=4.097 $Y=2.64
+ $X2=4.097 $Y2=2.485
r159 21 23 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=3.965 $Y=2.64
+ $X2=3.645 $Y2=2.64
r160 19 34 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=6.135 $Y=1.385
+ $X2=5.82 $Y2=1.385
r161 18 34 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=5.76 $Y=1.385
+ $X2=5.82 $Y2=1.385
r162 15 20 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=6.225 $Y=1.885
+ $X2=6.225 $Y2=1.73
r163 15 17 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.225 $Y=1.885
+ $X2=6.225 $Y2=2.46
r164 13 19 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.21 $Y=1.55
+ $X2=6.135 $Y2=1.385
r165 13 20 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.21 $Y=1.55
+ $X2=6.21 $Y2=1.73
r166 10 18 17.4878 $w=4.41e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.685 $Y=1.22
+ $X2=5.76 $Y2=1.385
r167 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.685 $Y=1.22
+ $X2=5.685 $Y2=0.74
r168 3 45 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=4.945
+ $Y=2.315 $X2=5.095 $Y2=2.525
r169 2 23 600 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=3.495
+ $Y=2.315 $X2=3.645 $Y2=2.61
r170 1 37 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.69 $X2=3.77 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_4%A_1678_395# 1 2 8 9 11 16 18 19 20 23 24 25
+ 28 31 32 36 41 43
c124 31 0 1.27304e-19 $X=9.86 $Y=1.875
c125 24 0 1.26505e-19 $X=9.775 $Y=1.96
c126 18 0 9.26151e-20 $X=8.492 $Y=1.975
r127 39 41 3.90026 $w=4.58e-07 $l=1.5e-07 $layer=LI1_cond $X=9.245 $Y=2.675
+ $X2=9.395 $Y2=2.675
r128 36 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.61 $Y=1.2
+ $X2=8.61 $Y2=1.365
r129 36 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.61 $Y=1.2
+ $X2=8.61 $Y2=1.035
r130 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.61
+ $Y=1.2 $X2=8.61 $Y2=1.2
r131 32 35 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.61 $Y=1.12 $X2=8.61
+ $Y2=1.2
r132 30 43 3.70735 $w=2.5e-07 $l=1.75425e-07 $layer=LI1_cond $X=9.86 $Y=1.205
+ $X2=9.722 $Y2=1.12
r133 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.86 $Y=1.205
+ $X2=9.86 $Y2=1.875
r134 26 43 3.70735 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.665 $Y=1.035
+ $X2=9.722 $Y2=1.12
r135 26 28 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=9.665 $Y=1.035
+ $X2=9.665 $Y2=0.615
r136 24 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.775 $Y=1.96
+ $X2=9.86 $Y2=1.875
r137 24 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.775 $Y=1.96
+ $X2=9.48 $Y2=1.96
r138 23 41 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=9.395 $Y=2.445
+ $X2=9.395 $Y2=2.675
r139 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.395 $Y=2.045
+ $X2=9.48 $Y2=1.96
r140 22 23 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=9.395 $Y=2.045
+ $X2=9.395 $Y2=2.445
r141 21 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.775 $Y=1.12
+ $X2=8.61 $Y2=1.12
r142 20 43 2.76166 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=9.5 $Y=1.12
+ $X2=9.722 $Y2=1.12
r143 20 21 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=9.5 $Y=1.12
+ $X2=8.775 $Y2=1.12
r144 18 19 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=8.492 $Y=1.975
+ $X2=8.492 $Y2=2.125
r145 18 46 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.52 $Y=1.975
+ $X2=8.52 $Y2=1.365
r146 16 45 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=8.55 $Y=0.615
+ $X2=8.55 $Y2=1.035
r147 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.48 $Y=2.39 $X2=8.48
+ $Y2=2.675
r148 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.48 $Y=2.3 $X2=8.48
+ $Y2=2.39
r149 8 19 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=8.48 $Y=2.3
+ $X2=8.48 $Y2=2.125
r150 2 39 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=9.095
+ $Y=2.465 $X2=9.245 $Y2=2.675
r151 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.525
+ $Y=0.405 $X2=9.665 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_4%A_1350_392# 1 2 9 12 13 15 16 19 20 22 23 26
+ 27 29 31 34 35 36 37 38 39 40 43 45 50 51 52 58 59
c166 50 0 1.00633e-19 $X=8.325 $Y=2.475
c167 38 0 1.07146e-19 $X=10.475 $Y=1.335
c168 27 0 5.64102e-20 $X=10.425 $Y=1.97
c169 26 0 1.97399e-19 $X=10.425 $Y=1.88
r170 65 66 24.9528 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.51 $Y=1.63
+ $X2=9.51 $Y2=1.705
r171 59 65 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.51 $Y=1.54 $X2=9.51
+ $Y2=1.63
r172 59 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.51 $Y=1.54
+ $X2=9.51 $Y2=1.375
r173 58 61 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=9.475 $Y=1.54
+ $X2=9.475 $Y2=1.62
r174 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.51
+ $Y=1.54 $X2=9.51 $Y2=1.54
r175 51 61 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.345 $Y=1.62
+ $X2=9.475 $Y2=1.62
r176 51 52 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=9.345 $Y=1.62 $X2=8.41
+ $Y2=1.62
r177 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.325 $Y=1.705
+ $X2=8.41 $Y2=1.62
r178 49 50 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=8.325 $Y=1.705
+ $X2=8.325 $Y2=2.475
r179 46 54 2.79691 $w=3.3e-07 $l=1.03e-07 $layer=LI1_cond $X=7.33 $Y=2.64
+ $X2=7.227 $Y2=2.64
r180 46 48 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=7.33 $Y=2.64
+ $X2=7.835 $Y2=2.64
r181 45 50 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.24 $Y=2.64
+ $X2=8.325 $Y2=2.475
r182 45 48 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=8.24 $Y=2.64
+ $X2=7.835 $Y2=2.64
r183 41 56 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.33 $Y=0.72
+ $X2=7.245 $Y2=0.72
r184 41 43 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=7.33 $Y=0.72
+ $X2=7.77 $Y2=0.72
r185 40 54 4.96927 $w=1.7e-07 $l=1.73767e-07 $layer=LI1_cond $X=7.245 $Y=2.475
+ $X2=7.227 $Y2=2.64
r186 39 56 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.245 $Y=0.845
+ $X2=7.245 $Y2=0.72
r187 39 40 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=7.245 $Y=0.845
+ $X2=7.245 $Y2=2.475
r188 37 38 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=10.475 $Y=1.185
+ $X2=10.475 $Y2=1.335
r189 34 37 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=10.51 $Y=0.74
+ $X2=10.51 $Y2=1.185
r190 31 36 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=10.44 $Y=1.555
+ $X2=10.425 $Y2=1.63
r191 31 38 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=10.44 $Y=1.555
+ $X2=10.44 $Y2=1.335
r192 27 29 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.425 $Y=1.97
+ $X2=10.425 $Y2=2.465
r193 26 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.425 $Y=1.88
+ $X2=10.425 $Y2=1.97
r194 25 36 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=10.425 $Y=1.705
+ $X2=10.425 $Y2=1.63
r195 25 26 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=10.425 $Y=1.705
+ $X2=10.425 $Y2=1.88
r196 24 35 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.065 $Y=1.63
+ $X2=9.975 $Y2=1.63
r197 23 36 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.335 $Y=1.63
+ $X2=10.425 $Y2=1.63
r198 23 24 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=10.335 $Y=1.63
+ $X2=10.065 $Y2=1.63
r199 20 22 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.975 $Y=1.97
+ $X2=9.975 $Y2=2.465
r200 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.975 $Y=1.88
+ $X2=9.975 $Y2=1.97
r201 18 35 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.975 $Y=1.705
+ $X2=9.975 $Y2=1.63
r202 18 19 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=9.975 $Y=1.705
+ $X2=9.975 $Y2=1.88
r203 17 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.675 $Y=1.63
+ $X2=9.51 $Y2=1.63
r204 16 35 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.885 $Y=1.63
+ $X2=9.975 $Y2=1.63
r205 16 17 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.885 $Y=1.63
+ $X2=9.675 $Y2=1.63
r206 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.47 $Y=2.39
+ $X2=9.47 $Y2=2.675
r207 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.47 $Y=2.3 $X2=9.47
+ $Y2=2.39
r208 12 66 231.282 $w=1.8e-07 $l=5.95e-07 $layer=POLY_cond $X=9.47 $Y=2.3
+ $X2=9.47 $Y2=1.705
r209 9 64 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=9.45 $Y=0.615
+ $X2=9.45 $Y2=1.375
r210 2 54 600 $w=1.7e-07 $l=8.93868e-07 $layer=licon1_PDIFF $count=1 $X=6.75
+ $Y=1.96 $X2=7.245 $Y2=2.64
r211 2 48 600 $w=1.7e-07 $l=1.38384e-06 $layer=licon1_PDIFF $count=1 $X=6.75
+ $Y=1.96 $X2=7.835 $Y2=2.64
r212 1 56 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=7.185
+ $Y=0.37 $X2=7.325 $Y2=0.68
r213 1 43 182 $w=1.7e-07 $l=7.23585e-07 $layer=licon1_NDIFF $count=1 $X=7.185
+ $Y=0.37 $X2=7.77 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_4%A_2010_409# 1 2 7 9 10 12 14 17 19 20 23 25
+ 27 30 32 34 37 39 43 45 46 49 56 59 67
c131 23 0 1.38275e-19 $X=12.025 $Y=0.74
r132 61 62 9.0375 $w=4e-07 $l=7.5e-08 $layer=POLY_cond $X=11.425 $Y=1.532
+ $X2=11.5 $Y2=1.532
r133 57 65 54.5473 $w=2.43e-07 $l=2.75e-07 $layer=POLY_cond $X=12.075 $Y=1.532
+ $X2=12.35 $Y2=1.532
r134 57 63 9.9177 $w=2.43e-07 $l=5e-08 $layer=POLY_cond $X=12.075 $Y=1.532
+ $X2=12.025 $Y2=1.532
r135 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=12.075
+ $Y=1.465 $X2=12.075 $Y2=1.465
r136 54 61 3.615 $w=4e-07 $l=3e-08 $layer=POLY_cond $X=11.395 $Y=1.532
+ $X2=11.425 $Y2=1.532
r137 53 56 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=11.395 $Y=1.465
+ $X2=12.075 $Y2=1.465
r138 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=11.395
+ $Y=1.465 $X2=11.395 $Y2=1.465
r139 51 59 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=10.89 $Y=1.465
+ $X2=10.725 $Y2=1.465
r140 51 53 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=10.89 $Y=1.465
+ $X2=11.395 $Y2=1.465
r141 47 59 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.725 $Y=1.3
+ $X2=10.725 $Y2=1.465
r142 47 49 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=10.725 $Y=1.3
+ $X2=10.725 $Y2=0.515
r143 45 59 6.46576 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=10.56 $Y=1.545
+ $X2=10.725 $Y2=1.465
r144 45 46 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=10.56 $Y=1.545
+ $X2=10.365 $Y2=1.545
r145 41 46 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.24 $Y=1.63
+ $X2=10.365 $Y2=1.545
r146 41 43 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=10.24 $Y=1.63
+ $X2=10.24 $Y2=2.19
r147 35 67 30.7449 $w=2.43e-07 $l=1.55e-07 $layer=POLY_cond $X=12.955 $Y=1.532
+ $X2=12.8 $Y2=1.532
r148 35 37 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=12.955 $Y=1.48
+ $X2=12.955 $Y2=0.74
r149 32 67 14.0634 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=12.8 $Y=1.765
+ $X2=12.8 $Y2=1.532
r150 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.8 $Y=1.765
+ $X2=12.8 $Y2=2.4
r151 28 67 54.5473 $w=2.43e-07 $l=2.75e-07 $layer=POLY_cond $X=12.525 $Y=1.532
+ $X2=12.8 $Y2=1.532
r152 28 65 34.7119 $w=2.43e-07 $l=1.75e-07 $layer=POLY_cond $X=12.525 $Y=1.532
+ $X2=12.35 $Y2=1.532
r153 28 30 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=12.525 $Y=1.48
+ $X2=12.525 $Y2=0.74
r154 25 65 14.0634 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=12.35 $Y=1.765
+ $X2=12.35 $Y2=1.532
r155 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.35 $Y=1.765
+ $X2=12.35 $Y2=2.4
r156 21 63 14.0634 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=12.025 $Y=1.3
+ $X2=12.025 $Y2=1.532
r157 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=12.025 $Y=1.3
+ $X2=12.025 $Y2=0.74
r158 20 62 10.6563 $w=4e-07 $l=1.03199e-07 $layer=POLY_cond $X=11.575 $Y=1.465
+ $X2=11.5 $Y2=1.532
r159 19 63 14.4 $w=3.3e-07 $l=1.03199e-07 $layer=POLY_cond $X=11.95 $Y=1.465
+ $X2=12.025 $Y2=1.532
r160 19 20 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=11.95 $Y=1.465
+ $X2=11.575 $Y2=1.465
r161 15 62 25.8619 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=11.5 $Y=1.3
+ $X2=11.5 $Y2=1.532
r162 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.5 $Y=1.3
+ $X2=11.5 $Y2=0.74
r163 12 61 25.8619 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=11.425 $Y=1.765
+ $X2=11.425 $Y2=1.532
r164 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.425 $Y=1.765
+ $X2=11.425 $Y2=2.4
r165 11 39 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=11.02 $Y=1.555
+ $X2=10.93 $Y2=1.555
r166 10 54 39.5853 $w=4e-07 $l=1.76125e-07 $layer=POLY_cond $X=11.23 $Y=1.555
+ $X2=11.395 $Y2=1.532
r167 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=11.23 $Y=1.555
+ $X2=11.02 $Y2=1.555
r168 7 39 83.7788 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=10.93 $Y=1.765
+ $X2=10.93 $Y2=1.555
r169 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.93 $Y=1.765
+ $X2=10.93 $Y2=2.4
r170 2 43 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=10.05
+ $Y=2.045 $X2=10.2 $Y2=2.19
r171 1 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.585
+ $Y=0.37 $X2=10.725 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 31 33 37 41 45 49
+ 53 57 61 65 67 69 74 75 77 78 80 81 82 84 89 94 102 120 124 133 136 139 142
+ 145 149
c172 149 0 2.33512e-20 $X=13.2 $Y=3.33
c173 102 0 1.50343e-19 $X=5.83 $Y=3.33
c174 84 0 1.97046e-19 $X=1 $Y=3.33
c175 61 0 1.07146e-19 $X=10.7 $Y=2.19
r176 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r177 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r178 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r179 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r180 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r181 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r182 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r183 128 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r184 128 146 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=11.76 $Y2=3.33
r185 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r186 125 145 13.7128 $w=1.7e-07 $l=3.53e-07 $layer=LI1_cond $X=12.24 $Y=3.33
+ $X2=11.887 $Y2=3.33
r187 125 127 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r188 124 148 4.57341 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=12.91 $Y=3.33
+ $X2=13.175 $Y2=3.33
r189 124 127 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=12.91 $Y=3.33
+ $X2=12.72 $Y2=3.33
r190 123 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r191 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r192 120 145 13.7128 $w=1.7e-07 $l=3.52e-07 $layer=LI1_cond $X=11.535 $Y=3.33
+ $X2=11.887 $Y2=3.33
r193 120 122 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.535 $Y=3.33
+ $X2=11.28 $Y2=3.33
r194 119 123 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r195 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r196 116 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r197 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r198 113 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r199 112 113 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r200 110 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r201 109 112 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=8.4 $Y2=3.33
r202 109 110 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r203 107 142 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=5.997 $Y2=3.33
r204 107 109 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=6.48 $Y2=3.33
r205 106 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r206 106 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r207 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r208 103 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=4.565 $Y2=3.33
r209 103 105 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=5.52 $Y2=3.33
r210 102 142 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=5.83 $Y=3.33
+ $X2=5.997 $Y2=3.33
r211 102 105 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.83 $Y=3.33
+ $X2=5.52 $Y2=3.33
r212 101 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r213 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r214 98 101 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r215 98 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r216 97 100 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r217 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r218 95 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.17 $Y2=3.33
r219 95 97 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.64 $Y2=3.33
r220 94 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=3.33
+ $X2=4.565 $Y2=3.33
r221 94 100 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.4 $Y=3.33
+ $X2=4.08 $Y2=3.33
r222 93 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r223 93 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r224 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r225 90 133 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.34 $Y=3.33
+ $X2=1.17 $Y2=3.33
r226 90 92 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.34 $Y=3.33
+ $X2=1.68 $Y2=3.33
r227 89 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=3.33
+ $X2=2.17 $Y2=3.33
r228 89 92 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.005 $Y=3.33
+ $X2=1.68 $Y2=3.33
r229 88 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r230 88 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r231 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r232 85 130 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=3.33
+ $X2=0.18 $Y2=3.33
r233 85 87 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.36 $Y=3.33
+ $X2=0.72 $Y2=3.33
r234 84 133 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1 $Y=3.33 $X2=1.17
+ $Y2=3.33
r235 84 87 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1 $Y=3.33 $X2=0.72
+ $Y2=3.33
r236 82 113 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=8.4 $Y2=3.33
r237 82 110 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.48 $Y2=3.33
r238 80 118 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.535 $Y=3.33
+ $X2=10.32 $Y2=3.33
r239 80 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.535 $Y=3.33
+ $X2=10.7 $Y2=3.33
r240 79 122 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=10.865 $Y=3.33
+ $X2=11.28 $Y2=3.33
r241 79 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.865 $Y=3.33
+ $X2=10.7 $Y2=3.33
r242 77 115 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=9.65 $Y=3.33
+ $X2=9.36 $Y2=3.33
r243 77 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.65 $Y=3.33
+ $X2=9.775 $Y2=3.33
r244 76 118 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.9 $Y=3.33
+ $X2=10.32 $Y2=3.33
r245 76 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.9 $Y=3.33
+ $X2=9.775 $Y2=3.33
r246 74 112 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.58 $Y=3.33
+ $X2=8.4 $Y2=3.33
r247 74 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.58 $Y=3.33
+ $X2=8.745 $Y2=3.33
r248 73 115 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.91 $Y=3.33
+ $X2=9.36 $Y2=3.33
r249 73 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.91 $Y=3.33
+ $X2=8.745 $Y2=3.33
r250 69 72 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=13.075 $Y=2.115
+ $X2=13.075 $Y2=2.815
r251 67 148 3.19276 $w=3.3e-07 $l=1.36015e-07 $layer=LI1_cond $X=13.075 $Y=3.245
+ $X2=13.175 $Y2=3.33
r252 67 72 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.075 $Y=3.245
+ $X2=13.075 $Y2=2.815
r253 63 145 2.87722 $w=7.05e-07 $l=8.5e-08 $layer=LI1_cond $X=11.887 $Y=3.245
+ $X2=11.887 $Y2=3.33
r254 63 65 15.9477 $w=7.03e-07 $l=9.4e-07 $layer=LI1_cond $X=11.887 $Y=3.245
+ $X2=11.887 $Y2=2.305
r255 59 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.7 $Y=3.245
+ $X2=10.7 $Y2=3.33
r256 59 61 36.8433 $w=3.28e-07 $l=1.055e-06 $layer=LI1_cond $X=10.7 $Y=3.245
+ $X2=10.7 $Y2=2.19
r257 55 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=3.245
+ $X2=9.775 $Y2=3.33
r258 55 57 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=9.775 $Y=3.245
+ $X2=9.775 $Y2=2.675
r259 51 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.745 $Y=3.245
+ $X2=8.745 $Y2=3.33
r260 51 53 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=8.745 $Y=3.245
+ $X2=8.745 $Y2=2.675
r261 47 142 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=5.997 $Y=3.245
+ $X2=5.997 $Y2=3.33
r262 47 49 14.2765 $w=3.33e-07 $l=4.15e-07 $layer=LI1_cond $X=5.997 $Y=3.245
+ $X2=5.997 $Y2=2.83
r263 43 139 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=3.245
+ $X2=4.565 $Y2=3.33
r264 43 45 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.565 $Y=3.245
+ $X2=4.565 $Y2=2.825
r265 39 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=3.33
r266 39 41 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=2.835
r267 35 133 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r268 35 37 13.8971 $w=3.38e-07 $l=4.1e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.835
r269 31 130 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.235 $Y=3.245
+ $X2=0.18 $Y2=3.33
r270 31 33 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.235 $Y=3.245
+ $X2=0.235 $Y2=2.75
r271 10 72 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=12.875
+ $Y=1.84 $X2=13.075 $Y2=2.815
r272 10 69 400 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=12.875
+ $Y=1.84 $X2=13.075 $Y2=2.115
r273 9 65 150 $w=1.7e-07 $l=8.20183e-07 $layer=licon1_PDIFF $count=4 $X=11.5
+ $Y=1.84 $X2=12.12 $Y2=2.305
r274 8 61 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=10.5
+ $Y=2.045 $X2=10.7 $Y2=2.19
r275 7 57 600 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_PDIFF $count=1 $X=9.545
+ $Y=2.465 $X2=9.735 $Y2=2.675
r276 6 53 600 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_PDIFF $count=1 $X=8.555
+ $Y=2.465 $X2=8.745 $Y2=2.675
r277 5 49 600 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_PDIFF $count=1 $X=5.81
+ $Y=2.7 $X2=5.995 $Y2=2.83
r278 4 45 600 $w=1.7e-07 $l=6.14329e-07 $layer=licon1_PDIFF $count=1 $X=4.335
+ $Y=2.315 $X2=4.565 $Y2=2.825
r279 3 41 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=2.02
+ $Y=1.96 $X2=2.17 $Y2=2.835
r280 2 37 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=2.54 $X2=1.165 $Y2=2.835
r281 1 33 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.275 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_4%A_37_78# 1 2 3 4 13 17 20 21 25 27 29 30 32
+ 34 38 40
c118 40 0 3.12839e-20 $X=3.17 $Y=2.495
c119 38 0 1.97046e-19 $X=0.56 $Y=2.52
c120 30 0 1.94359e-19 $X=3.435 $Y=1.305
c121 29 0 4.38676e-20 $X=3.625 $Y=1.305
r122 40 42 1.47581 $w=2.48e-07 $l=3e-08 $layer=LI1_cond $X=3.17 $Y=2.495
+ $X2=3.17 $Y2=2.525
r123 39 40 11.0685 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=3.17 $Y=2.27
+ $X2=3.17 $Y2=2.495
r124 34 36 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.33 $Y=0.6
+ $X2=0.33 $Y2=0.745
r125 31 32 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=3.71 $Y=1.39
+ $X2=3.71 $Y2=2.185
r126 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.625 $Y=1.305
+ $X2=3.71 $Y2=1.39
r127 29 30 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.625 $Y=1.305
+ $X2=3.435 $Y2=1.305
r128 28 39 2.94836 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.31 $Y=2.27
+ $X2=3.17 $Y2=2.27
r129 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.625 $Y=2.27
+ $X2=3.71 $Y2=2.185
r130 27 28 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.625 $Y=2.27
+ $X2=3.31 $Y2=2.27
r131 23 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.31 $Y=1.22
+ $X2=3.435 $Y2=1.305
r132 23 25 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=3.31 $Y=1.22
+ $X2=3.31 $Y2=0.9
r133 22 38 2.28545 $w=1.7e-07 $l=3.42272e-07 $layer=LI1_cond $X=0.89 $Y=2.495
+ $X2=0.56 $Y2=2.52
r134 21 40 2.94836 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.03 $Y=2.495
+ $X2=3.17 $Y2=2.495
r135 21 22 139.615 $w=1.68e-07 $l=2.14e-06 $layer=LI1_cond $X=3.03 $Y=2.495
+ $X2=0.89 $Y2=2.495
r136 20 38 4.14756 $w=2.2e-07 $l=2.5923e-07 $layer=LI1_cond $X=0.77 $Y=2.41
+ $X2=0.56 $Y2=2.52
r137 19 20 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=0.77 $Y=0.83
+ $X2=0.77 $Y2=2.41
r138 15 38 4.14756 $w=2.2e-07 $l=1.8554e-07 $layer=LI1_cond $X=0.695 $Y=2.64
+ $X2=0.56 $Y2=2.52
r139 15 17 4.69514 $w=2.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.695 $Y=2.64
+ $X2=0.695 $Y2=2.75
r140 14 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.495 $Y=0.745
+ $X2=0.33 $Y2=0.745
r141 13 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=0.745
+ $X2=0.77 $Y2=0.83
r142 13 14 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.685 $Y=0.745
+ $X2=0.495 $Y2=0.745
r143 4 42 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.055
+ $Y=2.315 $X2=3.195 $Y2=2.525
r144 3 17 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=2.54 $X2=0.725 $Y2=2.75
r145 2 25 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.135
+ $Y=0.69 $X2=3.27 $Y2=0.9
r146 1 34 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.39 $X2=0.33 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_4%Q 1 2 3 4 15 19 20 21 23 25 29 35 38 41 42
c73 42 0 1.38275e-19 $X=13.2 $Y=1.665
r74 44 45 2.94971 $w=5.17e-07 $l=1.25e-07 $layer=LI1_cond $X=12.575 $Y=1.62
+ $X2=12.7 $Y2=1.62
r75 42 45 11.7988 $w=5.17e-07 $l=5e-07 $layer=LI1_cond $X=13.2 $Y=1.62 $X2=12.7
+ $Y2=1.62
r76 38 45 5.00057 $w=2.5e-07 $l=3.5e-07 $layer=LI1_cond $X=12.7 $Y=1.27 $X2=12.7
+ $Y2=1.62
r77 37 41 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=12.7 $Y=1.13
+ $X2=12.7 $Y2=1.005
r78 37 38 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=12.7 $Y=1.13
+ $X2=12.7 $Y2=1.27
r79 33 41 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=12.7 $Y=0.88
+ $X2=12.7 $Y2=1.005
r80 33 35 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=12.7 $Y=0.88
+ $X2=12.7 $Y2=0.515
r81 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=12.575 $Y=1.985
+ $X2=12.575 $Y2=2.815
r82 27 44 3.36414 $w=3.3e-07 $l=3.5e-07 $layer=LI1_cond $X=12.575 $Y=1.97
+ $X2=12.575 $Y2=1.62
r83 27 29 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=12.575 $Y=1.97
+ $X2=12.575 $Y2=1.985
r84 26 40 3.87155 $w=2.5e-07 $l=1.58e-07 $layer=LI1_cond $X=11.91 $Y=1.005
+ $X2=11.752 $Y2=1.005
r85 25 41 1.34256 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=12.575 $Y=1.005
+ $X2=12.7 $Y2=1.005
r86 25 26 30.655 $w=2.48e-07 $l=6.65e-07 $layer=LI1_cond $X=12.575 $Y=1.005
+ $X2=11.91 $Y2=1.005
r87 21 40 3.06294 $w=3.15e-07 $l=1.25e-07 $layer=LI1_cond $X=11.752 $Y=0.88
+ $X2=11.752 $Y2=1.005
r88 21 23 12.8049 $w=3.13e-07 $l=3.5e-07 $layer=LI1_cond $X=11.752 $Y=0.88
+ $X2=11.752 $Y2=0.53
r89 19 44 9.81494 $w=5.17e-07 $l=3.37565e-07 $layer=LI1_cond $X=12.41 $Y=1.885
+ $X2=12.575 $Y2=1.62
r90 19 20 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=12.41 $Y=1.885
+ $X2=11.365 $Y2=1.885
r91 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=11.2 $Y=1.985
+ $X2=11.2 $Y2=2.815
r92 13 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.2 $Y=1.97
+ $X2=11.365 $Y2=1.885
r93 13 15 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=11.2 $Y=1.97
+ $X2=11.2 $Y2=1.985
r94 4 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12.425
+ $Y=1.84 $X2=12.575 $Y2=2.815
r95 4 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.425
+ $Y=1.84 $X2=12.575 $Y2=1.985
r96 3 17 400 $w=1.7e-07 $l=1.06806e-06 $layer=licon1_PDIFF $count=1 $X=11.005
+ $Y=1.84 $X2=11.2 $Y2=2.815
r97 3 15 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=11.005
+ $Y=1.84 $X2=11.2 $Y2=1.985
r98 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.6
+ $Y=0.37 $X2=12.74 $Y2=0.515
r99 1 40 182 $w=1.7e-07 $l=6.81249e-07 $layer=licon1_NDIFF $count=1 $X=11.575
+ $Y=0.37 $X2=11.76 $Y2=0.965
r100 1 23 182 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=1 $X=11.575
+ $Y=0.37 $X2=11.76 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LS__DFRTP_4%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 49 51
+ 54 55 57 58 59 65 69 77 89 93 98 104 108 114 117 120 124
c141 124 0 6.43803e-21 $X=13.2 $Y=0
r142 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r143 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r144 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r145 114 115 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r146 108 111 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.06 $Y=0
+ $X2=5.06 $Y2=0.285
r147 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r148 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r149 102 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r150 102 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r151 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r152 99 120 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=12.405 $Y=0
+ $X2=12.242 $Y2=0
r153 99 101 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.405 $Y=0
+ $X2=12.72 $Y2=0
r154 98 123 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=13.005 $Y=0
+ $X2=13.222 $Y2=0
r155 98 101 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.005 $Y=0
+ $X2=12.72 $Y2=0
r156 97 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r157 97 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r158 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r159 94 117 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.41 $Y=0
+ $X2=11.265 $Y2=0
r160 94 96 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=11.41 $Y=0
+ $X2=11.76 $Y2=0
r161 93 120 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=12.08 $Y=0
+ $X2=12.242 $Y2=0
r162 93 96 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=12.08 $Y=0 $X2=11.76
+ $Y2=0
r163 92 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r164 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r165 89 117 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.12 $Y=0
+ $X2=11.265 $Y2=0
r166 89 91 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=11.12 $Y=0 $X2=10.8
+ $Y2=0
r167 88 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=10.8
+ $Y2=0
r168 88 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=8.88 $Y2=0
r169 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r170 85 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.955 $Y=0
+ $X2=8.79 $Y2=0
r171 85 87 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=8.955 $Y=0 $X2=9.84
+ $Y2=0
r172 84 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r173 83 84 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r174 81 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r175 80 83 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=8.4
+ $Y2=0
r176 80 81 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r177 78 108 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.225 $Y=0
+ $X2=5.06 $Y2=0
r178 78 80 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.225 $Y=0 $X2=5.52
+ $Y2=0
r179 77 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.625 $Y=0
+ $X2=8.79 $Y2=0
r180 77 83 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.625 $Y=0 $X2=8.4
+ $Y2=0
r181 76 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r182 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r183 73 76 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r184 73 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r185 72 75 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r186 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r187 70 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.385 $Y=0
+ $X2=2.22 $Y2=0
r188 70 72 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.385 $Y=0
+ $X2=2.64 $Y2=0
r189 69 108 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.895 $Y=0
+ $X2=5.06 $Y2=0
r190 69 75 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.895 $Y=0
+ $X2=4.56 $Y2=0
r191 68 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r192 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r193 65 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.055 $Y=0
+ $X2=2.22 $Y2=0
r194 65 67 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.055 $Y=0
+ $X2=1.68 $Y2=0
r195 63 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r196 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r197 59 84 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=0 $X2=8.4
+ $Y2=0
r198 59 81 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=6.72 $Y=0 $X2=5.52
+ $Y2=0
r199 57 87 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=9.84 $Y2=0
r200 57 58 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=10.252 $Y2=0
r201 56 91 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=10.39 $Y=0 $X2=10.8
+ $Y2=0
r202 56 58 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=10.39 $Y=0
+ $X2=10.252 $Y2=0
r203 54 62 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.72
+ $Y2=0
r204 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.15
+ $Y2=0
r205 53 67 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.235 $Y=0
+ $X2=1.68 $Y2=0
r206 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.15
+ $Y2=0
r207 49 123 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=13.17 $Y=0.085
+ $X2=13.222 $Y2=0
r208 49 51 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.17 $Y=0.085
+ $X2=13.17 $Y2=0.515
r209 45 120 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=12.242 $Y=0.085
+ $X2=12.242 $Y2=0
r210 45 47 15.7796 $w=3.23e-07 $l=4.45e-07 $layer=LI1_cond $X=12.242 $Y=0.085
+ $X2=12.242 $Y2=0.53
r211 41 117 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=11.265 $Y=0.085
+ $X2=11.265 $Y2=0
r212 41 43 17.684 $w=2.88e-07 $l=4.45e-07 $layer=LI1_cond $X=11.265 $Y=0.085
+ $X2=11.265 $Y2=0.53
r213 37 58 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=10.252 $Y=0.085
+ $X2=10.252 $Y2=0
r214 37 39 18.02 $w=2.73e-07 $l=4.3e-07 $layer=LI1_cond $X=10.252 $Y=0.085
+ $X2=10.252 $Y2=0.515
r215 33 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.79 $Y=0.085
+ $X2=8.79 $Y2=0
r216 33 35 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=8.79 $Y=0.085
+ $X2=8.79 $Y2=0.615
r217 29 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=0.085
+ $X2=2.22 $Y2=0
r218 29 31 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=2.22 $Y=0.085
+ $X2=2.22 $Y2=0.715
r219 25 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0
r220 25 27 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0.6
r221 8 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.03
+ $Y=0.37 $X2=13.17 $Y2=0.515
r222 7 47 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=12.1
+ $Y=0.37 $X2=12.24 $Y2=0.53
r223 6 43 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=11.14
+ $Y=0.37 $X2=11.285 $Y2=0.53
r224 5 39 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.08
+ $Y=0.37 $X2=10.225 $Y2=0.515
r225 4 35 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=8.625
+ $Y=0.405 $X2=8.79 $Y2=0.615
r226 3 111 182 $w=1.7e-07 $l=5.03115e-07 $layer=licon1_NDIFF $count=1 $X=4.84
+ $Y=0.69 $X2=5.06 $Y2=0.285
r227 2 31 182 $w=1.7e-07 $l=2.32379e-07 $layer=licon1_NDIFF $count=1 $X=2.04
+ $Y=0.595 $X2=2.22 $Y2=0.715
r228 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.39 $X2=1.15 $Y2=0.6
.ends

