* File: sky130_fd_sc_ls__a311o_2.pex.spice
* Created: Fri Aug 28 12:57:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A311O_2%A_21_270# 1 2 3 10 12 15 17 18 20 21 23 26
+ 28 31 34 37 38 40 41 42 43 47 49 51 53 57 59 62
c149 21 0 1.22049e-19 $X=1.055 $Y=1.765
r150 59 60 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.25 $Y=2.035
+ $X2=1.25 $Y2=2.315
r151 55 57 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=3.875 $Y=0.92
+ $X2=3.875 $Y2=0.515
r152 51 64 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=2.12 $X2=3.87
+ $Y2=2.035
r153 51 53 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.87 $Y=2.12
+ $X2=3.87 $Y2=2.815
r154 50 62 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3 $Y=1.005
+ $X2=2.815 $Y2=1.005
r155 49 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.71 $Y=1.005
+ $X2=3.875 $Y2=0.92
r156 49 50 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.71 $Y=1.005 $X2=3
+ $Y2=1.005
r157 45 62 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.815 $Y=0.92
+ $X2=2.815 $Y2=1.005
r158 45 47 12.6146 $w=3.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.815 $Y=0.92
+ $X2=2.815 $Y2=0.515
r159 44 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.335 $Y=2.035
+ $X2=1.25 $Y2=2.035
r160 43 64 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=2.035
+ $X2=3.87 $Y2=2.035
r161 43 44 154.62 $w=1.68e-07 $l=2.37e-06 $layer=LI1_cond $X=3.705 $Y=2.035
+ $X2=1.335 $Y2=2.035
r162 41 62 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.63 $Y=1.005
+ $X2=2.815 $Y2=1.005
r163 41 42 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=2.63 $Y=1.005
+ $X2=1.335 $Y2=1.005
r164 40 59 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=1.95
+ $X2=1.25 $Y2=2.035
r165 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.25 $Y=1.09
+ $X2=1.335 $Y2=1.005
r166 39 40 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.25 $Y=1.09
+ $X2=1.25 $Y2=1.95
r167 37 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=2.315
+ $X2=1.25 $Y2=2.315
r168 37 38 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.165 $Y=2.315
+ $X2=0.435 $Y2=2.315
r169 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.515 $X2=0.27 $Y2=1.515
r170 32 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.27 $Y=2.23
+ $X2=0.435 $Y2=2.315
r171 32 34 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=0.27 $Y=2.23
+ $X2=0.27 $Y2=1.515
r172 29 30 9.19847 $w=3.93e-07 $l=7.5e-08 $layer=POLY_cond $X=0.605 $Y=1.557
+ $X2=0.68 $Y2=1.557
r173 28 35 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=0.515 $Y=1.515
+ $X2=0.27 $Y2=1.515
r174 28 29 12.4178 $w=3.93e-07 $l=1.08995e-07 $layer=POLY_cond $X=0.515 $Y=1.515
+ $X2=0.605 $Y2=1.557
r175 24 31 18.8402 $w=1.65e-07 $l=9.08295e-08 $layer=POLY_cond $X=1.11 $Y=1.35
+ $X2=1.075 $Y2=1.425
r176 24 26 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.11 $Y=1.35
+ $X2=1.11 $Y2=0.74
r177 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.055 $Y=1.765
+ $X2=1.055 $Y2=2.4
r178 20 21 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.055 $Y=1.675
+ $X2=1.055 $Y2=1.765
r179 19 31 18.8402 $w=1.65e-07 $l=8.44097e-08 $layer=POLY_cond $X=1.055 $Y=1.5
+ $X2=1.075 $Y2=1.425
r180 19 20 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=1.055 $Y=1.5
+ $X2=1.055 $Y2=1.675
r181 18 30 28.4128 $w=3.93e-07 $l=1.653e-07 $layer=POLY_cond $X=0.755 $Y=1.425
+ $X2=0.68 $Y2=1.557
r182 17 31 6.66866 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=0.965 $Y=1.425
+ $X2=1.075 $Y2=1.425
r183 17 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.965 $Y=1.425
+ $X2=0.755 $Y2=1.425
r184 13 30 25.4309 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.68 $Y=1.35
+ $X2=0.68 $Y2=1.557
r185 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.68 $Y=1.35
+ $X2=0.68 $Y2=0.74
r186 10 29 25.4309 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.605 $Y=1.765
+ $X2=0.605 $Y2=1.557
r187 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.605 $Y=1.765
+ $X2=0.605 $Y2=2.4
r188 3 64 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=3.72
+ $Y=1.96 $X2=3.87 $Y2=2.115
r189 3 53 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.72
+ $Y=1.96 $X2=3.87 $Y2=2.815
r190 2 57 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.735
+ $Y=0.37 $X2=3.875 $Y2=0.515
r191 1 47 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=2.655
+ $Y=0.37 $X2=2.815 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_2%A3 2 3 5 8 10 13 14
c40 13 0 1.61501e-19 $X=1.59 $Y=1.425
c41 8 0 9.80412e-20 $X=1.68 $Y=0.74
c42 2 0 1.95903e-19 $X=1.575 $Y=1.795
r43 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.425
+ $X2=1.59 $Y2=1.59
r44 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.425
+ $X2=1.59 $Y2=1.26
r45 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.59
+ $Y=1.425 $X2=1.59 $Y2=1.425
r46 10 14 9.53746 $w=2.88e-07 $l=2.4e-07 $layer=LI1_cond $X=1.65 $Y=1.665
+ $X2=1.65 $Y2=1.425
r47 8 15 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.68 $Y=0.74 $X2=1.68
+ $Y2=1.26
r48 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.575 $Y=1.885
+ $X2=1.575 $Y2=2.46
r49 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.575 $Y=1.795 $X2=1.575
+ $Y2=1.885
r50 2 16 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=1.575 $Y=1.795
+ $X2=1.575 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_2%A2 3 5 7 8
c30 8 0 3.57404e-19 $X=2.16 $Y=1.665
r31 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.615 $X2=2.13 $Y2=1.615
r32 5 11 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=2.055 $Y=1.885
+ $X2=2.13 $Y2=1.615
r33 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.055 $Y=1.885
+ $X2=2.055 $Y2=2.46
r34 1 11 38.5916 $w=2.93e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.04 $Y=1.45
+ $X2=2.13 $Y2=1.615
r35 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.04 $Y=1.45 $X2=2.04
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_2%A1 3 5 7 8
c33 8 0 3.55573e-19 $X=2.64 $Y=1.665
r34 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.615 $X2=2.67 $Y2=1.615
r35 5 11 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=2.745 $Y=1.885
+ $X2=2.67 $Y2=1.615
r36 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.745 $Y=1.885
+ $X2=2.745 $Y2=2.46
r37 1 11 38.5916 $w=2.93e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.58 $Y=1.45
+ $X2=2.67 $Y2=1.615
r38 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.58 $Y=1.45 $X2=2.58
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_2%B1 3 6 7 9 10 11 15
c38 15 0 2.32531e-19 $X=3.21 $Y=1.425
c39 6 0 2.78177e-19 $X=3.225 $Y=1.795
r40 15 18 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.425
+ $X2=3.21 $Y2=1.59
r41 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.425
+ $X2=3.21 $Y2=1.26
r42 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.21
+ $Y=1.425 $X2=3.21 $Y2=1.425
r43 11 16 8.97059 $w=5.18e-07 $l=3.9e-07 $layer=LI1_cond $X=3.6 $Y=1.52 $X2=3.21
+ $Y2=1.52
r44 10 16 2.07014 $w=5.18e-07 $l=9e-08 $layer=LI1_cond $X=3.12 $Y=1.52 $X2=3.21
+ $Y2=1.52
r45 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.225 $Y=1.885
+ $X2=3.225 $Y2=2.46
r46 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.225 $Y=1.795 $X2=3.225
+ $Y2=1.885
r47 6 18 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=3.225 $Y=1.795
+ $X2=3.225 $Y2=1.59
r48 3 17 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=3.12 $Y=0.74 $X2=3.12
+ $Y2=1.26
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_2%C1 1 3 6 9 10 13
c33 10 0 1.55135e-19 $X=4.08 $Y=1.665
r34 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.605 $X2=4.05 $Y2=1.605
r35 8 13 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=3.735 $Y=1.605
+ $X2=4.05 $Y2=1.605
r36 8 9 5.03009 $w=3.3e-07 $l=2.24499e-07 $layer=POLY_cond $X=3.735 $Y=1.605
+ $X2=3.555 $Y2=1.705
r37 4 9 37.0704 $w=1.5e-07 $l=3.13129e-07 $layer=POLY_cond $X=3.66 $Y=1.44
+ $X2=3.555 $Y2=1.705
r38 4 6 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=3.66 $Y=1.44 $X2=3.66
+ $Y2=0.74
r39 1 9 37.0704 $w=1.5e-07 $l=2.20454e-07 $layer=POLY_cond $X=3.645 $Y=1.885
+ $X2=3.555 $Y2=1.705
r40 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.645 $Y=1.885
+ $X2=3.645 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_2%VPWR 1 2 3 10 12 16 18 20 22 29 30 36 39
r57 42 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 39 42 11.3966 $w=5.28e-07 $l=5.05e-07 $layer=LI1_cond $X=2.4 $Y=2.825
+ $X2=2.4 $Y2=3.33
r59 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r60 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 30 45 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r62 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r63 27 42 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=2.665 $Y=3.33
+ $X2=2.4 $Y2=3.33
r64 27 29 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=2.665 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r66 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r67 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 23 33 4.54971 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=0.545 $Y=3.33
+ $X2=0.272 $Y2=3.33
r69 23 25 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.545 $Y=3.33
+ $X2=0.72 $Y2=3.33
r70 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.28 $Y2=3.33
r71 22 25 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 20 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r73 20 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r74 20 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r75 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.28 $Y2=3.33
r76 18 42 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=2.135 $Y=3.33
+ $X2=2.4 $Y2=3.33
r77 18 19 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.135 $Y=3.33
+ $X2=1.445 $Y2=3.33
r78 14 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=3.245
+ $X2=1.28 $Y2=3.33
r79 14 16 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.28 $Y=3.245
+ $X2=1.28 $Y2=2.735
r80 10 33 3.21646 $w=3.3e-07 $l=1.44375e-07 $layer=LI1_cond $X=0.38 $Y=3.245
+ $X2=0.272 $Y2=3.33
r81 10 12 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.38 $Y=3.245
+ $X2=0.38 $Y2=2.735
r82 3 39 600 $w=1.7e-07 $l=9.90846e-07 $layer=licon1_PDIFF $count=1 $X=2.13
+ $Y=1.96 $X2=2.4 $Y2=2.825
r83 2 16 600 $w=1.7e-07 $l=9.67096e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.84 $X2=1.28 $Y2=2.735
r84 1 12 600 $w=1.7e-07 $l=9.55458e-07 $layer=licon1_PDIFF $count=1 $X=0.255
+ $Y=1.84 $X2=0.38 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_2%X 1 2 10 12 15
c23 12 0 9.80412e-20 $X=0.895 $Y=0.495
r24 15 21 9.16044 $w=3.88e-07 $l=3.1e-07 $layer=LI1_cond $X=0.8 $Y=1.665 $X2=0.8
+ $Y2=1.975
r25 15 18 4.58901 $w=3.88e-07 $l=1.15e-07 $layer=LI1_cond $X=0.8 $Y=1.665
+ $X2=0.8 $Y2=1.55
r26 12 14 9.38574 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0.495
+ $X2=0.895 $Y2=0.75
r27 10 18 24.571 $w=2.63e-07 $l=5.65e-07 $layer=LI1_cond $X=0.862 $Y=0.985
+ $X2=0.862 $Y2=1.55
r28 10 14 10.2198 $w=2.63e-07 $l=2.35e-07 $layer=LI1_cond $X=0.862 $Y=0.985
+ $X2=0.862 $Y2=0.75
r29 2 21 600 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=0.68
+ $Y=1.84 $X2=0.83 $Y2=1.975
r30 1 12 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.755
+ $Y=0.37 $X2=0.895 $Y2=0.495
r31 1 10 182 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_NDIFF $count=1 $X=0.755
+ $Y=0.37 $X2=0.895 $Y2=0.985
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_2%A_330_392# 1 2 7 9 11 13 15
c33 9 0 1.22049e-19 $X=1.8 $Y=2.835
r34 13 20 3.1563 $w=3.3e-07 $l=1.4e-07 $layer=LI1_cond $X=3 $Y=2.57 $X2=3
+ $Y2=2.43
r35 13 15 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3 $Y=2.57 $X2=3
+ $Y2=2.835
r36 12 18 3.71993 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=2.43
+ $X2=1.8 $Y2=2.43
r37 11 20 3.71993 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=2.43 $X2=3
+ $Y2=2.43
r38 11 12 35.8081 $w=2.78e-07 $l=8.7e-07 $layer=LI1_cond $X=2.835 $Y=2.43
+ $X2=1.965 $Y2=2.43
r39 7 18 3.1563 $w=3.3e-07 $l=1.4e-07 $layer=LI1_cond $X=1.8 $Y=2.57 $X2=1.8
+ $Y2=2.43
r40 7 9 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.8 $Y=2.57 $X2=1.8
+ $Y2=2.835
r41 2 20 600 $w=1.7e-07 $l=5.27376e-07 $layer=licon1_PDIFF $count=1 $X=2.82
+ $Y=1.96 $X2=3 $Y2=2.405
r42 2 15 600 $w=1.7e-07 $l=9.60794e-07 $layer=licon1_PDIFF $count=1 $X=2.82
+ $Y=1.96 $X2=3 $Y2=2.835
r43 1 18 600 $w=1.7e-07 $l=5.14563e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=1.96 $X2=1.8 $Y2=2.405
r44 1 9 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=1.96 $X2=1.8 $Y2=2.835
.ends

.subckt PM_SKY130_FD_SC_LS__A311O_2%VGND 1 2 3 12 16 20 23 24 26 27 29 30 31 46
+ 47
r51 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r52 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r53 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r54 40 43 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r55 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r56 38 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r57 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r58 35 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r59 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r60 31 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r61 31 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r62 29 43 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.17 $Y=0 $X2=3.12
+ $Y2=0
r63 29 30 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.17 $Y=0 $X2=3.355
+ $Y2=0
r64 28 46 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.54 $Y=0 $X2=4.08
+ $Y2=0
r65 28 30 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.54 $Y=0 $X2=3.355
+ $Y2=0
r66 26 37 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.23 $Y=0 $X2=1.2
+ $Y2=0
r67 26 27 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.23 $Y=0 $X2=1.43
+ $Y2=0
r68 25 40 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.63 $Y=0 $X2=1.68
+ $Y2=0
r69 25 27 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.63 $Y=0 $X2=1.43
+ $Y2=0
r70 23 34 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=0.3 $Y=0 $X2=0.24 $Y2=0
r71 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.3 $Y=0 $X2=0.425
+ $Y2=0
r72 22 37 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=1.2
+ $Y2=0
r73 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.425
+ $Y2=0
r74 18 30 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=0.085
+ $X2=3.355 $Y2=0
r75 18 20 15.5736 $w=3.68e-07 $l=5e-07 $layer=LI1_cond $X=3.355 $Y=0.085
+ $X2=3.355 $Y2=0.585
r76 14 27 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.43 $Y=0.085 $X2=1.43
+ $Y2=0
r77 14 16 14.4055 $w=3.98e-07 $l=5e-07 $layer=LI1_cond $X=1.43 $Y=0.085 $X2=1.43
+ $Y2=0.585
r78 10 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.425 $Y=0.085
+ $X2=0.425 $Y2=0
r79 10 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.425 $Y=0.085
+ $X2=0.425 $Y2=0.515
r80 3 20 182 $w=1.7e-07 $l=2.83945e-07 $layer=licon1_NDIFF $count=1 $X=3.195
+ $Y=0.37 $X2=3.355 $Y2=0.585
r81 2 16 182 $w=1.7e-07 $l=3.35708e-07 $layer=licon1_NDIFF $count=1 $X=1.185
+ $Y=0.37 $X2=1.43 $Y2=0.585
r82 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.34
+ $Y=0.37 $X2=0.465 $Y2=0.515
.ends

