* File: sky130_fd_sc_ls__dfrtp_4.spice
* Created: Wed Sep  2 11:01:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dfrtp_4.pex.spice"
.subckt sky130_fd_sc_ls__dfrtp_4  VNB VPB D CLK RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1012 A_124_78# N_D_M1012_g N_A_37_78#_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_RESET_B_M1002_g A_124_78# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_CLK_M1008_g N_A_299_392#_M1008_s VNB NSHORT L=0.15
+ W=0.74 AD=0.141175 AS=0.24175 PD=1.125 PS=2.14 NRD=6.48 NRS=6.48 M=1 R=4.93333
+ SA=75000.2 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1004 N_A_494_392#_M1004_d N_A_299_392#_M1004_g N_VGND_M1008_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.20255 AS=0.141175 PD=2.07 PS=1.125 NRD=1.62 NRS=9.72 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1037 N_A_699_463#_M1037_d N_A_299_392#_M1037_g N_A_37_78#_M1037_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1155 PD=0.77 PS=1.39 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.6 A=0.063 P=1.14 MULT=1
MM1034 A_812_138# N_A_494_392#_M1034_g N_A_699_463#_M1037_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1018 A_890_138# N_A_834_355#_M1018_g A_812_138# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75003.7 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_RESET_B_M1029_g A_890_138# VNB NSHORT L=0.15 W=0.42
+ AD=0.221767 AS=0.0504 PD=1.26 PS=0.66 NRD=135.144 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1009 N_A_834_355#_M1009_d N_A_699_463#_M1009_g N_VGND_M1029_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.47175 AS=0.390733 PD=2.015 PS=2.22 NRD=0 NRS=76.704 M=1
+ R=4.93333 SA=75001.6 SB=75002.9 A=0.111 P=1.78 MULT=1
MM1001 N_A_1350_392#_M1001_d N_A_494_392#_M1001_g N_A_834_355#_M1009_d VNB
+ NSHORT L=0.15 W=0.74 AD=0.292172 AS=0.47175 PD=2.09241 PS=2.015 NRD=0
+ NRS=11.34 M=1 R=4.93333 SA=75003.1 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1035 A_1647_81# N_A_299_392#_M1035_g N_A_1350_392#_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.165828 PD=0.66 PS=1.18759 NRD=18.564 NRS=49.992 M=1
+ R=2.8 SA=75003.7 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_1678_395#_M1020_g A_1647_81# VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=7.14 NRS=18.564 M=1 R=2.8 SA=75004.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1033 A_1827_81# N_RESET_B_M1033_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=15.708 M=1 R=2.8 SA=75004.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1027 N_A_1678_395#_M1027_d N_A_1350_392#_M1027_g A_1827_81# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75005
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_2010_409#_M1013_d N_A_1350_392#_M1013_g N_VGND_M1013_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 M=1
+ R=4.93333 SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_A_2010_409#_M1000_g N_Q_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.13875 PD=2.05 PS=1.115 NRD=0 NRS=7.296 M=1 R=4.93333 SA=75000.2
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_A_2010_409#_M1016_g N_Q_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.13875 PD=1.09 PS=1.115 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1028 N_VGND_M1016_d N_A_2010_409#_M1028_g N_Q_M1028_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1036 N_VGND_M1036_d N_A_2010_409#_M1036_g N_Q_M1028_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2035 AS=0.1036 PD=2.03 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1021 N_A_37_78#_M1021_d N_D_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.063 AS=0.1218 PD=0.72 PS=1.42 NRD=4.6886 NRS=4.6886 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1022 N_VPWR_M1022_d N_RESET_B_M1022_g N_A_37_78#_M1021_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1197 AS=0.063 PD=1.41 PS=0.72 NRD=0 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_CLK_M1010_g N_A_299_392#_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.3223 PD=1.3 PS=2.75 NRD=1.9503 NRS=17.73 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1017 N_A_494_392#_M1017_d N_A_299_392#_M1017_g N_VPWR_M1010_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.285 AS=0.15 PD=2.57 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1006 N_A_699_463#_M1006_d N_A_494_392#_M1006_g N_A_37_78#_M1006_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.063 AS=0.1218 PD=0.72 PS=1.42 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1011 A_789_463# N_A_299_392#_M1011_g N_A_699_463#_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.063 PD=0.66 PS=0.72 NRD=30.4759 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1026 N_VPWR_M1026_d N_A_834_355#_M1026_g A_789_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1295 AS=0.0504 PD=1.115 PS=0.66 NRD=118.811 NRS=30.4759 M=1 R=2.8
+ SA=75001.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1025 N_A_699_463#_M1025_d N_RESET_B_M1025_g N_VPWR_M1026_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1218 AS=0.1295 PD=1.42 PS=1.115 NRD=4.6886 NRS=118.811 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 N_A_834_355#_M1015_d N_A_699_463#_M1015_g N_VPWR_M1015_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.2845 PD=1.3 PS=2.68 NRD=1.9503 NRS=2.9353 M=1
+ R=6.66667 SA=75000.2 SB=75003.2 A=0.15 P=2.3 MULT=1
MM1024 N_A_1350_392#_M1024_d N_A_299_392#_M1024_g N_A_834_355#_M1015_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.473521 AS=0.15 PD=3.14789 PS=1.3 NRD=69.9153
+ NRS=1.9503 M=1 R=6.66667 SA=75000.7 SB=75002.8 A=0.15 P=2.3 MULT=1
MM1007 A_1627_493# N_A_494_392#_M1007_g N_A_1350_392#_M1024_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.198879 PD=0.69 PS=1.32211 NRD=37.5088 NRS=4.6886 M=1
+ R=2.8 SA=75002.1 SB=75005 A=0.063 P=1.14 MULT=1
MM1038 N_VPWR_M1038_d N_A_1678_395#_M1038_g A_1627_493# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.0567 PD=0.81 PS=0.69 NRD=23.443 NRS=37.5088 M=1 R=2.8
+ SA=75002.5 SB=75004.6 A=0.063 P=1.14 MULT=1
MM1014 N_A_1678_395#_M1014_d N_RESET_B_M1014_g N_VPWR_M1038_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.063 AS=0.0819 PD=0.72 PS=0.81 NRD=4.6886 NRS=28.1316 M=1 R=2.8
+ SA=75003 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1023 N_VPWR_M1023_d N_A_1350_392#_M1023_g N_A_1678_395#_M1014_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0868 AS=0.063 PD=0.796667 PS=0.72 NRD=23.443 NRS=4.6886 M=1
+ R=2.8 SA=75003.5 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_2010_409#_M1003_d N_A_1350_392#_M1003_g N_VPWR_M1023_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.126 AS=0.1736 PD=1.14 PS=1.59333 NRD=2.3443 NRS=5.8509 M=1
+ R=5.6 SA=75002.1 SB=75003.1 A=0.126 P=1.98 MULT=1
MM1030 N_A_2010_409#_M1003_d N_A_1350_392#_M1030_g N_VPWR_M1030_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.126 AS=0.1596 PD=1.14 PS=1.26429 NRD=2.3443 NRS=14.0658 M=1
+ R=5.6 SA=75002.5 SB=75002.6 A=0.126 P=1.98 MULT=1
MM1005 N_VPWR_M1030_s N_A_2010_409#_M1005_g N_Q_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.2128 AS=0.1932 PD=1.68571 PS=1.465 NRD=2.6201 NRS=9.6727 M=1
+ R=7.46667 SA=75002.3 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1019 N_VPWR_M1019_d N_A_2010_409#_M1019_g N_Q_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.434 AS=0.1932 PD=1.895 PS=1.465 NRD=2.6201 NRS=1.7533 M=1
+ R=7.46667 SA=75002.8 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1031 N_VPWR_M1019_d N_A_2010_409#_M1031_g N_Q_M1031_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.434 AS=0.168 PD=1.895 PS=1.42 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75003.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1032 N_VPWR_M1032_d N_A_2010_409#_M1032_g N_Q_M1031_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75004.2 SB=75000.3 A=0.168 P=2.54 MULT=1
DX39_noxref VNB VPB NWDIODE A=25.4742 P=31.6
c_135 VNB 0 1.974e-19 $X=0 $Y=0
c_1947 A_1627_493# 0 1.00633e-19 $X=8.135 $Y=2.465
*
.include "sky130_fd_sc_ls__dfrtp_4.pxi.spice"
*
.ends
*
*
