* File: sky130_fd_sc_ls__nand2b_1.pex.spice
* Created: Wed Sep  2 11:11:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NAND2B_1%A_N 3 5 7 8 9 13
c32 5 0 3.22862e-20 $X=0.505 $Y=1.765
r33 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.465 $X2=0.61 $Y2=1.465
r34 13 15 13.8279 $w=3.66e-07 $l=1.05e-07 $layer=POLY_cond $X=0.505 $Y=1.532
+ $X2=0.61 $Y2=1.532
r35 12 13 1.31694 $w=3.66e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.532
+ $X2=0.505 $Y2=1.532
r36 9 16 2.74101 $w=4.78e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.54 $X2=0.61
+ $Y2=1.54
r37 8 16 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.54 $X2=0.61
+ $Y2=1.54
r38 5 13 23.7042 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.532
r39 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.26
r40 1 12 23.7042 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.532
r41 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__NAND2B_1%B 1 3 6 8 12
c35 12 0 3.22862e-20 $X=1.18 $Y=1.515
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.18
+ $Y=1.515 $X2=1.18 $Y2=1.515
r37 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.18 $Y=1.665
+ $X2=1.18 $Y2=1.515
r38 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.27 $Y=1.35
+ $X2=1.18 $Y2=1.515
r39 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.27 $Y=1.35 $X2=1.27
+ $Y2=0.74
r40 1 11 52.2586 $w=2.99e-07 $l=2.52488e-07 $layer=POLY_cond $X=1.175 $Y=1.765
+ $X2=1.18 $Y2=1.515
r41 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.175 $Y=1.765
+ $X2=1.175 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NAND2B_1%A_27_112# 1 2 9 11 13 16 20 21 22 27 29 31
+ 33
c69 27 0 1.74227e-19 $X=1.6 $Y=1.95
r70 31 34 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=1.465
+ $X2=1.715 $Y2=1.63
r71 31 33 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=1.465
+ $X2=1.715 $Y2=1.3
r72 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.75
+ $Y=1.465 $X2=1.75 $Y2=1.465
r73 27 34 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.6 $Y=1.95 $X2=1.6
+ $Y2=1.63
r74 24 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.6 $Y=1.13 $X2=1.6
+ $Y2=1.3
r75 23 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r76 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.515 $Y=2.035
+ $X2=1.6 $Y2=1.95
r77 22 23 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=1.515 $Y=2.035
+ $X2=0.445 $Y2=2.035
r78 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.515 $Y=1.045
+ $X2=1.6 $Y2=1.13
r79 20 21 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=1.515 $Y=1.045
+ $X2=0.38 $Y2=1.045
r80 14 21 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.247 $Y=0.96
+ $X2=0.38 $Y2=1.045
r81 14 16 5.43605 $w=2.63e-07 $l=1.25e-07 $layer=LI1_cond $X=0.247 $Y=0.96
+ $X2=0.247 $Y2=0.835
r82 11 32 61.4066 $w=2.86e-07 $l=3.3541e-07 $layer=POLY_cond $X=1.675 $Y=1.765
+ $X2=1.75 $Y2=1.465
r83 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.675 $Y=1.765
+ $X2=1.675 $Y2=2.4
r84 7 32 38.6549 $w=2.86e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.66 $Y=1.3
+ $X2=1.75 $Y2=1.465
r85 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.66 $Y=1.3 $X2=1.66
+ $Y2=0.74
r86 2 29 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r87 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__NAND2B_1%VPWR 1 2 11 17 20 21 22 29 30 33
r29 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 27 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r33 24 33 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=0.915 $Y=3.33
+ $X2=0.782 $Y2=3.33
r34 24 26 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.915 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 20 26 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 20 21 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.902 $Y2=3.33
r39 19 29 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.07 $Y=3.33 $X2=2.16
+ $Y2=3.33
r40 19 21 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.07 $Y=3.33
+ $X2=1.902 $Y2=3.33
r41 15 21 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.902 $Y=3.245
+ $X2=1.902 $Y2=3.33
r42 15 17 14.7926 $w=3.33e-07 $l=4.3e-07 $layer=LI1_cond $X=1.902 $Y=3.245
+ $X2=1.902 $Y2=2.815
r43 11 14 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=0.782 $Y=2.455
+ $X2=0.782 $Y2=2.795
r44 9 33 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.782 $Y=3.245
+ $X2=0.782 $Y2=3.33
r45 9 14 19.5698 $w=2.63e-07 $l=4.5e-07 $layer=LI1_cond $X=0.782 $Y=3.245
+ $X2=0.782 $Y2=2.795
r46 2 17 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=1.84 $X2=1.9 $Y2=2.815
r47 1 14 600 $w=1.7e-07 $l=1.06828e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.82 $Y2=2.795
r48 1 11 600 $w=1.7e-07 $l=7.25138e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.82 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__NAND2B_1%Y 1 2 7 11 14 15 16 17 21
r34 16 21 2.36995 $w=4.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.325 $Y=2.375
+ $X2=1.325 $Y2=2.46
r35 16 17 7.47549 $w=4.78e-07 $l=3e-07 $layer=LI1_cond $X=1.325 $Y=2.475
+ $X2=1.325 $Y2=2.775
r36 16 21 0.373774 $w=4.78e-07 $l=1.5e-08 $layer=LI1_cond $X=1.325 $Y=2.475
+ $X2=1.325 $Y2=2.46
r37 14 15 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=2.17 $Y=2.29
+ $X2=2.17 $Y2=1.13
r38 9 15 9.656 $w=3.98e-07 $l=2e-07 $layer=LI1_cond $X=2.055 $Y=0.93 $X2=2.055
+ $Y2=1.13
r39 9 11 11.9566 $w=3.98e-07 $l=4.15e-07 $layer=LI1_cond $X=2.055 $Y=0.93
+ $X2=2.055 $Y2=0.515
r40 8 16 6.69163 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=1.565 $Y=2.375
+ $X2=1.325 $Y2=2.375
r41 7 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.085 $Y=2.375
+ $X2=2.17 $Y2=2.29
r42 7 8 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.085 $Y=2.375
+ $X2=1.565 $Y2=2.375
r43 2 16 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.25
+ $Y=1.84 $X2=1.4 $Y2=2.455
r44 1 11 91 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=2 $X=1.735
+ $Y=0.37 $X2=1.94 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NAND2B_1%VGND 1 6 8 10 17 18 21
r22 21 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r23 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r24 15 21 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=0.885
+ $Y2=0
r25 15 17 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=2.16
+ $Y2=0
r26 13 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r27 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r28 10 21 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.885
+ $Y2=0
r29 10 12 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.24
+ $Y2=0
r30 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r31 8 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r32 8 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r33 4 21 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.885 $Y=0.085
+ $X2=0.885 $Y2=0
r34 4 6 11.0682 $w=6.68e-07 $l=6.2e-07 $layer=LI1_cond $X=0.885 $Y=0.085
+ $X2=0.885 $Y2=0.705
r35 1 6 91 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.56 $X2=1.055 $Y2=0.705
.ends

