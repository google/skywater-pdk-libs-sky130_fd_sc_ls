* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
X0 VPWR a_1021_97# a_1243_48# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 VGND a_1711_48# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 a_1243_48# a_828_74# a_1511_74# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X3 Q a_1711_48# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 a_301_74# a_828_74# a_1021_97# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_1021_97# a_828_74# a_1173_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_301_74# a_36_74# a_423_453# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_301_74# SCE a_450_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 Q_N a_2322_368# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 a_1691_508# a_1711_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VPWR SCE a_238_453# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_423_453# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 VPWR a_2322_368# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X13 a_1511_74# a_828_74# a_1691_508# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_1243_48# a_630_74# a_1511_74# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X15 a_1663_74# a_1711_48# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_2322_368# a_1711_48# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 Q a_1711_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X18 a_450_74# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_630_74# a_828_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X20 a_2322_368# a_1711_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VPWR a_630_74# a_828_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X22 a_223_74# D a_301_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VPWR CLK a_630_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X24 a_1021_97# a_630_74# a_1217_499# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 Q_N a_2322_368# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X26 a_1511_74# a_630_74# a_1663_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_36_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X28 a_1217_499# a_1243_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 a_301_74# a_630_74# a_1021_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_1173_97# a_1243_48# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_238_453# D a_301_74# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X32 VGND CLK a_630_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X33 VGND a_36_74# a_223_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 VPWR a_1511_74# a_1711_48# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 a_36_74# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 VGND a_1511_74# a_1711_48# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X37 VPWR a_1711_48# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X38 VGND a_1021_97# a_1243_48# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X39 VGND a_2322_368# Q_N VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
