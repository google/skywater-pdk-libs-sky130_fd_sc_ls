* File: sky130_fd_sc_ls__mux4_4.pxi.spice
* Created: Fri Aug 28 13:31:21 2020
* 
x_PM_SKY130_FD_SC_LS__MUX4_4%A1 N_A1_M1025_g N_A1_c_318_n N_A1_M1039_g
+ N_A1_M1028_g N_A1_c_319_n N_A1_M1041_g A1 A1 N_A1_c_317_n
+ PM_SKY130_FD_SC_LS__MUX4_4%A1
x_PM_SKY130_FD_SC_LS__MUX4_4%A0 N_A0_c_362_n N_A0_M1000_g N_A0_M1021_g
+ N_A0_M1022_g N_A0_c_363_n N_A0_M1008_g A0 A0 A0 N_A0_c_360_n N_A0_c_361_n
+ PM_SKY130_FD_SC_LS__MUX4_4%A0
x_PM_SKY130_FD_SC_LS__MUX4_4%A_758_306# N_A_758_306#_M1012_s
+ N_A_758_306#_M1030_s N_A_758_306#_c_431_n N_A_758_306#_M1023_g
+ N_A_758_306#_M1036_g N_A_758_306#_c_432_n N_A_758_306#_M1035_g
+ N_A_758_306#_M1042_g N_A_758_306#_c_421_n N_A_758_306#_c_422_n
+ N_A_758_306#_M1002_g N_A_758_306#_c_434_n N_A_758_306#_M1019_g
+ N_A_758_306#_c_423_n N_A_758_306#_M1051_g N_A_758_306#_c_435_n
+ N_A_758_306#_M1031_g N_A_758_306#_c_424_n N_A_758_306#_c_436_n
+ N_A_758_306#_c_425_n N_A_758_306#_c_533_p N_A_758_306#_c_426_n
+ N_A_758_306#_c_427_n N_A_758_306#_c_428_n N_A_758_306#_c_429_n
+ N_A_758_306#_c_430_n PM_SKY130_FD_SC_LS__MUX4_4%A_758_306#
x_PM_SKY130_FD_SC_LS__MUX4_4%S0 N_S0_c_556_n N_S0_c_578_n N_S0_M1003_g
+ N_S0_M1004_g N_S0_c_558_n N_S0_c_559_n N_S0_c_560_n N_S0_c_580_n N_S0_M1043_g
+ N_S0_M1047_g N_S0_c_562_n N_S0_M1012_g N_S0_c_564_n N_S0_c_565_n N_S0_c_582_n
+ N_S0_M1030_g N_S0_c_566_n N_S0_M1006_g N_S0_c_583_n N_S0_M1005_g N_S0_M1040_g
+ N_S0_c_584_n N_S0_M1045_g N_S0_c_569_n N_S0_c_570_n N_S0_c_571_n N_S0_c_572_n
+ N_S0_c_573_n N_S0_c_574_n S0 S0 S0 N_S0_c_576_n PM_SKY130_FD_SC_LS__MUX4_4%S0
x_PM_SKY130_FD_SC_LS__MUX4_4%A2 N_A2_c_732_n N_A2_c_739_n N_A2_M1007_g
+ N_A2_M1018_g N_A2_c_734_n N_A2_c_741_n N_A2_M1017_g N_A2_M1038_g A2 A2
+ N_A2_c_737_n PM_SKY130_FD_SC_LS__MUX4_4%A2
x_PM_SKY130_FD_SC_LS__MUX4_4%A3 N_A3_M1014_g N_A3_c_799_n N_A3_M1033_g
+ N_A3_c_794_n N_A3_M1027_g N_A3_c_800_n N_A3_M1046_g N_A3_c_795_n N_A3_c_796_n
+ A3 A3 N_A3_c_798_n PM_SKY130_FD_SC_LS__MUX4_4%A3
x_PM_SKY130_FD_SC_LS__MUX4_4%S1 N_S1_M1013_g N_S1_c_850_n N_S1_c_864_n
+ N_S1_M1001_g N_S1_M1015_g N_S1_c_852_n N_S1_c_866_n N_S1_M1044_g N_S1_c_853_n
+ N_S1_c_854_n N_S1_M1010_g N_S1_c_855_n N_S1_c_868_n N_S1_M1037_g N_S1_c_856_n
+ N_S1_c_857_n N_S1_c_858_n S1 N_S1_c_859_n N_S1_c_860_n S1 N_S1_c_861_n
+ N_S1_c_862_n PM_SKY130_FD_SC_LS__MUX4_4%S1
x_PM_SKY130_FD_SC_LS__MUX4_4%A_2489_347# N_A_2489_347#_M1010_s
+ N_A_2489_347#_M1037_s N_A_2489_347#_c_980_n N_A_2489_347#_M1011_g
+ N_A_2489_347#_M1009_g N_A_2489_347#_c_981_n N_A_2489_347#_M1020_g
+ N_A_2489_347#_M1048_g N_A_2489_347#_c_982_n N_A_2489_347#_c_983_n
+ N_A_2489_347#_c_976_n N_A_2489_347#_c_977_n N_A_2489_347#_c_978_n
+ N_A_2489_347#_c_987_n N_A_2489_347#_c_979_n
+ PM_SKY130_FD_SC_LS__MUX4_4%A_2489_347#
x_PM_SKY130_FD_SC_LS__MUX4_4%A_2199_74# N_A_2199_74#_M1013_s
+ N_A_2199_74#_M1015_s N_A_2199_74#_M1048_d N_A_2199_74#_M1001_d
+ N_A_2199_74#_M1044_d N_A_2199_74#_M1020_s N_A_2199_74#_c_1079_n
+ N_A_2199_74#_M1024_g N_A_2199_74#_M1016_g N_A_2199_74#_c_1080_n
+ N_A_2199_74#_M1032_g N_A_2199_74#_M1026_g N_A_2199_74#_c_1081_n
+ N_A_2199_74#_M1034_g N_A_2199_74#_M1029_g N_A_2199_74#_c_1082_n
+ N_A_2199_74#_M1049_g N_A_2199_74#_M1050_g N_A_2199_74#_c_1066_n
+ N_A_2199_74#_c_1098_n N_A_2199_74#_c_1084_n N_A_2199_74#_c_1085_n
+ N_A_2199_74#_c_1125_n N_A_2199_74#_c_1067_n N_A_2199_74#_c_1105_n
+ N_A_2199_74#_c_1068_n N_A_2199_74#_c_1086_n N_A_2199_74#_c_1087_n
+ N_A_2199_74#_c_1069_n N_A_2199_74#_c_1070_n N_A_2199_74#_c_1071_n
+ N_A_2199_74#_c_1072_n N_A_2199_74#_c_1073_n N_A_2199_74#_c_1074_n
+ N_A_2199_74#_c_1116_n N_A_2199_74#_c_1075_n N_A_2199_74#_c_1076_n
+ N_A_2199_74#_c_1077_n N_A_2199_74#_c_1078_n
+ PM_SKY130_FD_SC_LS__MUX4_4%A_2199_74#
x_PM_SKY130_FD_SC_LS__MUX4_4%VPWR N_VPWR_M1039_d N_VPWR_M1041_d N_VPWR_M1008_s
+ N_VPWR_M1030_d N_VPWR_M1007_s N_VPWR_M1017_s N_VPWR_M1046_d N_VPWR_M1037_d
+ N_VPWR_M1032_d N_VPWR_M1049_d N_VPWR_c_1271_n N_VPWR_c_1272_n N_VPWR_c_1273_n
+ N_VPWR_c_1274_n N_VPWR_c_1275_n N_VPWR_c_1276_n N_VPWR_c_1277_n
+ N_VPWR_c_1278_n N_VPWR_c_1279_n N_VPWR_c_1280_n N_VPWR_c_1281_n
+ N_VPWR_c_1282_n N_VPWR_c_1283_n N_VPWR_c_1284_n N_VPWR_c_1285_n
+ N_VPWR_c_1286_n N_VPWR_c_1287_n N_VPWR_c_1288_n VPWR N_VPWR_c_1289_n
+ N_VPWR_c_1290_n N_VPWR_c_1291_n N_VPWR_c_1292_n N_VPWR_c_1293_n
+ N_VPWR_c_1294_n N_VPWR_c_1295_n N_VPWR_c_1296_n N_VPWR_c_1297_n
+ N_VPWR_c_1270_n PM_SKY130_FD_SC_LS__MUX4_4%VPWR
x_PM_SKY130_FD_SC_LS__MUX4_4%A_116_392# N_A_116_392#_M1039_s
+ N_A_116_392#_M1023_d N_A_116_392#_c_1453_n N_A_116_392#_c_1454_n
+ N_A_116_392#_c_1455_n N_A_116_392#_c_1456_n N_A_116_392#_c_1451_n
+ N_A_116_392#_c_1452_n N_A_116_392#_c_1459_n
+ PM_SKY130_FD_SC_LS__MUX4_4%A_116_392#
x_PM_SKY130_FD_SC_LS__MUX4_4%A_296_392# N_A_296_392#_M1000_d
+ N_A_296_392#_M1003_d N_A_296_392#_c_1515_n N_A_296_392#_c_1516_n
+ N_A_296_392#_c_1517_n N_A_296_392#_c_1524_n
+ PM_SKY130_FD_SC_LS__MUX4_4%A_296_392#
x_PM_SKY130_FD_SC_LS__MUX4_4%A_509_392# N_A_509_392#_M1004_d
+ N_A_509_392#_M1047_d N_A_509_392#_M1042_s N_A_509_392#_M1009_s
+ N_A_509_392#_M1003_s N_A_509_392#_M1043_s N_A_509_392#_M1035_s
+ N_A_509_392#_M1001_s N_A_509_392#_c_1557_n N_A_509_392#_c_1545_n
+ N_A_509_392#_c_1558_n N_A_509_392#_c_1546_n N_A_509_392#_c_1547_n
+ N_A_509_392#_c_1559_n N_A_509_392#_c_1548_n N_A_509_392#_c_1560_n
+ N_A_509_392#_c_1549_n N_A_509_392#_c_1550_n N_A_509_392#_c_1630_n
+ N_A_509_392#_c_1561_n N_A_509_392#_c_1551_n N_A_509_392#_c_1562_n
+ N_A_509_392#_c_1552_n N_A_509_392#_c_1553_n N_A_509_392#_c_1554_n
+ N_A_509_392#_c_1635_n N_A_509_392#_c_1563_n N_A_509_392#_c_1564_n
+ N_A_509_392#_c_1565_n N_A_509_392#_c_1566_n N_A_509_392#_c_1555_n
+ N_A_509_392#_c_1556_n PM_SKY130_FD_SC_LS__MUX4_4%A_509_392#
x_PM_SKY130_FD_SC_LS__MUX4_4%A_1191_121# N_A_1191_121#_M1002_d
+ N_A_1191_121#_M1051_d N_A_1191_121#_M1040_s N_A_1191_121#_M1013_d
+ N_A_1191_121#_M1019_s N_A_1191_121#_M1031_s N_A_1191_121#_M1045_d
+ N_A_1191_121#_M1011_d N_A_1191_121#_c_1733_n N_A_1191_121#_c_1734_n
+ N_A_1191_121#_c_1743_n N_A_1191_121#_c_1744_n N_A_1191_121#_c_1761_n
+ N_A_1191_121#_c_1745_n N_A_1191_121#_c_1735_n N_A_1191_121#_c_1782_n
+ N_A_1191_121#_c_1736_n N_A_1191_121#_c_1773_n N_A_1191_121#_c_1737_n
+ N_A_1191_121#_c_1747_n N_A_1191_121#_c_1738_n N_A_1191_121#_c_1749_n
+ N_A_1191_121#_c_1739_n N_A_1191_121#_c_1740_n N_A_1191_121#_c_1750_n
+ N_A_1191_121#_c_1751_n N_A_1191_121#_c_1826_n N_A_1191_121#_c_1741_n
+ N_A_1191_121#_c_1752_n N_A_1191_121#_c_1742_n N_A_1191_121#_c_1753_n
+ PM_SKY130_FD_SC_LS__MUX4_4%A_1191_121#
x_PM_SKY130_FD_SC_LS__MUX4_4%A_1285_377# N_A_1285_377#_M1019_d
+ N_A_1285_377#_M1033_s N_A_1285_377#_c_1915_n N_A_1285_377#_c_1911_n
+ N_A_1285_377#_c_1912_n N_A_1285_377#_c_1913_n N_A_1285_377#_c_1926_n
+ N_A_1285_377#_c_1914_n PM_SKY130_FD_SC_LS__MUX4_4%A_1285_377#
x_PM_SKY130_FD_SC_LS__MUX4_4%A_1465_377# N_A_1465_377#_M1005_s
+ N_A_1465_377#_M1007_d N_A_1465_377#_c_1968_n N_A_1465_377#_c_1970_n
+ PM_SKY130_FD_SC_LS__MUX4_4%A_1465_377#
x_PM_SKY130_FD_SC_LS__MUX4_4%X N_X_M1016_d N_X_M1029_d N_X_M1024_s N_X_M1034_s
+ N_X_c_1996_n N_X_c_1989_n N_X_c_1997_n N_X_c_1998_n N_X_c_1990_n N_X_c_1991_n
+ N_X_c_1999_n N_X_c_1992_n N_X_c_2000_n N_X_c_1993_n N_X_c_2001_n N_X_c_1994_n
+ X X PM_SKY130_FD_SC_LS__MUX4_4%X
x_PM_SKY130_FD_SC_LS__MUX4_4%VGND N_VGND_M1025_d N_VGND_M1028_d N_VGND_M1022_s
+ N_VGND_M1012_d N_VGND_M1018_s N_VGND_M1038_s N_VGND_M1027_s N_VGND_M1010_d
+ N_VGND_M1026_s N_VGND_M1050_s N_VGND_c_2072_n N_VGND_c_2073_n N_VGND_c_2074_n
+ N_VGND_c_2075_n N_VGND_c_2076_n N_VGND_c_2114_n N_VGND_c_2077_n
+ N_VGND_c_2078_n N_VGND_c_2079_n N_VGND_c_2080_n N_VGND_c_2081_n
+ N_VGND_c_2082_n N_VGND_c_2083_n N_VGND_c_2084_n N_VGND_c_2085_n
+ N_VGND_c_2086_n N_VGND_c_2087_n N_VGND_c_2088_n N_VGND_c_2089_n
+ N_VGND_c_2090_n N_VGND_c_2091_n VGND N_VGND_c_2092_n N_VGND_c_2093_n
+ N_VGND_c_2094_n N_VGND_c_2095_n N_VGND_c_2096_n N_VGND_c_2097_n
+ N_VGND_c_2098_n N_VGND_c_2099_n N_VGND_c_2100_n
+ PM_SKY130_FD_SC_LS__MUX4_4%VGND
x_PM_SKY130_FD_SC_LS__MUX4_4%A_114_126# N_A_114_126#_M1025_s
+ N_A_114_126#_M1004_s N_A_114_126#_c_2274_n N_A_114_126#_c_2275_n
+ N_A_114_126#_c_2276_n N_A_114_126#_c_2277_n N_A_114_126#_c_2278_n
+ N_A_114_126#_c_2289_n N_A_114_126#_c_2279_n
+ PM_SKY130_FD_SC_LS__MUX4_4%A_114_126#
x_PM_SKY130_FD_SC_LS__MUX4_4%A_299_126# N_A_299_126#_M1021_d
+ N_A_299_126#_M1036_d N_A_299_126#_c_2324_n N_A_299_126#_c_2325_n
+ N_A_299_126#_c_2326_n N_A_299_126#_c_2327_n N_A_299_126#_c_2328_n
+ PM_SKY130_FD_SC_LS__MUX4_4%A_299_126#
x_PM_SKY130_FD_SC_LS__MUX4_4%A_1278_121# N_A_1278_121#_M1002_s
+ N_A_1278_121#_M1018_d N_A_1278_121#_c_2366_n N_A_1278_121#_c_2367_n
+ N_A_1278_121#_c_2368_n N_A_1278_121#_c_2369_n N_A_1278_121#_c_2370_n
+ N_A_1278_121#_c_2371_n N_A_1278_121#_c_2372_n
+ PM_SKY130_FD_SC_LS__MUX4_4%A_1278_121#
x_PM_SKY130_FD_SC_LS__MUX4_4%A_1450_121# N_A_1450_121#_M1006_d
+ N_A_1450_121#_M1014_d N_A_1450_121#_c_2419_n N_A_1450_121#_c_2420_n
+ N_A_1450_121#_c_2421_n N_A_1450_121#_c_2422_n N_A_1450_121#_c_2423_n
+ PM_SKY130_FD_SC_LS__MUX4_4%A_1450_121#
cc_1 VNB N_A1_M1025_g 0.0253008f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.95
cc_2 VNB N_A1_M1028_g 0.0200691f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.95
cc_3 VNB A1 0.00939308f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_A1_c_317_n 0.0368261f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.667
cc_5 VNB N_A0_M1021_g 0.0215995f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_6 VNB N_A0_M1022_g 0.0253354f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.95
cc_7 VNB A0 0.00608988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A0_c_360_n 0.0211455f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.667
cc_9 VNB N_A0_c_361_n 0.0196575f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.615
cc_10 VNB N_A_758_306#_M1036_g 0.0170312f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.885
cc_11 VNB N_A_758_306#_M1042_g 0.020382f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.667
cc_12 VNB N_A_758_306#_c_421_n 0.0246711f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.615
cc_13 VNB N_A_758_306#_c_422_n 0.0194199f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.615
cc_14 VNB N_A_758_306#_c_423_n 0.014905f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_15 VNB N_A_758_306#_c_424_n 0.0143874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_758_306#_c_425_n 0.00207742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_758_306#_c_426_n 0.0298973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_758_306#_c_427_n 0.00188816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_758_306#_c_428_n 0.0218401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_758_306#_c_429_n 0.0150421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_758_306#_c_430_n 0.0477444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_S0_c_556_n 0.0121349f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.95
cc_23 VNB N_S0_M1004_g 0.0240024f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.95
cc_24 VNB N_S0_c_558_n 0.0191625f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.95
cc_25 VNB N_S0_c_559_n 0.012611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_S0_c_560_n 0.0108562f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.46
cc_27 VNB N_S0_M1047_g 0.0228453f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.667
cc_28 VNB N_S0_c_562_n 0.124248f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.667
cc_29 VNB N_S0_M1012_g 0.0129586f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_30 VNB N_S0_c_564_n 0.00853501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_S0_c_565_n 0.0245856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_S0_c_566_n 0.210692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_S0_M1006_g 0.015698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_S0_M1040_g 0.0199871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_S0_c_569_n 0.0674609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_S0_c_570_n 0.0143757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_S0_c_571_n 0.0116326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_S0_c_572_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_S0_c_573_n 0.00732516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_S0_c_574_n 0.0258376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB S0 0.00433756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_S0_c_576_n 0.0270364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A2_c_732_n 0.00379398f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.95
cc_44 VNB N_A2_M1018_g 0.0272771f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.45
cc_45 VNB N_A2_c_734_n 0.00342908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A2_M1038_g 0.0232221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB A2 0.00398279f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.667
cc_48 VNB N_A2_c_737_n 0.0521472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A3_M1014_g 0.0343392f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.95
cc_50 VNB N_A3_c_794_n 0.0173391f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.45
cc_51 VNB N_A3_c_795_n 0.0127568f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_52 VNB N_A3_c_796_n 0.0149455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB A3 0.00455884f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.667
cc_54 VNB N_A3_c_798_n 0.0312433f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_55 VNB N_S1_M1013_g 0.0250832f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.95
cc_56 VNB N_S1_c_850_n 0.00889551f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_57 VNB N_S1_M1015_g 0.0246191f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.885
cc_58 VNB N_S1_c_852_n 0.00825093f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_59 VNB N_S1_c_853_n 0.0298116f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.667
cc_60 VNB N_S1_c_854_n 0.0209511f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.667
cc_61 VNB N_S1_c_855_n 0.0079111f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.667
cc_62 VNB N_S1_c_856_n 0.0550093f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_63 VNB N_S1_c_857_n 0.0130751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_S1_c_858_n 0.026117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_S1_c_859_n 0.0348594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_S1_c_860_n 0.0364686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_S1_c_861_n 0.00294663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_S1_c_862_n 0.00253735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_2489_347#_M1009_g 0.0350434f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=1.885
cc_70 VNB N_A_2489_347#_M1048_g 0.0395546f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.667
cc_71 VNB N_A_2489_347#_c_976_n 0.00698854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_2489_347#_c_977_n 7.73014e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_2489_347#_c_978_n 0.0268228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_2489_347#_c_979_n 0.00368999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_2199_74#_M1016_g 0.0242761f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.667
cc_76 VNB N_A_2199_74#_M1026_g 0.0203684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_2199_74#_M1029_g 0.0209263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_2199_74#_M1050_g 0.0232593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_2199_74#_c_1066_n 0.00856582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_2199_74#_c_1067_n 0.00365532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_2199_74#_c_1068_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_2199_74#_c_1069_n 0.00589658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2199_74#_c_1070_n 0.0160232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_2199_74#_c_1071_n 0.00273158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_2199_74#_c_1072_n 0.00150988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_2199_74#_c_1073_n 0.012286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2199_74#_c_1074_n 0.00378272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_2199_74#_c_1075_n 9.79592e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_2199_74#_c_1076_n 0.00151123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_2199_74#_c_1077_n 0.00325932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_2199_74#_c_1078_n 0.112672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VPWR_c_1270_n 0.701046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_116_392#_c_1451_n 0.00638497f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_94 VNB N_A_116_392#_c_1452_n 0.00221343f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_95 VNB N_A_509_392#_c_1545_n 0.00921432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_509_392#_c_1546_n 0.00340257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_509_392#_c_1547_n 0.016329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_509_392#_c_1548_n 0.00636936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_509_392#_c_1549_n 0.00281722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_509_392#_c_1550_n 5.89755e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_509_392#_c_1551_n 0.0108906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_509_392#_c_1552_n 2.82947e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_509_392#_c_1553_n 0.00167754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_509_392#_c_1554_n 0.00269263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_509_392#_c_1555_n 0.00133979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_509_392#_c_1556_n 0.00187902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1191_121#_c_1733_n 0.00217675f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=1.667
cc_108 VNB N_A_1191_121#_c_1734_n 0.00619748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1191_121#_c_1735_n 0.00140514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_1191_121#_c_1736_n 0.00347953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_1191_121#_c_1737_n 0.00196259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_1191_121#_c_1738_n 0.0279051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1191_121#_c_1739_n 0.0034847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1191_121#_c_1740_n 0.00905591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_1191_121#_c_1741_n 0.00101203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_1191_121#_c_1742_n 0.00157069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_X_c_1989_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.667
cc_118 VNB N_X_c_1990_n 0.00275044f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.667
cc_119 VNB N_X_c_1991_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_120 VNB N_X_c_1992_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_X_c_1993_n 0.0087474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_X_c_1994_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB X 0.026544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2072_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2073_n 0.0122963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2074_n 0.0415587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2075_n 0.00303884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2076_n 0.00401119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2077_n 0.0109437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2078_n 0.0136696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2079_n 0.00420208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2080_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2081_n 0.0109995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2082_n 0.00852643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2083_n 0.00420208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2084_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2085_n 0.0257769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2086_n 0.0134389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2087_n 0.0670697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2088_n 0.0163794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2089_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2090_n 0.0967389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2091_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2092_n 0.0391102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2093_n 0.0737216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2094_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2095_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2096_n 0.0063135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2097_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2098_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2099_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2100_n 0.831397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_A_114_126#_c_2274_n 0.00135554f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=0.95
cc_154 VNB N_A_114_126#_c_2275_n 0.0218796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_A_114_126#_c_2276_n 0.00488309f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=1.885
cc_156 VNB N_A_114_126#_c_2277_n 0.00331078f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.46
cc_157 VNB N_A_114_126#_c_2278_n 9.57738e-19 $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_158 VNB N_A_114_126#_c_2279_n 0.00821615f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=1.667
cc_159 VNB N_A_299_126#_c_2324_n 0.00949813f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.46
cc_160 VNB N_A_299_126#_c_2325_n 0.01887f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.95
cc_161 VNB N_A_299_126#_c_2326_n 0.00111857f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.46
cc_162 VNB N_A_299_126#_c_2327_n 0.00202937f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_163 VNB N_A_299_126#_c_2328_n 0.00574177f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=1.667
cc_164 VNB N_A_1278_121#_c_2366_n 0.00265586f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=0.95
cc_165 VNB N_A_1278_121#_c_2367_n 0.0291012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_A_1278_121#_c_2368_n 0.00341436f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=1.885
cc_167 VNB N_A_1278_121#_c_2369_n 0.00206083f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.46
cc_168 VNB N_A_1278_121#_c_2370_n 0.00409716f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_169 VNB N_A_1278_121#_c_2371_n 0.00151359f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_170 VNB N_A_1278_121#_c_2372_n 0.00204804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_A_1450_121#_c_2419_n 0.00529172f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.46
cc_172 VNB N_A_1450_121#_c_2420_n 0.027156f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=0.95
cc_173 VNB N_A_1450_121#_c_2421_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.46
cc_174 VNB N_A_1450_121#_c_2422_n 0.00187699f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_175 VNB N_A_1450_121#_c_2423_n 0.00310731f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=1.667
cc_176 VPB N_A1_c_318_n 0.0179601f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_177 VPB N_A1_c_319_n 0.0158878f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.885
cc_178 VPB A1 0.00572761f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_179 VPB N_A1_c_317_n 0.0456921f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.667
cc_180 VPB N_A0_c_362_n 0.0156304f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.45
cc_181 VPB N_A0_c_363_n 0.0173356f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.885
cc_182 VPB A0 0.00431663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A0_c_360_n 0.0321182f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.667
cc_184 VPB N_A0_c_361_n 0.0167624f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.615
cc_185 VPB N_A_758_306#_c_431_n 0.0149459f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_186 VPB N_A_758_306#_c_432_n 0.0174904f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_187 VPB N_A_758_306#_c_421_n 0.0303755f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.615
cc_188 VPB N_A_758_306#_c_434_n 0.0162802f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_189 VPB N_A_758_306#_c_435_n 0.0138187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_758_306#_c_436_n 0.0157165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_758_306#_c_425_n 5.65058e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_758_306#_c_426_n 0.012178f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_758_306#_c_427_n 5.97595e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_758_306#_c_429_n 0.00808002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_758_306#_c_430_n 0.0343925f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_S0_c_556_n 0.00729967f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.95
cc_197 VPB N_S0_c_578_n 0.0231052f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.95
cc_198 VPB N_S0_c_560_n 0.0065055f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_199 VPB N_S0_c_580_n 0.0220514f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_200 VPB N_S0_c_565_n 9.04465e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_S0_c_582_n 0.0288551f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_202 VPB N_S0_c_583_n 0.0141878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_S0_c_584_n 0.0178837f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_S0_c_574_n 0.019332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB S0 0.00850506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_S0_c_576_n 0.0252532f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A2_c_732_n 0.00794851f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.95
cc_208 VPB N_A2_c_739_n 0.0263561f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.95
cc_209 VPB N_A2_c_734_n 0.00686619f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A2_c_741_n 0.0232583f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.885
cc_211 VPB A2 0.00397864f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.667
cc_212 VPB N_A3_c_799_n 0.0168986f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_213 VPB N_A3_c_800_n 0.0164708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB A3 0.00245853f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.667
cc_215 VPB N_A3_c_798_n 0.0363067f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_216 VPB N_S1_c_850_n 0.00889551f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_217 VPB N_S1_c_864_n 0.0248709f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_218 VPB N_S1_c_852_n 0.0078279f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_219 VPB N_S1_c_866_n 0.0212458f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_220 VPB N_S1_c_855_n 8.6742e-19 $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.667
cc_221 VPB N_S1_c_868_n 0.026577f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_222 VPB N_S1_c_861_n 0.00376745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_2489_347#_c_980_n 0.0155129f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_224 VPB N_A_2489_347#_c_981_n 0.0207807f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_225 VPB N_A_2489_347#_c_982_n 0.0219737f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.667
cc_226 VPB N_A_2489_347#_c_983_n 0.0223434f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.667
cc_227 VPB N_A_2489_347#_c_976_n 0.00106366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_2489_347#_c_977_n 0.00203626f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_2489_347#_c_978_n 0.0496682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_2489_347#_c_987_n 0.00442592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_2199_74#_c_1079_n 0.0161953f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.667
cc_232 VPB N_A_2199_74#_c_1080_n 0.015621f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_233 VPB N_A_2199_74#_c_1081_n 0.0156183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_2199_74#_c_1082_n 0.0164169f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_2199_74#_c_1066_n 0.00977476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_2199_74#_c_1084_n 0.00187959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_2199_74#_c_1085_n 0.00232324f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_2199_74#_c_1086_n 0.00258185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_2199_74#_c_1087_n 0.0135482f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_2199_74#_c_1078_n 0.0270583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1271_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1272_n 0.0514046f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1273_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1274_n 0.0118293f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1275_n 0.022681f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1276_n 0.00831227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1277_n 0.0133578f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1278_n 0.0082016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1279_n 0.0131478f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1280_n 0.0438947f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1281_n 0.0141618f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1282_n 0.0195396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1283_n 0.0196689f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1284_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1285_n 0.09287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1286_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1287_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1288_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1289_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1290_n 0.0194914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1291_n 0.0753801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1292_n 0.0634408f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1293_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1294_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1295_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1296_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1297_n 0.0141964f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1270_n 0.187693f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_A_116_392#_c_1453_n 0.00183558f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_270 VPB N_A_116_392#_c_1454_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.95
cc_271 VPB N_A_116_392#_c_1455_n 0.00738029f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_A_116_392#_c_1456_n 0.00504555f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_273 VPB N_A_116_392#_c_1451_n 0.0102103f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_274 VPB N_A_116_392#_c_1452_n 0.00118275f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_275 VPB N_A_116_392#_c_1459_n 0.00293562f $X=-0.19 $Y=1.66 $X2=0.495
+ $Y2=1.667
cc_276 VPB N_A_296_392#_c_1515_n 0.00834688f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.95
cc_277 VPB N_A_296_392#_c_1516_n 0.00274988f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_278 VPB N_A_296_392#_c_1517_n 0.00289649f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_279 VPB N_A_509_392#_c_1557_n 0.00237811f $X=-0.19 $Y=1.66 $X2=0.955
+ $Y2=1.667
cc_280 VPB N_A_509_392#_c_1558_n 0.00290856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_509_392#_c_1559_n 0.0071671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_A_509_392#_c_1560_n 0.00716705f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_509_392#_c_1561_n 0.00688319f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_A_509_392#_c_1562_n 0.0022931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_509_392#_c_1563_n 0.0328248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_A_509_392#_c_1564_n 0.00237732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_A_509_392#_c_1565_n 0.00344421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_288 VPB N_A_509_392#_c_1566_n 0.00121179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_289 VPB N_A_509_392#_c_1555_n 0.0026961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_A_509_392#_c_1556_n 0.00248628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_291 VPB N_A_1191_121#_c_1743_n 0.00344446f $X=-0.19 $Y=1.66 $X2=0.72
+ $Y2=1.615
cc_292 VPB N_A_1191_121#_c_1744_n 0.0101364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_A_1191_121#_c_1745_n 0.00304938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_A_1191_121#_c_1736_n 0.00334157f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_A_1191_121#_c_1747_n 0.0393704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_A_1191_121#_c_1738_n 0.0068711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_A_1191_121#_c_1749_n 0.0176439f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_A_1191_121#_c_1750_n 0.0185971f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_299 VPB N_A_1191_121#_c_1751_n 0.00349119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_300 VPB N_A_1191_121#_c_1752_n 2.04274e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_301 VPB N_A_1191_121#_c_1753_n 0.0096214f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_302 VPB N_A_1285_377#_c_1911_n 0.0207262f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_303 VPB N_A_1285_377#_c_1912_n 0.00484594f $X=-0.19 $Y=1.66 $X2=0.955
+ $Y2=1.885
cc_304 VPB N_A_1285_377#_c_1913_n 0.00780705f $X=-0.19 $Y=1.66 $X2=0.955
+ $Y2=2.46
cc_305 VPB N_A_1285_377#_c_1914_n 0.00797734f $X=-0.19 $Y=1.66 $X2=0.495
+ $Y2=1.667
cc_306 VPB N_A_1465_377#_c_1968_n 0.00582192f $X=-0.19 $Y=1.66 $X2=0.925
+ $Y2=0.95
cc_307 VPB N_X_c_1996_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_308 VPB N_X_c_1997_n 0.00209566f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.615
cc_309 VPB N_X_c_1998_n 0.00183475f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.667
cc_310 VPB N_X_c_1999_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_311 VPB N_X_c_2000_n 0.0101857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_312 VPB N_X_c_2001_n 0.00183475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_313 VPB X 0.00736649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_314 N_A1_c_319_n N_A0_c_362_n 0.0216655f $X=0.955 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_315 N_A1_M1028_g N_A0_M1021_g 0.0115976f $X=0.925 $Y=0.95 $X2=0 $Y2=0
cc_316 N_A1_c_317_n N_A0_M1021_g 9.69146e-19 $X=0.925 $Y=1.667 $X2=0 $Y2=0
cc_317 A1 A0 0.0247408f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_318 N_A1_c_317_n A0 0.00388845f $X=0.925 $Y=1.667 $X2=0 $Y2=0
cc_319 A1 N_A0_c_360_n 2.15092e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_320 N_A1_c_317_n N_A0_c_360_n 0.0201224f $X=0.925 $Y=1.667 $X2=0 $Y2=0
cc_321 N_A1_c_318_n N_VPWR_c_1272_n 0.00850369f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_322 A1 N_VPWR_c_1272_n 0.0205478f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_323 N_A1_c_317_n N_VPWR_c_1272_n 0.00335457f $X=0.925 $Y=1.667 $X2=0 $Y2=0
cc_324 N_A1_c_319_n N_VPWR_c_1273_n 0.0051932f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_325 N_A1_c_318_n N_VPWR_c_1289_n 0.00445602f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_326 N_A1_c_319_n N_VPWR_c_1289_n 0.00445602f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_327 N_A1_c_318_n N_VPWR_c_1270_n 0.00861084f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_328 N_A1_c_319_n N_VPWR_c_1270_n 0.00857673f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_329 N_A1_c_318_n N_A_116_392#_c_1453_n 0.00238159f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_330 N_A1_c_319_n N_A_116_392#_c_1453_n 9.95967e-19 $X=0.955 $Y=1.885 $X2=0
+ $Y2=0
cc_331 A1 N_A_116_392#_c_1453_n 0.0272953f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_332 N_A1_c_317_n N_A_116_392#_c_1453_n 0.0078875f $X=0.925 $Y=1.667 $X2=0
+ $Y2=0
cc_333 N_A1_c_318_n N_A_116_392#_c_1454_n 0.00939341f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_334 N_A1_c_319_n N_A_116_392#_c_1454_n 0.0101905f $X=0.955 $Y=1.885 $X2=0
+ $Y2=0
cc_335 N_A1_c_319_n N_A_116_392#_c_1455_n 0.0159795f $X=0.955 $Y=1.885 $X2=0
+ $Y2=0
cc_336 A1 N_VGND_c_2073_n 0.0206322f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_337 N_A1_c_317_n N_VGND_c_2073_n 0.00337787f $X=0.925 $Y=1.667 $X2=0 $Y2=0
cc_338 N_A1_M1025_g N_VGND_c_2074_n 0.00290289f $X=0.495 $Y=0.95 $X2=0 $Y2=0
cc_339 N_A1_M1025_g N_VGND_c_2075_n 0.0145041f $X=0.495 $Y=0.95 $X2=0 $Y2=0
cc_340 N_A1_M1028_g N_VGND_c_2075_n 0.0154359f $X=0.925 $Y=0.95 $X2=0 $Y2=0
cc_341 A1 N_VGND_c_2075_n 0.0398625f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_342 N_A1_c_317_n N_VGND_c_2075_n 0.00539292f $X=0.925 $Y=1.667 $X2=0 $Y2=0
cc_343 N_A1_M1025_g N_VGND_c_2092_n 0.00354577f $X=0.495 $Y=0.95 $X2=0 $Y2=0
cc_344 N_A1_M1028_g N_VGND_c_2092_n 2.33667e-19 $X=0.925 $Y=0.95 $X2=0 $Y2=0
cc_345 N_A1_M1025_g N_VGND_c_2100_n 0.00391696f $X=0.495 $Y=0.95 $X2=0 $Y2=0
cc_346 N_A1_M1025_g N_A_114_126#_c_2274_n 0.00626483f $X=0.495 $Y=0.95 $X2=0
+ $Y2=0
cc_347 N_A1_M1028_g N_A_114_126#_c_2274_n 0.00727484f $X=0.925 $Y=0.95 $X2=0
+ $Y2=0
cc_348 N_A1_M1028_g N_A_114_126#_c_2275_n 0.00455657f $X=0.925 $Y=0.95 $X2=0
+ $Y2=0
cc_349 A0 N_S0_c_556_n 8.62325e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_350 N_A0_c_361_n N_S0_c_556_n 0.006687f $X=2.19 $Y=1.635 $X2=0 $Y2=0
cc_351 N_A0_c_362_n N_VPWR_c_1273_n 0.0101085f $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_352 N_A0_c_363_n N_VPWR_c_1273_n 6.87135e-19 $X=1.905 $Y=1.885 $X2=0 $Y2=0
cc_353 N_A0_c_363_n N_VPWR_c_1274_n 0.00590397f $X=1.905 $Y=1.885 $X2=0 $Y2=0
cc_354 N_A0_c_362_n N_VPWR_c_1290_n 0.00413917f $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_355 N_A0_c_363_n N_VPWR_c_1290_n 0.00445602f $X=1.905 $Y=1.885 $X2=0 $Y2=0
cc_356 N_A0_c_362_n N_VPWR_c_1270_n 0.00818187f $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_357 N_A0_c_363_n N_VPWR_c_1270_n 0.00460221f $X=1.905 $Y=1.885 $X2=0 $Y2=0
cc_358 N_A0_c_362_n N_A_116_392#_c_1454_n 9.51579e-19 $X=1.405 $Y=1.885 $X2=0
+ $Y2=0
cc_359 N_A0_c_362_n N_A_116_392#_c_1455_n 0.0151078f $X=1.405 $Y=1.885 $X2=0
+ $Y2=0
cc_360 N_A0_c_363_n N_A_116_392#_c_1455_n 0.0128867f $X=1.905 $Y=1.885 $X2=0
+ $Y2=0
cc_361 A0 N_A_116_392#_c_1455_n 0.0857078f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_362 N_A0_c_360_n N_A_116_392#_c_1455_n 0.00785707f $X=1.995 $Y=1.635 $X2=0
+ $Y2=0
cc_363 N_A0_c_361_n N_A_116_392#_c_1455_n 0.00795903f $X=2.19 $Y=1.635 $X2=0
+ $Y2=0
cc_364 N_A0_c_363_n N_A_116_392#_c_1456_n 0.00194432f $X=1.905 $Y=1.885 $X2=0
+ $Y2=0
cc_365 A0 N_A_116_392#_c_1456_n 0.00227977f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_366 N_A0_c_360_n N_A_116_392#_c_1456_n 0.00203925f $X=1.995 $Y=1.635 $X2=0
+ $Y2=0
cc_367 A0 N_A_116_392#_c_1452_n 0.0151563f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_368 N_A0_c_361_n N_A_116_392#_c_1452_n 7.73608e-19 $X=2.19 $Y=1.635 $X2=0
+ $Y2=0
cc_369 N_A0_c_363_n N_A_296_392#_c_1515_n 0.0111269f $X=1.905 $Y=1.885 $X2=0
+ $Y2=0
cc_370 N_A0_c_362_n N_A_296_392#_c_1517_n 0.00272481f $X=1.405 $Y=1.885 $X2=0
+ $Y2=0
cc_371 N_A0_c_363_n N_A_296_392#_c_1517_n 0.0115156f $X=1.905 $Y=1.885 $X2=0
+ $Y2=0
cc_372 N_A0_M1022_g N_A_509_392#_c_1551_n 0.00280676f $X=1.85 $Y=0.95 $X2=0
+ $Y2=0
cc_373 N_A0_M1021_g N_VGND_c_2076_n 0.00308767f $X=1.42 $Y=0.95 $X2=0 $Y2=0
cc_374 A0 N_VGND_c_2076_n 0.0228477f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_375 N_A0_c_360_n N_VGND_c_2076_n 7.63156e-19 $X=1.995 $Y=1.635 $X2=0 $Y2=0
cc_376 N_A0_M1021_g N_VGND_c_2114_n 0.00569723f $X=1.42 $Y=0.95 $X2=0 $Y2=0
cc_377 N_A0_M1022_g N_VGND_c_2114_n 5.68292e-19 $X=1.85 $Y=0.95 $X2=0 $Y2=0
cc_378 N_A0_M1022_g N_VGND_c_2092_n 0.00258164f $X=1.85 $Y=0.95 $X2=0 $Y2=0
cc_379 N_A0_M1022_g N_VGND_c_2100_n 0.00360493f $X=1.85 $Y=0.95 $X2=0 $Y2=0
cc_380 N_A0_M1021_g N_A_114_126#_c_2274_n 6.3983e-19 $X=1.42 $Y=0.95 $X2=0 $Y2=0
cc_381 N_A0_M1021_g N_A_114_126#_c_2275_n 0.00692429f $X=1.42 $Y=0.95 $X2=0
+ $Y2=0
cc_382 N_A0_M1021_g N_A_114_126#_c_2277_n 0.0029318f $X=1.42 $Y=0.95 $X2=0 $Y2=0
cc_383 N_A0_M1022_g N_A_114_126#_c_2277_n 0.0067325f $X=1.85 $Y=0.95 $X2=0 $Y2=0
cc_384 N_A0_M1021_g N_A_114_126#_c_2278_n 0.00180292f $X=1.42 $Y=0.95 $X2=0
+ $Y2=0
cc_385 N_A0_M1022_g N_A_114_126#_c_2278_n 0.0117504f $X=1.85 $Y=0.95 $X2=0 $Y2=0
cc_386 N_A0_M1022_g N_A_299_126#_c_2324_n 0.0106426f $X=1.85 $Y=0.95 $X2=0 $Y2=0
cc_387 A0 N_A_299_126#_c_2324_n 0.0412064f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_388 N_A0_c_360_n N_A_299_126#_c_2324_n 0.00985359f $X=1.995 $Y=1.635 $X2=0
+ $Y2=0
cc_389 N_A0_M1021_g N_A_299_126#_c_2327_n 5.84569e-19 $X=1.42 $Y=0.95 $X2=0
+ $Y2=0
cc_390 N_A0_M1022_g N_A_299_126#_c_2327_n 0.00900763f $X=1.85 $Y=0.95 $X2=0
+ $Y2=0
cc_391 A0 N_A_299_126#_c_2327_n 0.0196736f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_392 N_A0_c_360_n N_A_299_126#_c_2327_n 0.00228163f $X=1.995 $Y=1.635 $X2=0
+ $Y2=0
cc_393 N_A0_M1022_g N_A_299_126#_c_2328_n 0.00320159f $X=1.85 $Y=0.95 $X2=0
+ $Y2=0
cc_394 N_A_758_306#_c_421_n N_S0_c_560_n 0.0197631f $X=4.42 $Y=1.547 $X2=0 $Y2=0
cc_395 N_A_758_306#_c_431_n N_S0_c_580_n 0.00773369f $X=3.88 $Y=1.885 $X2=0
+ $Y2=0
cc_396 N_A_758_306#_M1036_g N_S0_M1047_g 0.0126979f $X=3.905 $Y=0.915 $X2=0
+ $Y2=0
cc_397 N_A_758_306#_M1036_g N_S0_c_562_n 0.00882199f $X=3.905 $Y=0.915 $X2=0
+ $Y2=0
cc_398 N_A_758_306#_M1042_g N_S0_c_562_n 0.00903828f $X=4.335 $Y=0.915 $X2=0
+ $Y2=0
cc_399 N_A_758_306#_c_424_n N_S0_c_562_n 0.00506365f $X=5.11 $Y=0.515 $X2=0
+ $Y2=0
cc_400 N_A_758_306#_c_424_n N_S0_M1012_g 0.0111534f $X=5.11 $Y=0.515 $X2=0 $Y2=0
cc_401 N_A_758_306#_c_425_n N_S0_c_565_n 8.03098e-19 $X=6.365 $Y=1.53 $X2=0
+ $Y2=0
cc_402 N_A_758_306#_c_426_n N_S0_c_565_n 0.0205345f $X=4.875 $Y=1.515 $X2=0
+ $Y2=0
cc_403 N_A_758_306#_c_427_n N_S0_c_565_n 0.00452077f $X=5.2 $Y=1.515 $X2=0 $Y2=0
cc_404 N_A_758_306#_c_428_n N_S0_c_565_n 0.0174642f $X=6.035 $Y=1.53 $X2=0 $Y2=0
cc_405 N_A_758_306#_c_430_n N_S0_c_565_n 0.00463574f $X=6.745 $Y=1.587 $X2=0
+ $Y2=0
cc_406 N_A_758_306#_c_436_n N_S0_c_582_n 0.0113473f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_407 N_A_758_306#_c_422_n N_S0_c_566_n 0.00980793f $X=6.315 $Y=1.365 $X2=0
+ $Y2=0
cc_408 N_A_758_306#_c_423_n N_S0_c_566_n 0.00844637f $X=6.745 $Y=1.365 $X2=0
+ $Y2=0
cc_409 N_A_758_306#_c_423_n N_S0_M1006_g 0.0106844f $X=6.745 $Y=1.365 $X2=0
+ $Y2=0
cc_410 N_A_758_306#_c_430_n N_S0_M1006_g 0.011768f $X=6.745 $Y=1.587 $X2=0 $Y2=0
cc_411 N_A_758_306#_c_435_n N_S0_c_583_n 0.0176919f $X=6.8 $Y=1.81 $X2=0 $Y2=0
cc_412 N_A_758_306#_c_421_n N_S0_c_571_n 0.0126979f $X=4.42 $Y=1.547 $X2=0 $Y2=0
cc_413 N_A_758_306#_c_430_n N_S0_c_576_n 0.0114652f $X=6.745 $Y=1.587 $X2=0
+ $Y2=0
cc_414 N_A_758_306#_c_434_n N_VPWR_c_1275_n 0.00560884f $X=6.35 $Y=1.81 $X2=0
+ $Y2=0
cc_415 N_A_758_306#_c_436_n N_VPWR_c_1275_n 0.0763693f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_416 N_A_758_306#_c_428_n N_VPWR_c_1275_n 0.0171257f $X=6.035 $Y=1.53 $X2=0
+ $Y2=0
cc_417 N_A_758_306#_c_431_n N_VPWR_c_1291_n 0.00278257f $X=3.88 $Y=1.885 $X2=0
+ $Y2=0
cc_418 N_A_758_306#_c_432_n N_VPWR_c_1291_n 0.00278242f $X=4.33 $Y=1.885 $X2=0
+ $Y2=0
cc_419 N_A_758_306#_c_436_n N_VPWR_c_1291_n 0.011066f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_420 N_A_758_306#_c_434_n N_VPWR_c_1292_n 0.00479747f $X=6.35 $Y=1.81 $X2=0
+ $Y2=0
cc_421 N_A_758_306#_c_435_n N_VPWR_c_1292_n 8.35168e-19 $X=6.8 $Y=1.81 $X2=0
+ $Y2=0
cc_422 N_A_758_306#_c_431_n N_VPWR_c_1270_n 0.00354126f $X=3.88 $Y=1.885 $X2=0
+ $Y2=0
cc_423 N_A_758_306#_c_432_n N_VPWR_c_1270_n 0.00358622f $X=4.33 $Y=1.885 $X2=0
+ $Y2=0
cc_424 N_A_758_306#_c_434_n N_VPWR_c_1270_n 0.00469908f $X=6.35 $Y=1.81 $X2=0
+ $Y2=0
cc_425 N_A_758_306#_c_436_n N_VPWR_c_1270_n 0.00915947f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_426 N_A_758_306#_c_421_n N_A_116_392#_c_1451_n 0.0237362f $X=4.42 $Y=1.547
+ $X2=0 $Y2=0
cc_427 N_A_758_306#_c_431_n N_A_116_392#_c_1459_n 0.00422968f $X=3.88 $Y=1.885
+ $X2=0 $Y2=0
cc_428 N_A_758_306#_c_432_n N_A_116_392#_c_1459_n 0.00315068f $X=4.33 $Y=1.885
+ $X2=0 $Y2=0
cc_429 N_A_758_306#_c_421_n N_A_116_392#_c_1459_n 0.00358644f $X=4.42 $Y=1.547
+ $X2=0 $Y2=0
cc_430 N_A_758_306#_c_431_n N_A_509_392#_c_1558_n 0.0114074f $X=3.88 $Y=1.885
+ $X2=0 $Y2=0
cc_431 N_A_758_306#_c_432_n N_A_509_392#_c_1558_n 6.74657e-19 $X=4.33 $Y=1.885
+ $X2=0 $Y2=0
cc_432 N_A_758_306#_c_421_n N_A_509_392#_c_1558_n 4.08005e-19 $X=4.42 $Y=1.547
+ $X2=0 $Y2=0
cc_433 N_A_758_306#_M1036_g N_A_509_392#_c_1546_n 0.00203728f $X=3.905 $Y=0.915
+ $X2=0 $Y2=0
cc_434 N_A_758_306#_M1036_g N_A_509_392#_c_1547_n 0.00330666f $X=3.905 $Y=0.915
+ $X2=0 $Y2=0
cc_435 N_A_758_306#_M1042_g N_A_509_392#_c_1547_n 0.00283033f $X=4.335 $Y=0.915
+ $X2=0 $Y2=0
cc_436 N_A_758_306#_c_424_n N_A_509_392#_c_1547_n 0.00526842f $X=5.11 $Y=0.515
+ $X2=0 $Y2=0
cc_437 N_A_758_306#_c_431_n N_A_509_392#_c_1559_n 0.0108414f $X=3.88 $Y=1.885
+ $X2=0 $Y2=0
cc_438 N_A_758_306#_c_432_n N_A_509_392#_c_1559_n 0.0128044f $X=4.33 $Y=1.885
+ $X2=0 $Y2=0
cc_439 N_A_758_306#_c_436_n N_A_509_392#_c_1559_n 0.00526106f $X=5.115 $Y=1.985
+ $X2=0 $Y2=0
cc_440 N_A_758_306#_M1036_g N_A_509_392#_c_1548_n 7.22399e-19 $X=3.905 $Y=0.915
+ $X2=0 $Y2=0
cc_441 N_A_758_306#_M1042_g N_A_509_392#_c_1548_n 0.0098936f $X=4.335 $Y=0.915
+ $X2=0 $Y2=0
cc_442 N_A_758_306#_c_424_n N_A_509_392#_c_1548_n 0.0499741f $X=5.11 $Y=0.515
+ $X2=0 $Y2=0
cc_443 N_A_758_306#_c_432_n N_A_509_392#_c_1560_n 0.0100434f $X=4.33 $Y=1.885
+ $X2=0 $Y2=0
cc_444 N_A_758_306#_c_431_n N_A_509_392#_c_1562_n 0.00180969f $X=3.88 $Y=1.885
+ $X2=0 $Y2=0
cc_445 N_A_758_306#_M1042_g N_A_509_392#_c_1553_n 0.00183387f $X=4.335 $Y=0.915
+ $X2=0 $Y2=0
cc_446 N_A_758_306#_c_429_n N_A_509_392#_c_1553_n 0.00666801f $X=4.71 $Y=1.515
+ $X2=0 $Y2=0
cc_447 N_A_758_306#_M1030_s N_A_509_392#_c_1563_n 0.00456387f $X=4.97 $Y=1.84
+ $X2=0 $Y2=0
cc_448 N_A_758_306#_c_434_n N_A_509_392#_c_1563_n 0.00611384f $X=6.35 $Y=1.81
+ $X2=0 $Y2=0
cc_449 N_A_758_306#_c_435_n N_A_509_392#_c_1563_n 0.00611384f $X=6.8 $Y=1.81
+ $X2=0 $Y2=0
cc_450 N_A_758_306#_c_436_n N_A_509_392#_c_1563_n 0.023829f $X=5.115 $Y=1.985
+ $X2=0 $Y2=0
cc_451 N_A_758_306#_c_425_n N_A_509_392#_c_1563_n 0.00395434f $X=6.365 $Y=1.53
+ $X2=0 $Y2=0
cc_452 N_A_758_306#_c_426_n N_A_509_392#_c_1563_n 0.00523275f $X=4.875 $Y=1.515
+ $X2=0 $Y2=0
cc_453 N_A_758_306#_c_427_n N_A_509_392#_c_1563_n 0.0100335f $X=5.2 $Y=1.515
+ $X2=0 $Y2=0
cc_454 N_A_758_306#_c_428_n N_A_509_392#_c_1563_n 0.0143906f $X=6.035 $Y=1.53
+ $X2=0 $Y2=0
cc_455 N_A_758_306#_c_436_n N_A_509_392#_c_1564_n 6.54704e-19 $X=5.115 $Y=1.985
+ $X2=0 $Y2=0
cc_456 N_A_758_306#_c_432_n N_A_509_392#_c_1565_n 0.00265935f $X=4.33 $Y=1.885
+ $X2=0 $Y2=0
cc_457 N_A_758_306#_c_436_n N_A_509_392#_c_1565_n 0.062652f $X=5.115 $Y=1.985
+ $X2=0 $Y2=0
cc_458 N_A_758_306#_c_429_n N_A_509_392#_c_1565_n 0.00572494f $X=4.71 $Y=1.515
+ $X2=0 $Y2=0
cc_459 N_A_758_306#_c_431_n N_A_509_392#_c_1556_n 6.94525e-19 $X=3.88 $Y=1.885
+ $X2=0 $Y2=0
cc_460 N_A_758_306#_c_432_n N_A_509_392#_c_1556_n 0.00115539f $X=4.33 $Y=1.885
+ $X2=0 $Y2=0
cc_461 N_A_758_306#_M1042_g N_A_509_392#_c_1556_n 0.00492997f $X=4.335 $Y=0.915
+ $X2=0 $Y2=0
cc_462 N_A_758_306#_c_421_n N_A_509_392#_c_1556_n 0.0164572f $X=4.42 $Y=1.547
+ $X2=0 $Y2=0
cc_463 N_A_758_306#_c_424_n N_A_509_392#_c_1556_n 0.00515416f $X=5.11 $Y=0.515
+ $X2=0 $Y2=0
cc_464 N_A_758_306#_c_436_n N_A_509_392#_c_1556_n 0.00809031f $X=5.115 $Y=1.985
+ $X2=0 $Y2=0
cc_465 N_A_758_306#_c_426_n N_A_509_392#_c_1556_n 4.37509e-19 $X=4.875 $Y=1.515
+ $X2=0 $Y2=0
cc_466 N_A_758_306#_c_427_n N_A_509_392#_c_1556_n 0.0248912f $X=5.2 $Y=1.515
+ $X2=0 $Y2=0
cc_467 N_A_758_306#_c_429_n N_A_509_392#_c_1556_n 0.0126905f $X=4.71 $Y=1.515
+ $X2=0 $Y2=0
cc_468 N_A_758_306#_c_428_n N_A_1191_121#_c_1733_n 0.0208194f $X=6.035 $Y=1.53
+ $X2=0 $Y2=0
cc_469 N_A_758_306#_c_430_n N_A_1191_121#_c_1733_n 0.00347152f $X=6.745 $Y=1.587
+ $X2=0 $Y2=0
cc_470 N_A_758_306#_c_422_n N_A_1191_121#_c_1734_n 4.43891e-19 $X=6.315 $Y=1.365
+ $X2=0 $Y2=0
cc_471 N_A_758_306#_c_425_n N_A_1191_121#_c_1743_n 0.013784f $X=6.365 $Y=1.53
+ $X2=0 $Y2=0
cc_472 N_A_758_306#_c_428_n N_A_1191_121#_c_1743_n 0.00116029f $X=6.035 $Y=1.53
+ $X2=0 $Y2=0
cc_473 N_A_758_306#_c_430_n N_A_1191_121#_c_1743_n 0.00407674f $X=6.745 $Y=1.587
+ $X2=0 $Y2=0
cc_474 N_A_758_306#_c_434_n N_A_1191_121#_c_1744_n 0.0061053f $X=6.35 $Y=1.81
+ $X2=0 $Y2=0
cc_475 N_A_758_306#_c_422_n N_A_1191_121#_c_1761_n 0.0119972f $X=6.315 $Y=1.365
+ $X2=0 $Y2=0
cc_476 N_A_758_306#_c_423_n N_A_1191_121#_c_1761_n 0.0114803f $X=6.745 $Y=1.365
+ $X2=0 $Y2=0
cc_477 N_A_758_306#_c_425_n N_A_1191_121#_c_1761_n 0.0317383f $X=6.365 $Y=1.53
+ $X2=0 $Y2=0
cc_478 N_A_758_306#_c_430_n N_A_1191_121#_c_1761_n 0.00224206f $X=6.745 $Y=1.587
+ $X2=0 $Y2=0
cc_479 N_A_758_306#_c_434_n N_A_1191_121#_c_1745_n 0.0102328f $X=6.35 $Y=1.81
+ $X2=0 $Y2=0
cc_480 N_A_758_306#_c_435_n N_A_1191_121#_c_1745_n 0.0121432f $X=6.8 $Y=1.81
+ $X2=0 $Y2=0
cc_481 N_A_758_306#_c_425_n N_A_1191_121#_c_1745_n 0.0337976f $X=6.365 $Y=1.53
+ $X2=0 $Y2=0
cc_482 N_A_758_306#_c_430_n N_A_1191_121#_c_1745_n 0.00988402f $X=6.745 $Y=1.587
+ $X2=0 $Y2=0
cc_483 N_A_758_306#_c_423_n N_A_1191_121#_c_1736_n 0.00221303f $X=6.745 $Y=1.365
+ $X2=0 $Y2=0
cc_484 N_A_758_306#_c_435_n N_A_1191_121#_c_1736_n 0.00130706f $X=6.8 $Y=1.81
+ $X2=0 $Y2=0
cc_485 N_A_758_306#_c_533_p N_A_1191_121#_c_1736_n 0.0206343f $X=6.54 $Y=1.53
+ $X2=0 $Y2=0
cc_486 N_A_758_306#_c_430_n N_A_1191_121#_c_1736_n 0.005835f $X=6.745 $Y=1.587
+ $X2=0 $Y2=0
cc_487 N_A_758_306#_c_435_n N_A_1191_121#_c_1773_n 0.00412619f $X=6.8 $Y=1.81
+ $X2=0 $Y2=0
cc_488 N_A_758_306#_c_423_n N_A_1191_121#_c_1741_n 4.93723e-19 $X=6.745 $Y=1.365
+ $X2=0 $Y2=0
cc_489 N_A_758_306#_c_430_n N_A_1191_121#_c_1741_n 5.04279e-19 $X=6.745 $Y=1.587
+ $X2=0 $Y2=0
cc_490 N_A_758_306#_c_434_n N_A_1285_377#_c_1915_n 0.00836448f $X=6.35 $Y=1.81
+ $X2=0 $Y2=0
cc_491 N_A_758_306#_c_435_n N_A_1285_377#_c_1915_n 0.00924488f $X=6.8 $Y=1.81
+ $X2=0 $Y2=0
cc_492 N_A_758_306#_c_435_n N_A_1285_377#_c_1911_n 0.0106926f $X=6.8 $Y=1.81
+ $X2=0 $Y2=0
cc_493 N_A_758_306#_c_434_n N_A_1285_377#_c_1912_n 0.0067217f $X=6.35 $Y=1.81
+ $X2=0 $Y2=0
cc_494 N_A_758_306#_c_435_n N_A_1285_377#_c_1912_n 0.00177695f $X=6.8 $Y=1.81
+ $X2=0 $Y2=0
cc_495 N_A_758_306#_c_422_n N_VGND_c_2078_n 0.00251838f $X=6.315 $Y=1.365 $X2=0
+ $Y2=0
cc_496 N_A_758_306#_c_424_n N_VGND_c_2078_n 0.0300842f $X=5.11 $Y=0.515 $X2=0
+ $Y2=0
cc_497 N_A_758_306#_c_428_n N_VGND_c_2078_n 0.0217489f $X=6.035 $Y=1.53 $X2=0
+ $Y2=0
cc_498 N_A_758_306#_c_424_n N_VGND_c_2093_n 0.0112807f $X=5.11 $Y=0.515 $X2=0
+ $Y2=0
cc_499 N_A_758_306#_c_422_n N_VGND_c_2100_n 7.88433e-19 $X=6.315 $Y=1.365 $X2=0
+ $Y2=0
cc_500 N_A_758_306#_c_424_n N_VGND_c_2100_n 0.0083297f $X=5.11 $Y=0.515 $X2=0
+ $Y2=0
cc_501 N_A_758_306#_M1036_g N_A_299_126#_c_2325_n 0.0108159f $X=3.905 $Y=0.915
+ $X2=0 $Y2=0
cc_502 N_A_758_306#_M1042_g N_A_299_126#_c_2325_n 0.00124776f $X=4.335 $Y=0.915
+ $X2=0 $Y2=0
cc_503 N_A_758_306#_c_421_n N_A_299_126#_c_2325_n 0.0103225f $X=4.42 $Y=1.547
+ $X2=0 $Y2=0
cc_504 N_A_758_306#_M1036_g N_A_299_126#_c_2326_n 0.00848904f $X=3.905 $Y=0.915
+ $X2=0 $Y2=0
cc_505 N_A_758_306#_c_422_n N_A_1278_121#_c_2366_n 0.00749799f $X=6.315 $Y=1.365
+ $X2=0 $Y2=0
cc_506 N_A_758_306#_c_423_n N_A_1278_121#_c_2366_n 0.00699059f $X=6.745 $Y=1.365
+ $X2=0 $Y2=0
cc_507 N_A_758_306#_c_423_n N_A_1278_121#_c_2367_n 0.00163034f $X=6.745 $Y=1.365
+ $X2=0 $Y2=0
cc_508 N_S0_c_574_n N_A2_c_732_n 0.00720075f $X=8.155 $Y=1.56 $X2=0 $Y2=0
cc_509 N_S0_c_566_n N_A2_M1018_g 0.016973f $X=8.155 $Y=0.18 $X2=0 $Y2=0
cc_510 N_S0_c_569_n A2 0.00102397f $X=8.23 $Y=1.395 $X2=0 $Y2=0
cc_511 N_S0_c_574_n A2 2.4966e-19 $X=8.155 $Y=1.56 $X2=0 $Y2=0
cc_512 S0 A2 0.0225759f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_513 N_S0_c_569_n N_A2_c_737_n 0.00720075f $X=8.23 $Y=1.395 $X2=0 $Y2=0
cc_514 S0 N_A2_c_737_n 0.00383373f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_515 N_S0_c_578_n N_VPWR_c_1274_n 0.00121376f $X=2.93 $Y=1.885 $X2=0 $Y2=0
cc_516 N_S0_c_582_n N_VPWR_c_1275_n 0.0215552f $X=5.34 $Y=1.765 $X2=0 $Y2=0
cc_517 N_S0_c_578_n N_VPWR_c_1291_n 0.00279489f $X=2.93 $Y=1.885 $X2=0 $Y2=0
cc_518 N_S0_c_580_n N_VPWR_c_1291_n 0.00278271f $X=3.405 $Y=1.885 $X2=0 $Y2=0
cc_519 N_S0_c_582_n N_VPWR_c_1291_n 0.00413917f $X=5.34 $Y=1.765 $X2=0 $Y2=0
cc_520 N_S0_c_583_n N_VPWR_c_1292_n 8.16603e-19 $X=7.25 $Y=1.81 $X2=0 $Y2=0
cc_521 N_S0_c_584_n N_VPWR_c_1292_n 8.16603e-19 $X=7.7 $Y=1.81 $X2=0 $Y2=0
cc_522 N_S0_c_578_n N_VPWR_c_1270_n 0.00354316f $X=2.93 $Y=1.885 $X2=0 $Y2=0
cc_523 N_S0_c_580_n N_VPWR_c_1270_n 0.00354363f $X=3.405 $Y=1.885 $X2=0 $Y2=0
cc_524 N_S0_c_582_n N_VPWR_c_1270_n 0.00822528f $X=5.34 $Y=1.765 $X2=0 $Y2=0
cc_525 N_S0_c_578_n N_A_116_392#_c_1455_n 0.00377865f $X=2.93 $Y=1.885 $X2=0
+ $Y2=0
cc_526 N_S0_c_556_n N_A_116_392#_c_1456_n 0.00373913f $X=2.93 $Y=1.795 $X2=0
+ $Y2=0
cc_527 N_S0_c_578_n N_A_116_392#_c_1456_n 0.00250565f $X=2.93 $Y=1.885 $X2=0
+ $Y2=0
cc_528 N_S0_c_556_n N_A_116_392#_c_1451_n 0.0139099f $X=2.93 $Y=1.795 $X2=0
+ $Y2=0
cc_529 N_S0_c_560_n N_A_116_392#_c_1451_n 0.0170835f $X=3.405 $Y=1.795 $X2=0
+ $Y2=0
cc_530 N_S0_c_570_n N_A_116_392#_c_1451_n 0.00150122f $X=2.957 $Y=1.46 $X2=0
+ $Y2=0
cc_531 N_S0_c_571_n N_A_116_392#_c_1451_n 0.00150122f $X=3.432 $Y=1.46 $X2=0
+ $Y2=0
cc_532 N_S0_c_578_n N_A_296_392#_c_1515_n 0.0125185f $X=2.93 $Y=1.885 $X2=0
+ $Y2=0
cc_533 N_S0_c_578_n N_A_296_392#_c_1516_n 0.0107603f $X=2.93 $Y=1.885 $X2=0
+ $Y2=0
cc_534 N_S0_c_580_n N_A_296_392#_c_1516_n 2.22151e-19 $X=3.405 $Y=1.885 $X2=0
+ $Y2=0
cc_535 N_S0_c_578_n N_A_296_392#_c_1524_n 0.00127391f $X=2.93 $Y=1.885 $X2=0
+ $Y2=0
cc_536 N_S0_c_578_n N_A_509_392#_c_1557_n 0.00909697f $X=2.93 $Y=1.885 $X2=0
+ $Y2=0
cc_537 N_S0_c_580_n N_A_509_392#_c_1557_n 0.0134615f $X=3.405 $Y=1.885 $X2=0
+ $Y2=0
cc_538 N_S0_M1004_g N_A_509_392#_c_1545_n 0.0125911f $X=3 $Y=0.915 $X2=0 $Y2=0
cc_539 N_S0_c_558_n N_A_509_392#_c_1545_n 0.0034051f $X=3.4 $Y=0.18 $X2=0 $Y2=0
cc_540 N_S0_M1047_g N_A_509_392#_c_1545_n 0.0165579f $X=3.475 $Y=0.915 $X2=0
+ $Y2=0
cc_541 N_S0_M1047_g N_A_509_392#_c_1546_n 0.00505756f $X=3.475 $Y=0.915 $X2=0
+ $Y2=0
cc_542 N_S0_c_562_n N_A_509_392#_c_1547_n 0.01748f $X=5.25 $Y=0.18 $X2=0 $Y2=0
cc_543 N_S0_M1012_g N_A_509_392#_c_1547_n 0.00174103f $X=5.325 $Y=0.74 $X2=0
+ $Y2=0
cc_544 N_S0_c_582_n N_A_509_392#_c_1559_n 0.00279287f $X=5.34 $Y=1.765 $X2=0
+ $Y2=0
cc_545 N_S0_c_578_n N_A_509_392#_c_1561_n 0.00673207f $X=2.93 $Y=1.885 $X2=0
+ $Y2=0
cc_546 N_S0_c_580_n N_A_509_392#_c_1561_n 5.40419e-19 $X=3.405 $Y=1.885 $X2=0
+ $Y2=0
cc_547 N_S0_M1004_g N_A_509_392#_c_1551_n 0.009152f $X=3 $Y=0.915 $X2=0 $Y2=0
cc_548 N_S0_c_562_n N_A_509_392#_c_1552_n 0.00470837f $X=5.25 $Y=0.18 $X2=0
+ $Y2=0
cc_549 N_S0_c_582_n N_A_509_392#_c_1563_n 0.00761327f $X=5.34 $Y=1.765 $X2=0
+ $Y2=0
cc_550 S0 N_A_509_392#_c_1563_n 0.00940257f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_551 N_S0_M1012_g N_A_1191_121#_c_1733_n 0.00179375f $X=5.325 $Y=0.74 $X2=0
+ $Y2=0
cc_552 N_S0_c_564_n N_A_1191_121#_c_1733_n 2.94405e-19 $X=5.34 $Y=1.275 $X2=0
+ $Y2=0
cc_553 N_S0_M1012_g N_A_1191_121#_c_1734_n 8.46248e-19 $X=5.325 $Y=0.74 $X2=0
+ $Y2=0
cc_554 N_S0_c_566_n N_A_1191_121#_c_1734_n 0.00494503f $X=8.155 $Y=0.18 $X2=0
+ $Y2=0
cc_555 N_S0_c_582_n N_A_1191_121#_c_1744_n 0.00145255f $X=5.34 $Y=1.765 $X2=0
+ $Y2=0
cc_556 N_S0_M1006_g N_A_1191_121#_c_1735_n 6.552e-19 $X=7.175 $Y=0.925 $X2=0
+ $Y2=0
cc_557 N_S0_M1006_g N_A_1191_121#_c_1782_n 0.00407014f $X=7.175 $Y=0.925 $X2=0
+ $Y2=0
cc_558 N_S0_M1040_g N_A_1191_121#_c_1782_n 4.70674e-19 $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_559 N_S0_M1006_g N_A_1191_121#_c_1736_n 0.00313646f $X=7.175 $Y=0.925 $X2=0
+ $Y2=0
cc_560 N_S0_c_583_n N_A_1191_121#_c_1736_n 0.0013323f $X=7.25 $Y=1.81 $X2=0
+ $Y2=0
cc_561 N_S0_M1040_g N_A_1191_121#_c_1736_n 6.31438e-19 $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_562 S0 N_A_1191_121#_c_1736_n 0.0267619f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_563 N_S0_c_576_n N_A_1191_121#_c_1736_n 0.00802909f $X=7.79 $Y=1.56 $X2=0
+ $Y2=0
cc_564 N_S0_M1006_g N_A_1191_121#_c_1737_n 0.0103465f $X=7.175 $Y=0.925 $X2=0
+ $Y2=0
cc_565 N_S0_M1040_g N_A_1191_121#_c_1737_n 0.00968335f $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_566 N_S0_c_583_n N_A_1191_121#_c_1747_n 0.0163197f $X=7.25 $Y=1.81 $X2=0
+ $Y2=0
cc_567 N_S0_c_584_n N_A_1191_121#_c_1747_n 0.00846974f $X=7.7 $Y=1.81 $X2=0
+ $Y2=0
cc_568 N_S0_c_574_n N_A_1191_121#_c_1747_n 0.00305792f $X=8.155 $Y=1.56 $X2=0
+ $Y2=0
cc_569 S0 N_A_1191_121#_c_1747_n 0.0792113f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_570 N_S0_c_576_n N_A_1191_121#_c_1747_n 0.00148072f $X=7.79 $Y=1.56 $X2=0
+ $Y2=0
cc_571 N_S0_M1006_g N_A_1191_121#_c_1741_n 0.00265737f $X=7.175 $Y=0.925 $X2=0
+ $Y2=0
cc_572 N_S0_c_583_n N_A_1191_121#_c_1752_n 6.14512e-19 $X=7.25 $Y=1.81 $X2=0
+ $Y2=0
cc_573 N_S0_M1040_g N_A_1191_121#_c_1742_n 5.15987e-19 $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_574 N_S0_c_569_n N_A_1191_121#_c_1742_n 0.00476489f $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_575 N_S0_c_583_n N_A_1285_377#_c_1915_n 9.00086e-19 $X=7.25 $Y=1.81 $X2=0
+ $Y2=0
cc_576 N_S0_c_583_n N_A_1285_377#_c_1911_n 0.012727f $X=7.25 $Y=1.81 $X2=0 $Y2=0
cc_577 N_S0_c_584_n N_A_1285_377#_c_1911_n 0.0105678f $X=7.7 $Y=1.81 $X2=0 $Y2=0
cc_578 N_S0_c_584_n N_A_1285_377#_c_1914_n 0.00833356f $X=7.7 $Y=1.81 $X2=0
+ $Y2=0
cc_579 N_S0_c_584_n N_A_1465_377#_c_1968_n 0.012095f $X=7.7 $Y=1.81 $X2=0 $Y2=0
cc_580 N_S0_c_583_n N_A_1465_377#_c_1970_n 0.00566403f $X=7.25 $Y=1.81 $X2=0
+ $Y2=0
cc_581 N_S0_c_584_n N_A_1465_377#_c_1970_n 0.0108408f $X=7.7 $Y=1.81 $X2=0 $Y2=0
cc_582 N_S0_c_559_n N_VGND_c_2077_n 0.00227104f $X=3.075 $Y=0.18 $X2=0 $Y2=0
cc_583 N_S0_M1012_g N_VGND_c_2078_n 0.0147983f $X=5.325 $Y=0.74 $X2=0 $Y2=0
cc_584 N_S0_c_564_n N_VGND_c_2078_n 9.58393e-19 $X=5.34 $Y=1.275 $X2=0 $Y2=0
cc_585 N_S0_c_566_n N_VGND_c_2078_n 0.0187754f $X=8.155 $Y=0.18 $X2=0 $Y2=0
cc_586 N_S0_c_573_n N_VGND_c_2078_n 0.00460513f $X=5.325 $Y=0.18 $X2=0 $Y2=0
cc_587 N_S0_c_566_n N_VGND_c_2086_n 0.00443934f $X=8.155 $Y=0.18 $X2=0 $Y2=0
cc_588 N_S0_c_569_n N_VGND_c_2086_n 6.29386e-19 $X=8.23 $Y=1.395 $X2=0 $Y2=0
cc_589 N_S0_c_566_n N_VGND_c_2087_n 0.0604235f $X=8.155 $Y=0.18 $X2=0 $Y2=0
cc_590 N_S0_c_559_n N_VGND_c_2093_n 0.0586296f $X=3.075 $Y=0.18 $X2=0 $Y2=0
cc_591 N_S0_c_558_n N_VGND_c_2100_n 0.00777952f $X=3.4 $Y=0.18 $X2=0 $Y2=0
cc_592 N_S0_c_559_n N_VGND_c_2100_n 0.00604517f $X=3.075 $Y=0.18 $X2=0 $Y2=0
cc_593 N_S0_c_562_n N_VGND_c_2100_n 0.0489771f $X=5.25 $Y=0.18 $X2=0 $Y2=0
cc_594 N_S0_c_566_n N_VGND_c_2100_n 0.0737993f $X=8.155 $Y=0.18 $X2=0 $Y2=0
cc_595 N_S0_c_572_n N_VGND_c_2100_n 0.00370846f $X=3.475 $Y=0.18 $X2=0 $Y2=0
cc_596 N_S0_c_573_n N_VGND_c_2100_n 0.00749832f $X=5.325 $Y=0.18 $X2=0 $Y2=0
cc_597 N_S0_M1004_g N_A_114_126#_c_2289_n 0.0155442f $X=3 $Y=0.915 $X2=0 $Y2=0
cc_598 N_S0_c_571_n N_A_114_126#_c_2289_n 3.37014e-19 $X=3.432 $Y=1.46 $X2=0
+ $Y2=0
cc_599 N_S0_M1004_g N_A_114_126#_c_2279_n 0.00991756f $X=3 $Y=0.915 $X2=0 $Y2=0
cc_600 N_S0_c_570_n N_A_114_126#_c_2279_n 3.26692e-19 $X=2.957 $Y=1.46 $X2=0
+ $Y2=0
cc_601 N_S0_M1004_g N_A_299_126#_c_2325_n 0.00490473f $X=3 $Y=0.915 $X2=0 $Y2=0
cc_602 N_S0_M1047_g N_A_299_126#_c_2325_n 0.00850432f $X=3.475 $Y=0.915 $X2=0
+ $Y2=0
cc_603 N_S0_c_570_n N_A_299_126#_c_2325_n 0.00997967f $X=2.957 $Y=1.46 $X2=0
+ $Y2=0
cc_604 N_S0_c_571_n N_A_299_126#_c_2325_n 0.00925259f $X=3.432 $Y=1.46 $X2=0
+ $Y2=0
cc_605 N_S0_M1047_g N_A_299_126#_c_2326_n 9.78227e-19 $X=3.475 $Y=0.915 $X2=0
+ $Y2=0
cc_606 N_S0_M1004_g N_A_299_126#_c_2328_n 0.00440371f $X=3 $Y=0.915 $X2=0 $Y2=0
cc_607 N_S0_c_570_n N_A_299_126#_c_2328_n 6.41487e-19 $X=2.957 $Y=1.46 $X2=0
+ $Y2=0
cc_608 N_S0_M1006_g N_A_1278_121#_c_2366_n 6.67018e-19 $X=7.175 $Y=0.925 $X2=0
+ $Y2=0
cc_609 N_S0_c_566_n N_A_1278_121#_c_2367_n 0.0264241f $X=8.155 $Y=0.18 $X2=0
+ $Y2=0
cc_610 N_S0_M1006_g N_A_1278_121#_c_2367_n 0.00115636f $X=7.175 $Y=0.925 $X2=0
+ $Y2=0
cc_611 N_S0_M1040_g N_A_1278_121#_c_2367_n 0.00115673f $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_612 N_S0_c_569_n N_A_1278_121#_c_2367_n 0.00580058f $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_613 N_S0_c_566_n N_A_1278_121#_c_2368_n 0.00727301f $X=8.155 $Y=0.18 $X2=0
+ $Y2=0
cc_614 N_S0_M1040_g N_A_1278_121#_c_2369_n 5.73967e-19 $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_615 N_S0_c_569_n N_A_1278_121#_c_2369_n 0.0068488f $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_616 N_S0_c_569_n N_A_1278_121#_c_2371_n 0.00783294f $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_617 N_S0_M1040_g N_A_1450_121#_c_2419_n 0.00950725f $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_618 N_S0_c_569_n N_A_1450_121#_c_2419_n 0.0012418f $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_619 S0 N_A_1450_121#_c_2419_n 0.0446554f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_620 N_S0_c_576_n N_A_1450_121#_c_2419_n 0.00694924f $X=7.79 $Y=1.56 $X2=0
+ $Y2=0
cc_621 N_S0_c_569_n N_A_1450_121#_c_2420_n 0.0010042f $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_622 S0 N_A_1450_121#_c_2420_n 0.00925546f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_623 N_S0_M1040_g N_A_1450_121#_c_2422_n 0.00485385f $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_624 N_S0_c_569_n N_A_1450_121#_c_2422_n 5.67881e-19 $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_625 S0 N_A_1450_121#_c_2422_n 0.0196697f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_626 N_S0_c_576_n N_A_1450_121#_c_2422_n 0.00239105f $X=7.79 $Y=1.56 $X2=0
+ $Y2=0
cc_627 N_S0_M1040_g N_A_1450_121#_c_2423_n 7.7137e-19 $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_628 N_S0_c_569_n N_A_1450_121#_c_2423_n 0.0153513f $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_629 S0 N_A_1450_121#_c_2423_n 0.0129022f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_630 N_A2_M1038_g N_A3_M1014_g 0.0219085f $X=9.385 $Y=0.69 $X2=0 $Y2=0
cc_631 A2 N_A3_M1014_g 0.00454402f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_632 N_A2_c_741_n N_A3_c_799_n 0.0287768f $X=9.245 $Y=1.885 $X2=0 $Y2=0
cc_633 N_A2_c_734_n A3 6.45648e-19 $X=9.245 $Y=1.795 $X2=0 $Y2=0
cc_634 A2 A3 0.0235668f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_635 N_A2_c_737_n A3 6.12354e-19 $X=9.385 $Y=1.425 $X2=0 $Y2=0
cc_636 N_A2_c_734_n N_A3_c_798_n 0.00878274f $X=9.245 $Y=1.795 $X2=0 $Y2=0
cc_637 A2 N_A3_c_798_n 0.00144227f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_638 N_A2_c_737_n N_A3_c_798_n 0.0219085f $X=9.385 $Y=1.425 $X2=0 $Y2=0
cc_639 N_A2_c_741_n N_VPWR_c_1281_n 0.00361052f $X=9.245 $Y=1.885 $X2=0 $Y2=0
cc_640 N_A2_c_739_n N_VPWR_c_1282_n 0.00314961f $X=8.795 $Y=1.885 $X2=0 $Y2=0
cc_641 N_A2_c_741_n N_VPWR_c_1282_n 0.00314961f $X=9.245 $Y=1.885 $X2=0 $Y2=0
cc_642 N_A2_c_739_n N_VPWR_c_1297_n 0.0051324f $X=8.795 $Y=1.885 $X2=0 $Y2=0
cc_643 N_A2_c_739_n N_VPWR_c_1270_n 0.00395154f $X=8.795 $Y=1.885 $X2=0 $Y2=0
cc_644 N_A2_c_741_n N_VPWR_c_1270_n 0.00391819f $X=9.245 $Y=1.885 $X2=0 $Y2=0
cc_645 A2 N_A_509_392#_c_1563_n 0.00557945f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_646 N_A2_c_739_n N_A_1191_121#_c_1747_n 0.0151577f $X=8.795 $Y=1.885 $X2=0
+ $Y2=0
cc_647 N_A2_c_741_n N_A_1191_121#_c_1747_n 0.0139074f $X=9.245 $Y=1.885 $X2=0
+ $Y2=0
cc_648 A2 N_A_1191_121#_c_1747_n 0.0505729f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_649 N_A2_c_737_n N_A_1191_121#_c_1747_n 9.6499e-19 $X=9.385 $Y=1.425 $X2=0
+ $Y2=0
cc_650 N_A2_c_739_n N_A_1285_377#_c_1913_n 0.0131108f $X=8.795 $Y=1.885 $X2=0
+ $Y2=0
cc_651 N_A2_c_741_n N_A_1285_377#_c_1913_n 0.0143307f $X=9.245 $Y=1.885 $X2=0
+ $Y2=0
cc_652 N_A2_c_741_n N_A_1285_377#_c_1926_n 0.00147616f $X=9.245 $Y=1.885 $X2=0
+ $Y2=0
cc_653 N_A2_c_739_n N_A_1285_377#_c_1914_n 0.00432465f $X=8.795 $Y=1.885 $X2=0
+ $Y2=0
cc_654 N_A2_c_739_n N_A_1465_377#_c_1968_n 0.0104079f $X=8.795 $Y=1.885 $X2=0
+ $Y2=0
cc_655 N_A2_c_741_n N_A_1465_377#_c_1968_n 0.00412569f $X=9.245 $Y=1.885 $X2=0
+ $Y2=0
cc_656 N_A2_M1018_g N_VGND_c_2079_n 4.68597e-19 $X=8.955 $Y=0.69 $X2=0 $Y2=0
cc_657 N_A2_M1038_g N_VGND_c_2079_n 0.00822569f $X=9.385 $Y=0.69 $X2=0 $Y2=0
cc_658 N_A2_M1018_g N_VGND_c_2086_n 0.00240369f $X=8.955 $Y=0.69 $X2=0 $Y2=0
cc_659 N_A2_M1018_g N_VGND_c_2088_n 0.00316493f $X=8.955 $Y=0.69 $X2=0 $Y2=0
cc_660 N_A2_M1038_g N_VGND_c_2088_n 0.00383152f $X=9.385 $Y=0.69 $X2=0 $Y2=0
cc_661 N_A2_M1018_g N_VGND_c_2100_n 0.00394055f $X=8.955 $Y=0.69 $X2=0 $Y2=0
cc_662 N_A2_M1038_g N_VGND_c_2100_n 0.0075754f $X=9.385 $Y=0.69 $X2=0 $Y2=0
cc_663 N_A2_M1018_g N_A_1278_121#_c_2367_n 5.24269e-19 $X=8.955 $Y=0.69 $X2=0
+ $Y2=0
cc_664 N_A2_M1018_g N_A_1278_121#_c_2369_n 0.00226665f $X=8.955 $Y=0.69 $X2=0
+ $Y2=0
cc_665 N_A2_M1018_g N_A_1278_121#_c_2370_n 0.00981813f $X=8.955 $Y=0.69 $X2=0
+ $Y2=0
cc_666 N_A2_M1018_g N_A_1278_121#_c_2372_n 0.00953282f $X=8.955 $Y=0.69 $X2=0
+ $Y2=0
cc_667 N_A2_M1018_g N_A_1450_121#_c_2420_n 0.0115689f $X=8.955 $Y=0.69 $X2=0
+ $Y2=0
cc_668 N_A2_M1038_g N_A_1450_121#_c_2420_n 0.0142932f $X=9.385 $Y=0.69 $X2=0
+ $Y2=0
cc_669 A2 N_A_1450_121#_c_2420_n 0.054183f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_670 N_A2_c_737_n N_A_1450_121#_c_2420_n 0.00812717f $X=9.385 $Y=1.425 $X2=0
+ $Y2=0
cc_671 N_A2_M1038_g N_A_1450_121#_c_2421_n 9.61031e-19 $X=9.385 $Y=0.69 $X2=0
+ $Y2=0
cc_672 N_A2_M1018_g N_A_1450_121#_c_2423_n 0.00262376f $X=8.955 $Y=0.69 $X2=0
+ $Y2=0
cc_673 N_A3_c_800_n N_VPWR_c_1276_n 0.00675985f $X=10.325 $Y=1.885 $X2=0 $Y2=0
cc_674 N_A3_c_799_n N_VPWR_c_1281_n 0.00332626f $X=9.875 $Y=1.885 $X2=0 $Y2=0
cc_675 N_A3_c_799_n N_VPWR_c_1283_n 0.00312616f $X=9.875 $Y=1.885 $X2=0 $Y2=0
cc_676 N_A3_c_800_n N_VPWR_c_1283_n 0.00444469f $X=10.325 $Y=1.885 $X2=0 $Y2=0
cc_677 N_A3_c_799_n N_VPWR_c_1270_n 0.0038866f $X=9.875 $Y=1.885 $X2=0 $Y2=0
cc_678 N_A3_c_800_n N_VPWR_c_1270_n 0.00858722f $X=10.325 $Y=1.885 $X2=0 $Y2=0
cc_679 A3 N_A_509_392#_c_1563_n 0.00519452f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_680 N_A3_c_799_n N_A_1191_121#_c_1747_n 0.0130063f $X=9.875 $Y=1.885 $X2=0
+ $Y2=0
cc_681 N_A3_c_800_n N_A_1191_121#_c_1747_n 0.0166408f $X=10.325 $Y=1.885 $X2=0
+ $Y2=0
cc_682 A3 N_A_1191_121#_c_1747_n 0.0475163f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_683 N_A3_c_798_n N_A_1191_121#_c_1747_n 0.00932914f $X=10.325 $Y=1.665 $X2=0
+ $Y2=0
cc_684 N_A3_c_794_n N_A_1191_121#_c_1738_n 0.00188304f $X=10.245 $Y=1.085 $X2=0
+ $Y2=0
cc_685 N_A3_c_800_n N_A_1191_121#_c_1738_n 0.00173042f $X=10.325 $Y=1.885 $X2=0
+ $Y2=0
cc_686 N_A3_c_796_n N_A_1191_121#_c_1738_n 0.0108756f $X=10.335 $Y=1.16 $X2=0
+ $Y2=0
cc_687 A3 N_A_1191_121#_c_1738_n 0.0196213f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_688 N_A3_c_798_n N_A_1191_121#_c_1738_n 0.00534737f $X=10.325 $Y=1.665 $X2=0
+ $Y2=0
cc_689 N_A3_c_800_n N_A_1191_121#_c_1749_n 0.00500195f $X=10.325 $Y=1.885 $X2=0
+ $Y2=0
cc_690 N_A3_c_794_n N_A_1191_121#_c_1739_n 6.63977e-19 $X=10.245 $Y=1.085 $X2=0
+ $Y2=0
cc_691 N_A3_c_799_n N_A_1285_377#_c_1913_n 0.0149608f $X=9.875 $Y=1.885 $X2=0
+ $Y2=0
cc_692 N_A3_c_800_n N_A_1285_377#_c_1913_n 0.00415864f $X=10.325 $Y=1.885 $X2=0
+ $Y2=0
cc_693 N_A3_c_799_n N_A_1285_377#_c_1926_n 0.007143f $X=9.875 $Y=1.885 $X2=0
+ $Y2=0
cc_694 N_A3_c_800_n N_A_1285_377#_c_1926_n 0.0038234f $X=10.325 $Y=1.885 $X2=0
+ $Y2=0
cc_695 N_A3_c_799_n N_A_1465_377#_c_1968_n 7.25313e-19 $X=9.875 $Y=1.885 $X2=0
+ $Y2=0
cc_696 N_A3_M1014_g N_VGND_c_2079_n 0.00160688f $X=9.815 $Y=0.69 $X2=0 $Y2=0
cc_697 N_A3_M1014_g N_VGND_c_2080_n 0.00434272f $X=9.815 $Y=0.69 $X2=0 $Y2=0
cc_698 N_A3_c_794_n N_VGND_c_2080_n 0.00383152f $X=10.245 $Y=1.085 $X2=0 $Y2=0
cc_699 N_A3_M1014_g N_VGND_c_2081_n 5.59381e-19 $X=9.815 $Y=0.69 $X2=0 $Y2=0
cc_700 N_A3_c_794_n N_VGND_c_2081_n 0.0129152f $X=10.245 $Y=1.085 $X2=0 $Y2=0
cc_701 N_A3_c_796_n N_VGND_c_2081_n 0.00323003f $X=10.335 $Y=1.16 $X2=0 $Y2=0
cc_702 A3 N_VGND_c_2081_n 0.00601406f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_703 N_A3_M1014_g N_VGND_c_2100_n 0.00820382f $X=9.815 $Y=0.69 $X2=0 $Y2=0
cc_704 N_A3_c_794_n N_VGND_c_2100_n 0.0075754f $X=10.245 $Y=1.085 $X2=0 $Y2=0
cc_705 N_A3_M1014_g N_A_1450_121#_c_2420_n 0.0135496f $X=9.815 $Y=0.69 $X2=0
+ $Y2=0
cc_706 N_A3_c_794_n N_A_1450_121#_c_2420_n 0.00109283f $X=10.245 $Y=1.085 $X2=0
+ $Y2=0
cc_707 A3 N_A_1450_121#_c_2420_n 0.0177215f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_708 N_A3_c_798_n N_A_1450_121#_c_2420_n 0.00281218f $X=10.325 $Y=1.665 $X2=0
+ $Y2=0
cc_709 N_A3_M1014_g N_A_1450_121#_c_2421_n 0.00754481f $X=9.815 $Y=0.69 $X2=0
+ $Y2=0
cc_710 N_S1_c_866_n N_A_2489_347#_c_980_n 0.02595f $X=12.035 $Y=1.885 $X2=0
+ $Y2=0
cc_711 N_S1_M1015_g N_A_2489_347#_M1009_g 0.00828914f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_712 N_S1_c_858_n N_A_2489_347#_M1009_g 0.00438971f $X=13.54 $Y=1.215 $X2=0
+ $Y2=0
cc_713 N_S1_c_859_n N_A_2489_347#_M1009_g 0.0182158f $X=12.315 $Y=1.36 $X2=0
+ $Y2=0
cc_714 N_S1_c_862_n N_A_2489_347#_M1009_g 0.0109898f $X=12.835 $Y=1.455 $X2=0
+ $Y2=0
cc_715 N_S1_c_858_n N_A_2489_347#_M1048_g 0.01631f $X=13.54 $Y=1.215 $X2=0 $Y2=0
cc_716 N_S1_c_860_n N_A_2489_347#_M1048_g 0.0145818f $X=13.87 $Y=1.385 $X2=0
+ $Y2=0
cc_717 N_S1_c_862_n N_A_2489_347#_M1048_g 9.7513e-19 $X=12.835 $Y=1.455 $X2=0
+ $Y2=0
cc_718 N_S1_c_858_n N_A_2489_347#_c_982_n 0.0333171f $X=13.54 $Y=1.215 $X2=0
+ $Y2=0
cc_719 N_S1_c_860_n N_A_2489_347#_c_982_n 0.00250238f $X=13.87 $Y=1.385 $X2=0
+ $Y2=0
cc_720 N_S1_c_868_n N_A_2489_347#_c_983_n 0.00145993f $X=14.3 $Y=1.765 $X2=0
+ $Y2=0
cc_721 N_S1_c_853_n N_A_2489_347#_c_976_n 0.0209844f $X=14.21 $Y=1.37 $X2=0
+ $Y2=0
cc_722 N_S1_c_854_n N_A_2489_347#_c_976_n 0.00537771f $X=14.285 $Y=1.22 $X2=0
+ $Y2=0
cc_723 N_S1_c_855_n N_A_2489_347#_c_976_n 0.00632146f $X=14.3 $Y=1.675 $X2=0
+ $Y2=0
cc_724 N_S1_c_858_n N_A_2489_347#_c_976_n 0.0307762f $X=13.54 $Y=1.215 $X2=0
+ $Y2=0
cc_725 N_S1_c_860_n N_A_2489_347#_c_976_n 2.10237e-19 $X=13.87 $Y=1.385 $X2=0
+ $Y2=0
cc_726 N_S1_c_858_n N_A_2489_347#_c_977_n 0.0293493f $X=13.54 $Y=1.215 $X2=0
+ $Y2=0
cc_727 N_S1_c_860_n N_A_2489_347#_c_977_n 3.06382e-19 $X=13.87 $Y=1.385 $X2=0
+ $Y2=0
cc_728 N_S1_c_862_n N_A_2489_347#_c_977_n 0.0246532f $X=12.835 $Y=1.455 $X2=0
+ $Y2=0
cc_729 N_S1_c_852_n N_A_2489_347#_c_978_n 0.00888992f $X=12.035 $Y=1.795 $X2=0
+ $Y2=0
cc_730 N_S1_c_858_n N_A_2489_347#_c_978_n 0.00280142f $X=13.54 $Y=1.215 $X2=0
+ $Y2=0
cc_731 N_S1_c_859_n N_A_2489_347#_c_978_n 0.00227232f $X=12.315 $Y=1.36 $X2=0
+ $Y2=0
cc_732 N_S1_c_860_n N_A_2489_347#_c_978_n 0.00530331f $X=13.87 $Y=1.385 $X2=0
+ $Y2=0
cc_733 N_S1_c_861_n N_A_2489_347#_c_978_n 0.0096783f $X=12.665 $Y=1.455 $X2=0
+ $Y2=0
cc_734 N_S1_c_862_n N_A_2489_347#_c_978_n 0.0159807f $X=12.835 $Y=1.455 $X2=0
+ $Y2=0
cc_735 N_S1_c_853_n N_A_2489_347#_c_987_n 0.00681687f $X=14.21 $Y=1.37 $X2=0
+ $Y2=0
cc_736 N_S1_c_868_n N_A_2489_347#_c_987_n 0.00506949f $X=14.3 $Y=1.765 $X2=0
+ $Y2=0
cc_737 N_S1_c_853_n N_A_2489_347#_c_979_n 0.00474764f $X=14.21 $Y=1.37 $X2=0
+ $Y2=0
cc_738 N_S1_c_868_n N_A_2199_74#_c_1079_n 0.0191387f $X=14.3 $Y=1.765 $X2=0
+ $Y2=0
cc_739 N_S1_c_854_n N_A_2199_74#_M1016_g 0.00759404f $X=14.285 $Y=1.22 $X2=0
+ $Y2=0
cc_740 N_S1_c_857_n N_A_2199_74#_M1016_g 0.00421747f $X=14.3 $Y=1.37 $X2=0 $Y2=0
cc_741 N_S1_M1013_g N_A_2199_74#_c_1066_n 0.00631046f $X=11.355 $Y=0.69 $X2=0
+ $Y2=0
cc_742 N_S1_c_850_n N_A_2199_74#_c_1066_n 0.00843503f $X=11.535 $Y=1.795 $X2=0
+ $Y2=0
cc_743 N_S1_c_864_n N_A_2199_74#_c_1066_n 0.0146742f $X=11.535 $Y=1.885 $X2=0
+ $Y2=0
cc_744 N_S1_c_852_n N_A_2199_74#_c_1066_n 2.39988e-19 $X=12.035 $Y=1.795 $X2=0
+ $Y2=0
cc_745 N_S1_c_866_n N_A_2199_74#_c_1066_n 6.80971e-19 $X=12.035 $Y=1.885 $X2=0
+ $Y2=0
cc_746 N_S1_c_856_n N_A_2199_74#_c_1066_n 0.0182011f $X=12.125 $Y=1.36 $X2=0
+ $Y2=0
cc_747 N_S1_c_864_n N_A_2199_74#_c_1098_n 0.00917562f $X=11.535 $Y=1.885 $X2=0
+ $Y2=0
cc_748 N_S1_c_866_n N_A_2199_74#_c_1098_n 0.0153402f $X=12.035 $Y=1.885 $X2=0
+ $Y2=0
cc_749 N_S1_c_864_n N_A_2199_74#_c_1084_n 4.09683e-19 $X=11.535 $Y=1.885 $X2=0
+ $Y2=0
cc_750 N_S1_c_866_n N_A_2199_74#_c_1085_n 0.00152337f $X=12.035 $Y=1.885 $X2=0
+ $Y2=0
cc_751 N_S1_c_859_n N_A_2199_74#_c_1085_n 0.00151241f $X=12.315 $Y=1.36 $X2=0
+ $Y2=0
cc_752 N_S1_c_861_n N_A_2199_74#_c_1085_n 0.0294528f $X=12.665 $Y=1.455 $X2=0
+ $Y2=0
cc_753 N_S1_c_859_n N_A_2199_74#_c_1067_n 5.84221e-19 $X=12.315 $Y=1.36 $X2=0
+ $Y2=0
cc_754 N_S1_c_861_n N_A_2199_74#_c_1105_n 0.0171013f $X=12.665 $Y=1.455 $X2=0
+ $Y2=0
cc_755 N_S1_c_854_n N_A_2199_74#_c_1069_n 0.00475331f $X=14.285 $Y=1.22 $X2=0
+ $Y2=0
cc_756 N_S1_c_858_n N_A_2199_74#_c_1069_n 0.0274492f $X=13.54 $Y=1.215 $X2=0
+ $Y2=0
cc_757 N_S1_c_860_n N_A_2199_74#_c_1069_n 8.35195e-19 $X=13.87 $Y=1.385 $X2=0
+ $Y2=0
cc_758 N_S1_c_854_n N_A_2199_74#_c_1070_n 0.0160644f $X=14.285 $Y=1.22 $X2=0
+ $Y2=0
cc_759 N_S1_c_854_n N_A_2199_74#_c_1071_n 0.00694011f $X=14.285 $Y=1.22 $X2=0
+ $Y2=0
cc_760 N_S1_c_857_n N_A_2199_74#_c_1071_n 0.00251159f $X=14.3 $Y=1.37 $X2=0
+ $Y2=0
cc_761 N_S1_c_855_n N_A_2199_74#_c_1072_n 0.00276866f $X=14.3 $Y=1.675 $X2=0
+ $Y2=0
cc_762 N_S1_c_857_n N_A_2199_74#_c_1072_n 0.00746893f $X=14.3 $Y=1.37 $X2=0
+ $Y2=0
cc_763 N_S1_M1013_g N_A_2199_74#_c_1074_n 0.0123838f $X=11.355 $Y=0.69 $X2=0
+ $Y2=0
cc_764 N_S1_M1015_g N_A_2199_74#_c_1074_n 4.89925e-19 $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_765 N_S1_M1015_g N_A_2199_74#_c_1116_n 0.00816632f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_766 N_S1_c_856_n N_A_2199_74#_c_1116_n 0.00448287f $X=12.125 $Y=1.36 $X2=0
+ $Y2=0
cc_767 N_S1_M1013_g N_A_2199_74#_c_1075_n 8.90513e-19 $X=11.355 $Y=0.69 $X2=0
+ $Y2=0
cc_768 N_S1_M1015_g N_A_2199_74#_c_1075_n 0.00988861f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_769 N_S1_c_857_n N_A_2199_74#_c_1078_n 0.0107014f $X=14.3 $Y=1.37 $X2=0 $Y2=0
cc_770 N_S1_c_868_n N_VPWR_c_1277_n 0.0043835f $X=14.3 $Y=1.765 $X2=0 $Y2=0
cc_771 N_S1_c_864_n N_VPWR_c_1285_n 0.00278271f $X=11.535 $Y=1.885 $X2=0 $Y2=0
cc_772 N_S1_c_866_n N_VPWR_c_1285_n 0.00278271f $X=12.035 $Y=1.885 $X2=0 $Y2=0
cc_773 N_S1_c_868_n N_VPWR_c_1285_n 0.00460063f $X=14.3 $Y=1.765 $X2=0 $Y2=0
cc_774 N_S1_c_864_n N_VPWR_c_1270_n 0.00359085f $X=11.535 $Y=1.885 $X2=0 $Y2=0
cc_775 N_S1_c_866_n N_VPWR_c_1270_n 0.00354798f $X=12.035 $Y=1.885 $X2=0 $Y2=0
cc_776 N_S1_c_868_n N_VPWR_c_1270_n 0.00912933f $X=14.3 $Y=1.765 $X2=0 $Y2=0
cc_777 N_S1_M1015_g N_A_509_392#_c_1549_n 0.00609692f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_778 N_S1_c_856_n N_A_509_392#_c_1549_n 0.0100662f $X=12.125 $Y=1.36 $X2=0
+ $Y2=0
cc_779 N_S1_c_861_n N_A_509_392#_c_1549_n 0.0135925f $X=12.665 $Y=1.455 $X2=0
+ $Y2=0
cc_780 N_S1_M1013_g N_A_509_392#_c_1550_n 6.78751e-19 $X=11.355 $Y=0.69 $X2=0
+ $Y2=0
cc_781 N_S1_M1015_g N_A_509_392#_c_1550_n 0.00528673f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_782 N_S1_c_861_n N_A_509_392#_c_1630_n 0.00877217f $X=12.665 $Y=1.455 $X2=0
+ $Y2=0
cc_783 N_S1_c_862_n N_A_509_392#_c_1630_n 0.0128809f $X=12.835 $Y=1.455 $X2=0
+ $Y2=0
cc_784 N_S1_M1015_g N_A_509_392#_c_1554_n 0.00323735f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_785 N_S1_c_859_n N_A_509_392#_c_1554_n 0.00385917f $X=12.315 $Y=1.36 $X2=0
+ $Y2=0
cc_786 N_S1_c_861_n N_A_509_392#_c_1554_n 0.0137977f $X=12.665 $Y=1.455 $X2=0
+ $Y2=0
cc_787 N_S1_c_858_n N_A_509_392#_c_1635_n 0.0196914f $X=13.54 $Y=1.215 $X2=0
+ $Y2=0
cc_788 N_S1_c_864_n N_A_509_392#_c_1563_n 0.00803139f $X=11.535 $Y=1.885 $X2=0
+ $Y2=0
cc_789 N_S1_c_864_n N_A_509_392#_c_1566_n 0.00191803f $X=11.535 $Y=1.885 $X2=0
+ $Y2=0
cc_790 N_S1_M1013_g N_A_509_392#_c_1555_n 3.16363e-19 $X=11.355 $Y=0.69 $X2=0
+ $Y2=0
cc_791 N_S1_c_850_n N_A_509_392#_c_1555_n 0.00315355f $X=11.535 $Y=1.795 $X2=0
+ $Y2=0
cc_792 N_S1_c_864_n N_A_509_392#_c_1555_n 0.00309587f $X=11.535 $Y=1.885 $X2=0
+ $Y2=0
cc_793 N_S1_M1015_g N_A_509_392#_c_1555_n 0.00546568f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_794 N_S1_c_852_n N_A_509_392#_c_1555_n 0.00632518f $X=12.035 $Y=1.795 $X2=0
+ $Y2=0
cc_795 N_S1_c_866_n N_A_509_392#_c_1555_n 0.0105858f $X=12.035 $Y=1.885 $X2=0
+ $Y2=0
cc_796 N_S1_c_856_n N_A_509_392#_c_1555_n 0.0281339f $X=12.125 $Y=1.36 $X2=0
+ $Y2=0
cc_797 N_S1_c_861_n N_A_509_392#_c_1555_n 0.0403568f $X=12.665 $Y=1.455 $X2=0
+ $Y2=0
cc_798 N_S1_M1013_g N_A_1191_121#_c_1738_n 0.00687329f $X=11.355 $Y=0.69 $X2=0
+ $Y2=0
cc_799 N_S1_c_864_n N_A_1191_121#_c_1738_n 2.12928e-19 $X=11.535 $Y=1.885 $X2=0
+ $Y2=0
cc_800 N_S1_c_856_n N_A_1191_121#_c_1738_n 0.00197547f $X=12.125 $Y=1.36 $X2=0
+ $Y2=0
cc_801 N_S1_c_864_n N_A_1191_121#_c_1749_n 0.00434988f $X=11.535 $Y=1.885 $X2=0
+ $Y2=0
cc_802 N_S1_M1013_g N_A_1191_121#_c_1740_n 0.0115258f $X=11.355 $Y=0.69 $X2=0
+ $Y2=0
cc_803 N_S1_M1015_g N_A_1191_121#_c_1740_n 0.00147484f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_804 N_S1_c_864_n N_A_1191_121#_c_1750_n 0.0115217f $X=11.535 $Y=1.885 $X2=0
+ $Y2=0
cc_805 N_S1_c_866_n N_A_1191_121#_c_1750_n 0.00991323f $X=12.035 $Y=1.885 $X2=0
+ $Y2=0
cc_806 N_S1_c_864_n N_A_1191_121#_c_1753_n 2.15315e-19 $X=11.535 $Y=1.885 $X2=0
+ $Y2=0
cc_807 N_S1_c_854_n N_VGND_c_2082_n 0.00177323f $X=14.285 $Y=1.22 $X2=0 $Y2=0
cc_808 N_S1_M1013_g N_VGND_c_2090_n 0.00278271f $X=11.355 $Y=0.69 $X2=0 $Y2=0
cc_809 N_S1_M1015_g N_VGND_c_2090_n 0.00311652f $X=11.945 $Y=0.69 $X2=0 $Y2=0
cc_810 N_S1_c_854_n N_VGND_c_2090_n 0.00278271f $X=14.285 $Y=1.22 $X2=0 $Y2=0
cc_811 N_S1_M1013_g N_VGND_c_2100_n 0.00359811f $X=11.355 $Y=0.69 $X2=0 $Y2=0
cc_812 N_S1_M1015_g N_VGND_c_2100_n 0.00396569f $X=11.945 $Y=0.69 $X2=0 $Y2=0
cc_813 N_S1_c_854_n N_VGND_c_2100_n 0.00360685f $X=14.285 $Y=1.22 $X2=0 $Y2=0
cc_814 N_A_2489_347#_c_980_n N_A_2199_74#_c_1098_n 0.00182789f $X=12.535
+ $Y=1.885 $X2=0 $Y2=0
cc_815 N_A_2489_347#_c_980_n N_A_2199_74#_c_1085_n 0.00259032f $X=12.535
+ $Y=1.885 $X2=0 $Y2=0
cc_816 N_A_2489_347#_c_981_n N_A_2199_74#_c_1085_n 5.11707e-19 $X=13.035
+ $Y=1.885 $X2=0 $Y2=0
cc_817 N_A_2489_347#_c_978_n N_A_2199_74#_c_1085_n 3.41183e-19 $X=13.165
+ $Y=1.635 $X2=0 $Y2=0
cc_818 N_A_2489_347#_c_980_n N_A_2199_74#_c_1125_n 0.00611081f $X=12.535
+ $Y=1.885 $X2=0 $Y2=0
cc_819 N_A_2489_347#_c_981_n N_A_2199_74#_c_1125_n 2.69714e-19 $X=13.035
+ $Y=1.885 $X2=0 $Y2=0
cc_820 N_A_2489_347#_c_980_n N_A_2199_74#_c_1105_n 0.0107323f $X=12.535 $Y=1.885
+ $X2=0 $Y2=0
cc_821 N_A_2489_347#_c_981_n N_A_2199_74#_c_1105_n 0.0178859f $X=13.035 $Y=1.885
+ $X2=0 $Y2=0
cc_822 N_A_2489_347#_c_977_n N_A_2199_74#_c_1105_n 0.00913123f $X=13.165
+ $Y=1.635 $X2=0 $Y2=0
cc_823 N_A_2489_347#_c_978_n N_A_2199_74#_c_1105_n 0.00500631f $X=13.165
+ $Y=1.635 $X2=0 $Y2=0
cc_824 N_A_2489_347#_M1009_g N_A_2199_74#_c_1068_n 0.0116317f $X=12.795 $Y=0.69
+ $X2=0 $Y2=0
cc_825 N_A_2489_347#_M1048_g N_A_2199_74#_c_1068_n 0.0137009f $X=13.225 $Y=0.69
+ $X2=0 $Y2=0
cc_826 N_A_2489_347#_c_982_n N_A_2199_74#_c_1086_n 0.0120254f $X=13.875 $Y=1.805
+ $X2=0 $Y2=0
cc_827 N_A_2489_347#_c_983_n N_A_2199_74#_c_1086_n 0.00830695f $X=14.04 $Y=1.985
+ $X2=0 $Y2=0
cc_828 N_A_2489_347#_c_977_n N_A_2199_74#_c_1086_n 0.0153206f $X=13.165 $Y=1.635
+ $X2=0 $Y2=0
cc_829 N_A_2489_347#_c_978_n N_A_2199_74#_c_1086_n 0.0013544f $X=13.165 $Y=1.635
+ $X2=0 $Y2=0
cc_830 N_A_2489_347#_c_981_n N_A_2199_74#_c_1087_n 0.0147503f $X=13.035 $Y=1.885
+ $X2=0 $Y2=0
cc_831 N_A_2489_347#_c_983_n N_A_2199_74#_c_1087_n 0.0345589f $X=14.04 $Y=1.985
+ $X2=0 $Y2=0
cc_832 N_A_2489_347#_c_979_n N_A_2199_74#_c_1069_n 0.0244318f $X=14.07 $Y=0.775
+ $X2=0 $Y2=0
cc_833 N_A_2489_347#_M1010_s N_A_2199_74#_c_1070_n 0.00273752f $X=13.925 $Y=0.37
+ $X2=0 $Y2=0
cc_834 N_A_2489_347#_c_979_n N_A_2199_74#_c_1070_n 0.0184007f $X=14.07 $Y=0.775
+ $X2=0 $Y2=0
cc_835 N_A_2489_347#_c_976_n N_A_2199_74#_c_1071_n 0.0135902f $X=14.12 $Y=1.72
+ $X2=0 $Y2=0
cc_836 N_A_2489_347#_c_976_n N_A_2199_74#_c_1072_n 0.0255059f $X=14.12 $Y=1.72
+ $X2=0 $Y2=0
cc_837 N_A_2489_347#_M1009_g N_A_2199_74#_c_1075_n 0.00280783f $X=12.795 $Y=0.69
+ $X2=0 $Y2=0
cc_838 N_A_2489_347#_c_983_n N_VPWR_c_1277_n 0.044017f $X=14.04 $Y=1.985 $X2=0
+ $Y2=0
cc_839 N_A_2489_347#_c_987_n N_VPWR_c_1277_n 0.00376845f $X=14.04 $Y=1.805 $X2=0
+ $Y2=0
cc_840 N_A_2489_347#_c_980_n N_VPWR_c_1285_n 0.00278271f $X=12.535 $Y=1.885
+ $X2=0 $Y2=0
cc_841 N_A_2489_347#_c_981_n N_VPWR_c_1285_n 0.0044313f $X=13.035 $Y=1.885 $X2=0
+ $Y2=0
cc_842 N_A_2489_347#_c_983_n N_VPWR_c_1285_n 0.0146357f $X=14.04 $Y=1.985 $X2=0
+ $Y2=0
cc_843 N_A_2489_347#_c_980_n N_VPWR_c_1270_n 0.00354798f $X=12.535 $Y=1.885
+ $X2=0 $Y2=0
cc_844 N_A_2489_347#_c_981_n N_VPWR_c_1270_n 0.00859385f $X=13.035 $Y=1.885
+ $X2=0 $Y2=0
cc_845 N_A_2489_347#_c_983_n N_VPWR_c_1270_n 0.0121141f $X=14.04 $Y=1.985 $X2=0
+ $Y2=0
cc_846 N_A_2489_347#_M1009_g N_A_509_392#_c_1630_n 0.010582f $X=12.795 $Y=0.69
+ $X2=0 $Y2=0
cc_847 N_A_2489_347#_M1009_g N_A_509_392#_c_1554_n 0.00360839f $X=12.795 $Y=0.69
+ $X2=0 $Y2=0
cc_848 N_A_2489_347#_M1009_g N_A_509_392#_c_1635_n 0.00828563f $X=12.795 $Y=0.69
+ $X2=0 $Y2=0
cc_849 N_A_2489_347#_M1048_g N_A_509_392#_c_1635_n 0.00453241f $X=13.225 $Y=0.69
+ $X2=0 $Y2=0
cc_850 N_A_2489_347#_c_980_n N_A_509_392#_c_1555_n 4.42243e-19 $X=12.535
+ $Y=1.885 $X2=0 $Y2=0
cc_851 N_A_2489_347#_c_978_n N_A_509_392#_c_1555_n 6.11957e-19 $X=13.165
+ $Y=1.635 $X2=0 $Y2=0
cc_852 N_A_2489_347#_c_980_n N_A_1191_121#_c_1750_n 0.0119779f $X=12.535
+ $Y=1.885 $X2=0 $Y2=0
cc_853 N_A_2489_347#_c_981_n N_A_1191_121#_c_1750_n 0.00685456f $X=13.035
+ $Y=1.885 $X2=0 $Y2=0
cc_854 N_A_2489_347#_c_981_n N_A_1191_121#_c_1826_n 0.00520993f $X=13.035
+ $Y=1.885 $X2=0 $Y2=0
cc_855 N_A_2489_347#_c_987_n N_X_c_1998_n 6.16447e-19 $X=14.04 $Y=1.805 $X2=0
+ $Y2=0
cc_856 N_A_2489_347#_M1009_g N_VGND_c_2090_n 0.00278271f $X=12.795 $Y=0.69 $X2=0
+ $Y2=0
cc_857 N_A_2489_347#_M1048_g N_VGND_c_2090_n 0.00278271f $X=13.225 $Y=0.69 $X2=0
+ $Y2=0
cc_858 N_A_2489_347#_M1009_g N_VGND_c_2100_n 0.0035536f $X=12.795 $Y=0.69 $X2=0
+ $Y2=0
cc_859 N_A_2489_347#_M1048_g N_VGND_c_2100_n 0.00358427f $X=13.225 $Y=0.69 $X2=0
+ $Y2=0
cc_860 N_A_2199_74#_c_1079_n N_VPWR_c_1277_n 0.00967877f $X=14.815 $Y=1.765
+ $X2=0 $Y2=0
cc_861 N_A_2199_74#_c_1072_n N_VPWR_c_1277_n 0.0145645f $X=14.545 $Y=1.465 $X2=0
+ $Y2=0
cc_862 N_A_2199_74#_c_1073_n N_VPWR_c_1277_n 0.0129622f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_863 N_A_2199_74#_c_1080_n N_VPWR_c_1278_n 0.00646055f $X=15.265 $Y=1.765
+ $X2=0 $Y2=0
cc_864 N_A_2199_74#_c_1081_n N_VPWR_c_1278_n 0.00620497f $X=15.765 $Y=1.765
+ $X2=0 $Y2=0
cc_865 N_A_2199_74#_c_1082_n N_VPWR_c_1280_n 0.0198182f $X=16.215 $Y=1.765 $X2=0
+ $Y2=0
cc_866 N_A_2199_74#_c_1087_n N_VPWR_c_1285_n 0.0146357f $X=13.31 $Y=2.485 $X2=0
+ $Y2=0
cc_867 N_A_2199_74#_c_1079_n N_VPWR_c_1287_n 0.00445602f $X=14.815 $Y=1.765
+ $X2=0 $Y2=0
cc_868 N_A_2199_74#_c_1080_n N_VPWR_c_1287_n 0.00445602f $X=15.265 $Y=1.765
+ $X2=0 $Y2=0
cc_869 N_A_2199_74#_c_1081_n N_VPWR_c_1293_n 0.00445602f $X=15.765 $Y=1.765
+ $X2=0 $Y2=0
cc_870 N_A_2199_74#_c_1082_n N_VPWR_c_1293_n 0.00445602f $X=16.215 $Y=1.765
+ $X2=0 $Y2=0
cc_871 N_A_2199_74#_c_1079_n N_VPWR_c_1270_n 0.00857553f $X=14.815 $Y=1.765
+ $X2=0 $Y2=0
cc_872 N_A_2199_74#_c_1080_n N_VPWR_c_1270_n 0.0085805f $X=15.265 $Y=1.765 $X2=0
+ $Y2=0
cc_873 N_A_2199_74#_c_1081_n N_VPWR_c_1270_n 0.00857378f $X=15.765 $Y=1.765
+ $X2=0 $Y2=0
cc_874 N_A_2199_74#_c_1082_n N_VPWR_c_1270_n 0.00860648f $X=16.215 $Y=1.765
+ $X2=0 $Y2=0
cc_875 N_A_2199_74#_c_1087_n N_VPWR_c_1270_n 0.0121141f $X=13.31 $Y=2.485 $X2=0
+ $Y2=0
cc_876 N_A_2199_74#_c_1068_n N_A_509_392#_M1009_s 0.00176461f $X=13.345 $Y=0.34
+ $X2=0 $Y2=0
cc_877 N_A_2199_74#_c_1098_n N_A_509_392#_M1001_s 0.00481926f $X=12.145 $Y=2.65
+ $X2=0 $Y2=0
cc_878 N_A_2199_74#_M1015_s N_A_509_392#_c_1549_n 0.00394438f $X=12.02 $Y=0.37
+ $X2=0 $Y2=0
cc_879 N_A_2199_74#_c_1067_n N_A_509_392#_c_1549_n 0.00829606f $X=12.493
+ $Y=0.437 $X2=0 $Y2=0
cc_880 N_A_2199_74#_c_1116_n N_A_509_392#_c_1549_n 0.00937046f $X=11.985 $Y=0.51
+ $X2=0 $Y2=0
cc_881 N_A_2199_74#_c_1074_n N_A_509_392#_c_1550_n 0.0117142f $X=11.265 $Y=0.68
+ $X2=0 $Y2=0
cc_882 N_A_2199_74#_c_1116_n N_A_509_392#_c_1550_n 0.0216666f $X=11.985 $Y=0.51
+ $X2=0 $Y2=0
cc_883 N_A_2199_74#_M1015_s N_A_509_392#_c_1630_n 0.00500868f $X=12.02 $Y=0.37
+ $X2=0 $Y2=0
cc_884 N_A_2199_74#_c_1068_n N_A_509_392#_c_1630_n 0.00445011f $X=13.345 $Y=0.34
+ $X2=0 $Y2=0
cc_885 N_A_2199_74#_c_1076_n N_A_509_392#_c_1630_n 0.0125748f $X=12.675 $Y=0.437
+ $X2=0 $Y2=0
cc_886 N_A_2199_74#_M1015_s N_A_509_392#_c_1554_n 0.00692408f $X=12.02 $Y=0.37
+ $X2=0 $Y2=0
cc_887 N_A_2199_74#_c_1067_n N_A_509_392#_c_1554_n 0.0131573f $X=12.493 $Y=0.437
+ $X2=0 $Y2=0
cc_888 N_A_2199_74#_c_1068_n N_A_509_392#_c_1635_n 0.0142275f $X=13.345 $Y=0.34
+ $X2=0 $Y2=0
cc_889 N_A_2199_74#_c_1066_n N_A_509_392#_c_1563_n 0.0386176f $X=11.31 $Y=2.105
+ $X2=0 $Y2=0
cc_890 N_A_2199_74#_c_1098_n N_A_509_392#_c_1563_n 0.00383998f $X=12.145 $Y=2.65
+ $X2=0 $Y2=0
cc_891 N_A_2199_74#_c_1066_n N_A_509_392#_c_1566_n 0.00265576f $X=11.31 $Y=2.105
+ $X2=0 $Y2=0
cc_892 N_A_2199_74#_c_1098_n N_A_509_392#_c_1566_n 0.00226942f $X=12.145 $Y=2.65
+ $X2=0 $Y2=0
cc_893 N_A_2199_74#_c_1085_n N_A_509_392#_c_1566_n 0.00133571f $X=12.31 $Y=2.23
+ $X2=0 $Y2=0
cc_894 N_A_2199_74#_c_1066_n N_A_509_392#_c_1555_n 0.0846651f $X=11.31 $Y=2.105
+ $X2=0 $Y2=0
cc_895 N_A_2199_74#_c_1098_n N_A_509_392#_c_1555_n 0.019415f $X=12.145 $Y=2.65
+ $X2=0 $Y2=0
cc_896 N_A_2199_74#_c_1085_n N_A_509_392#_c_1555_n 0.0108722f $X=12.31 $Y=2.23
+ $X2=0 $Y2=0
cc_897 N_A_2199_74#_c_1116_n N_A_1191_121#_M1013_d 0.00871026f $X=11.985 $Y=0.51
+ $X2=0 $Y2=0
cc_898 N_A_2199_74#_c_1105_n N_A_1191_121#_M1011_d 0.0060005f $X=13.145 $Y=2.145
+ $X2=0 $Y2=0
cc_899 N_A_2199_74#_c_1066_n N_A_1191_121#_c_1738_n 0.0539165f $X=11.31 $Y=2.105
+ $X2=0 $Y2=0
cc_900 N_A_2199_74#_c_1074_n N_A_1191_121#_c_1738_n 0.0344938f $X=11.265 $Y=0.68
+ $X2=0 $Y2=0
cc_901 N_A_2199_74#_c_1066_n N_A_1191_121#_c_1749_n 0.0355988f $X=11.31 $Y=2.105
+ $X2=0 $Y2=0
cc_902 N_A_2199_74#_c_1084_n N_A_1191_121#_c_1749_n 0.0143582f $X=11.475 $Y=2.65
+ $X2=0 $Y2=0
cc_903 N_A_2199_74#_M1013_s N_A_1191_121#_c_1740_n 0.00441657f $X=10.995 $Y=0.37
+ $X2=0 $Y2=0
cc_904 N_A_2199_74#_c_1074_n N_A_1191_121#_c_1740_n 0.0231725f $X=11.265 $Y=0.68
+ $X2=0 $Y2=0
cc_905 N_A_2199_74#_c_1116_n N_A_1191_121#_c_1740_n 0.0222818f $X=11.985 $Y=0.51
+ $X2=0 $Y2=0
cc_906 N_A_2199_74#_c_1075_n N_A_1191_121#_c_1740_n 0.012401f $X=12.155 $Y=0.51
+ $X2=0 $Y2=0
cc_907 N_A_2199_74#_M1001_d N_A_1191_121#_c_1750_n 0.00287371f $X=11.165 $Y=1.96
+ $X2=0 $Y2=0
cc_908 N_A_2199_74#_M1044_d N_A_1191_121#_c_1750_n 0.00250873f $X=12.11 $Y=1.96
+ $X2=0 $Y2=0
cc_909 N_A_2199_74#_c_1098_n N_A_1191_121#_c_1750_n 0.0532727f $X=12.145 $Y=2.65
+ $X2=0 $Y2=0
cc_910 N_A_2199_74#_c_1084_n N_A_1191_121#_c_1750_n 0.0206482f $X=11.475 $Y=2.65
+ $X2=0 $Y2=0
cc_911 N_A_2199_74#_c_1105_n N_A_1191_121#_c_1750_n 0.00287635f $X=13.145
+ $Y=2.145 $X2=0 $Y2=0
cc_912 N_A_2199_74#_c_1087_n N_A_1191_121#_c_1750_n 0.00395311f $X=13.31
+ $Y=2.485 $X2=0 $Y2=0
cc_913 N_A_2199_74#_c_1105_n N_A_1191_121#_c_1826_n 0.0202127f $X=13.145
+ $Y=2.145 $X2=0 $Y2=0
cc_914 N_A_2199_74#_c_1066_n N_A_1191_121#_c_1753_n 0.0129149f $X=11.31 $Y=2.105
+ $X2=0 $Y2=0
cc_915 N_A_2199_74#_c_1079_n N_X_c_1996_n 0.0106573f $X=14.815 $Y=1.765 $X2=0
+ $Y2=0
cc_916 N_A_2199_74#_c_1080_n N_X_c_1996_n 0.0127555f $X=15.265 $Y=1.765 $X2=0
+ $Y2=0
cc_917 N_A_2199_74#_c_1081_n N_X_c_1996_n 7.39949e-19 $X=15.765 $Y=1.765 $X2=0
+ $Y2=0
cc_918 N_A_2199_74#_M1016_g N_X_c_1989_n 0.00760419f $X=15.015 $Y=0.74 $X2=0
+ $Y2=0
cc_919 N_A_2199_74#_M1026_g N_X_c_1989_n 3.97481e-19 $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_920 N_A_2199_74#_c_1080_n N_X_c_1997_n 0.0122806f $X=15.265 $Y=1.765 $X2=0
+ $Y2=0
cc_921 N_A_2199_74#_c_1081_n N_X_c_1997_n 0.0122806f $X=15.765 $Y=1.765 $X2=0
+ $Y2=0
cc_922 N_A_2199_74#_c_1073_n N_X_c_1997_n 0.0455181f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_923 N_A_2199_74#_c_1078_n N_X_c_1997_n 0.00906657f $X=16.215 $Y=1.532 $X2=0
+ $Y2=0
cc_924 N_A_2199_74#_c_1079_n N_X_c_1998_n 0.00254313f $X=14.815 $Y=1.765 $X2=0
+ $Y2=0
cc_925 N_A_2199_74#_c_1080_n N_X_c_1998_n 9.3899e-19 $X=15.265 $Y=1.765 $X2=0
+ $Y2=0
cc_926 N_A_2199_74#_c_1073_n N_X_c_1998_n 0.0276943f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_927 N_A_2199_74#_c_1078_n N_X_c_1998_n 0.00795526f $X=16.215 $Y=1.532 $X2=0
+ $Y2=0
cc_928 N_A_2199_74#_M1026_g N_X_c_1990_n 0.0124899f $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_929 N_A_2199_74#_M1029_g N_X_c_1990_n 0.01115f $X=15.875 $Y=0.74 $X2=0 $Y2=0
cc_930 N_A_2199_74#_c_1073_n N_X_c_1990_n 0.0447482f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_931 N_A_2199_74#_c_1078_n N_X_c_1990_n 0.00234554f $X=16.215 $Y=1.532 $X2=0
+ $Y2=0
cc_932 N_A_2199_74#_M1016_g N_X_c_1991_n 0.00245337f $X=15.015 $Y=0.74 $X2=0
+ $Y2=0
cc_933 N_A_2199_74#_c_1073_n N_X_c_1991_n 0.0209731f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_934 N_A_2199_74#_c_1078_n N_X_c_1991_n 0.00270102f $X=16.215 $Y=1.532 $X2=0
+ $Y2=0
cc_935 N_A_2199_74#_c_1080_n N_X_c_1999_n 6.39139e-19 $X=15.265 $Y=1.765 $X2=0
+ $Y2=0
cc_936 N_A_2199_74#_c_1081_n N_X_c_1999_n 0.0121613f $X=15.765 $Y=1.765 $X2=0
+ $Y2=0
cc_937 N_A_2199_74#_c_1082_n N_X_c_1999_n 0.0165744f $X=16.215 $Y=1.765 $X2=0
+ $Y2=0
cc_938 N_A_2199_74#_M1026_g N_X_c_1992_n 6.20738e-19 $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_939 N_A_2199_74#_M1029_g N_X_c_1992_n 0.00866629f $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_940 N_A_2199_74#_M1050_g N_X_c_1992_n 3.97481e-19 $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_941 N_A_2199_74#_c_1082_n N_X_c_2000_n 0.0146401f $X=16.215 $Y=1.765 $X2=0
+ $Y2=0
cc_942 N_A_2199_74#_c_1073_n N_X_c_2000_n 0.0038938f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_943 N_A_2199_74#_c_1078_n N_X_c_2000_n 0.00290392f $X=16.215 $Y=1.532 $X2=0
+ $Y2=0
cc_944 N_A_2199_74#_M1050_g N_X_c_1993_n 0.0158508f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_945 N_A_2199_74#_c_1073_n N_X_c_1993_n 0.0025934f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_946 N_A_2199_74#_c_1081_n N_X_c_2001_n 9.3899e-19 $X=15.765 $Y=1.765 $X2=0
+ $Y2=0
cc_947 N_A_2199_74#_c_1082_n N_X_c_2001_n 9.3899e-19 $X=16.215 $Y=1.765 $X2=0
+ $Y2=0
cc_948 N_A_2199_74#_c_1073_n N_X_c_2001_n 0.0276943f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_949 N_A_2199_74#_c_1078_n N_X_c_2001_n 0.00794155f $X=16.215 $Y=1.532 $X2=0
+ $Y2=0
cc_950 N_A_2199_74#_M1029_g N_X_c_1994_n 9.7541e-19 $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_951 N_A_2199_74#_c_1073_n N_X_c_1994_n 0.0209731f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_952 N_A_2199_74#_c_1078_n N_X_c_1994_n 0.00235428f $X=16.215 $Y=1.532 $X2=0
+ $Y2=0
cc_953 N_A_2199_74#_c_1082_n X 0.00122632f $X=16.215 $Y=1.765 $X2=0 $Y2=0
cc_954 N_A_2199_74#_M1050_g X 0.0169854f $X=16.305 $Y=0.74 $X2=0 $Y2=0
cc_955 N_A_2199_74#_c_1073_n X 0.0209823f $X=16.125 $Y=1.465 $X2=0 $Y2=0
cc_956 N_A_2199_74#_c_1078_n X 0.00504915f $X=16.215 $Y=1.532 $X2=0 $Y2=0
cc_957 N_A_2199_74#_c_1070_n N_VGND_M1010_d 5.37942e-19 $X=14.375 $Y=0.34 $X2=0
+ $Y2=0
cc_958 N_A_2199_74#_c_1071_n N_VGND_M1010_d 0.00934994f $X=14.46 $Y=1.3 $X2=0
+ $Y2=0
cc_959 N_A_2199_74#_M1016_g N_VGND_c_2082_n 0.00262092f $X=15.015 $Y=0.74 $X2=0
+ $Y2=0
cc_960 N_A_2199_74#_c_1070_n N_VGND_c_2082_n 0.014187f $X=14.375 $Y=0.34 $X2=0
+ $Y2=0
cc_961 N_A_2199_74#_c_1071_n N_VGND_c_2082_n 0.0512232f $X=14.46 $Y=1.3 $X2=0
+ $Y2=0
cc_962 N_A_2199_74#_c_1073_n N_VGND_c_2082_n 0.0148609f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_963 N_A_2199_74#_c_1078_n N_VGND_c_2082_n 8.1907e-19 $X=16.215 $Y=1.532 $X2=0
+ $Y2=0
cc_964 N_A_2199_74#_M1016_g N_VGND_c_2083_n 5.05592e-19 $X=15.015 $Y=0.74 $X2=0
+ $Y2=0
cc_965 N_A_2199_74#_M1026_g N_VGND_c_2083_n 0.00914496f $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_966 N_A_2199_74#_M1029_g N_VGND_c_2083_n 0.00183835f $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_967 N_A_2199_74#_M1029_g N_VGND_c_2085_n 5.04273e-19 $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_968 N_A_2199_74#_M1050_g N_VGND_c_2085_n 0.0112604f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_969 N_A_2199_74#_c_1070_n N_VGND_c_2090_n 0.0567846f $X=14.375 $Y=0.34 $X2=0
+ $Y2=0
cc_970 N_A_2199_74#_c_1116_n N_VGND_c_2090_n 0.00265664f $X=11.985 $Y=0.51 $X2=0
+ $Y2=0
cc_971 N_A_2199_74#_c_1075_n N_VGND_c_2090_n 0.089252f $X=12.155 $Y=0.51 $X2=0
+ $Y2=0
cc_972 N_A_2199_74#_c_1077_n N_VGND_c_2090_n 0.0237213f $X=13.51 $Y=0.34 $X2=0
+ $Y2=0
cc_973 N_A_2199_74#_M1016_g N_VGND_c_2094_n 0.00434272f $X=15.015 $Y=0.74 $X2=0
+ $Y2=0
cc_974 N_A_2199_74#_M1026_g N_VGND_c_2094_n 0.00383152f $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_975 N_A_2199_74#_M1029_g N_VGND_c_2095_n 0.00434272f $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_976 N_A_2199_74#_M1050_g N_VGND_c_2095_n 0.00383152f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_977 N_A_2199_74#_M1016_g N_VGND_c_2100_n 0.00822542f $X=15.015 $Y=0.74 $X2=0
+ $Y2=0
cc_978 N_A_2199_74#_M1026_g N_VGND_c_2100_n 0.0075754f $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_979 N_A_2199_74#_M1029_g N_VGND_c_2100_n 0.00820284f $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_980 N_A_2199_74#_M1050_g N_VGND_c_2100_n 0.0075754f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_981 N_A_2199_74#_c_1070_n N_VGND_c_2100_n 0.032237f $X=14.375 $Y=0.34 $X2=0
+ $Y2=0
cc_982 N_A_2199_74#_c_1116_n N_VGND_c_2100_n 0.00514655f $X=11.985 $Y=0.51 $X2=0
+ $Y2=0
cc_983 N_A_2199_74#_c_1075_n N_VGND_c_2100_n 0.0500945f $X=12.155 $Y=0.51 $X2=0
+ $Y2=0
cc_984 N_A_2199_74#_c_1077_n N_VGND_c_2100_n 0.0128418f $X=13.51 $Y=0.34 $X2=0
+ $Y2=0
cc_985 N_VPWR_c_1272_n N_A_116_392#_c_1453_n 0.013464f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_986 N_VPWR_c_1272_n N_A_116_392#_c_1454_n 0.0563195f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_987 N_VPWR_c_1273_n N_A_116_392#_c_1454_n 0.0449538f $X=1.18 $Y=2.475 $X2=0
+ $Y2=0
cc_988 N_VPWR_c_1289_n N_A_116_392#_c_1454_n 0.014552f $X=1.095 $Y=3.33 $X2=0
+ $Y2=0
cc_989 N_VPWR_c_1270_n N_A_116_392#_c_1454_n 0.0119791f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_990 N_VPWR_M1041_d N_A_116_392#_c_1455_n 0.00420698f $X=1.03 $Y=1.96 $X2=0
+ $Y2=0
cc_991 N_VPWR_M1008_s N_A_116_392#_c_1455_n 0.00554645f $X=1.98 $Y=1.96 $X2=0
+ $Y2=0
cc_992 N_VPWR_c_1273_n N_A_116_392#_c_1455_n 0.0154248f $X=1.18 $Y=2.475 $X2=0
+ $Y2=0
cc_993 N_VPWR_M1008_s N_A_296_392#_c_1515_n 0.00591595f $X=1.98 $Y=1.96 $X2=0
+ $Y2=0
cc_994 N_VPWR_c_1274_n N_A_296_392#_c_1515_n 0.0198092f $X=2.13 $Y=2.815 $X2=0
+ $Y2=0
cc_995 N_VPWR_c_1270_n N_A_296_392#_c_1515_n 0.0154502f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_996 N_VPWR_c_1273_n N_A_296_392#_c_1517_n 0.0187702f $X=1.18 $Y=2.475 $X2=0
+ $Y2=0
cc_997 N_VPWR_c_1274_n N_A_296_392#_c_1517_n 0.0221564f $X=2.13 $Y=2.815 $X2=0
+ $Y2=0
cc_998 N_VPWR_c_1290_n N_A_296_392#_c_1517_n 0.0145781f $X=2.045 $Y=3.33 $X2=0
+ $Y2=0
cc_999 N_VPWR_c_1270_n N_A_296_392#_c_1517_n 0.0120405f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1000 N_VPWR_c_1291_n N_A_509_392#_c_1557_n 0.0396956f $X=5.4 $Y=3.33 $X2=0
+ $Y2=0
cc_1001 N_VPWR_c_1270_n N_A_509_392#_c_1557_n 0.0223402f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1002 N_VPWR_c_1291_n N_A_509_392#_c_1559_n 0.0595512f $X=5.4 $Y=3.33 $X2=0
+ $Y2=0
cc_1003 N_VPWR_c_1270_n N_A_509_392#_c_1559_n 0.0329703f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1004 N_VPWR_c_1274_n N_A_509_392#_c_1561_n 0.0280959f $X=2.13 $Y=2.815 $X2=0
+ $Y2=0
cc_1005 N_VPWR_c_1291_n N_A_509_392#_c_1561_n 0.0230359f $X=5.4 $Y=3.33 $X2=0
+ $Y2=0
cc_1006 N_VPWR_c_1270_n N_A_509_392#_c_1561_n 0.0127743f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1007 N_VPWR_c_1291_n N_A_509_392#_c_1562_n 0.0236039f $X=5.4 $Y=3.33 $X2=0
+ $Y2=0
cc_1008 N_VPWR_c_1270_n N_A_509_392#_c_1562_n 0.012761f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1009 N_VPWR_c_1275_n N_A_509_392#_c_1563_n 0.0309855f $X=5.565 $Y=1.985 $X2=0
+ $Y2=0
cc_1010 N_VPWR_c_1276_n N_A_509_392#_c_1563_n 0.00142931f $X=10.55 $Y=2.45 $X2=0
+ $Y2=0
cc_1011 N_VPWR_c_1275_n N_A_1191_121#_c_1743_n 0.010962f $X=5.565 $Y=1.985 $X2=0
+ $Y2=0
cc_1012 N_VPWR_c_1275_n N_A_1191_121#_c_1744_n 0.0565308f $X=5.565 $Y=1.985
+ $X2=0 $Y2=0
cc_1013 N_VPWR_c_1292_n N_A_1191_121#_c_1744_n 0.00849124f $X=8.32 $Y=3.33 $X2=0
+ $Y2=0
cc_1014 N_VPWR_c_1270_n N_A_1191_121#_c_1744_n 0.00873398f $X=16.56 $Y=3.33
+ $X2=0 $Y2=0
cc_1015 N_VPWR_M1007_s N_A_1191_121#_c_1747_n 0.00514671f $X=8.34 $Y=1.96 $X2=0
+ $Y2=0
cc_1016 N_VPWR_M1017_s N_A_1191_121#_c_1747_n 0.00770399f $X=9.32 $Y=1.96 $X2=0
+ $Y2=0
cc_1017 N_VPWR_M1046_d N_A_1191_121#_c_1747_n 0.00543701f $X=10.4 $Y=1.96 $X2=0
+ $Y2=0
cc_1018 N_VPWR_c_1276_n N_A_1191_121#_c_1747_n 0.0122803f $X=10.55 $Y=2.45 $X2=0
+ $Y2=0
cc_1019 N_VPWR_c_1276_n N_A_1191_121#_c_1749_n 0.0458208f $X=10.55 $Y=2.45 $X2=0
+ $Y2=0
cc_1020 N_VPWR_c_1285_n N_A_1191_121#_c_1750_n 0.129801f $X=14.375 $Y=3.33 $X2=0
+ $Y2=0
cc_1021 N_VPWR_c_1270_n N_A_1191_121#_c_1750_n 0.0734911f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1022 N_VPWR_c_1276_n N_A_1191_121#_c_1751_n 0.0142847f $X=10.55 $Y=2.45 $X2=0
+ $Y2=0
cc_1023 N_VPWR_c_1285_n N_A_1191_121#_c_1751_n 0.0121867f $X=14.375 $Y=3.33
+ $X2=0 $Y2=0
cc_1024 N_VPWR_c_1270_n N_A_1191_121#_c_1751_n 0.00660921f $X=16.56 $Y=3.33
+ $X2=0 $Y2=0
cc_1025 N_VPWR_c_1292_n N_A_1285_377#_c_1911_n 0.0798496f $X=8.32 $Y=3.33 $X2=0
+ $Y2=0
cc_1026 N_VPWR_c_1270_n N_A_1285_377#_c_1911_n 0.0466173f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1027 N_VPWR_c_1292_n N_A_1285_377#_c_1912_n 0.0236566f $X=8.32 $Y=3.33 $X2=0
+ $Y2=0
cc_1028 N_VPWR_c_1270_n N_A_1285_377#_c_1912_n 0.0128296f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1029 N_VPWR_M1007_s N_A_1285_377#_c_1913_n 0.00851715f $X=8.34 $Y=1.96 $X2=0
+ $Y2=0
cc_1030 N_VPWR_M1017_s N_A_1285_377#_c_1913_n 0.0112556f $X=9.32 $Y=1.96 $X2=0
+ $Y2=0
cc_1031 N_VPWR_c_1276_n N_A_1285_377#_c_1913_n 0.0239056f $X=10.55 $Y=2.45 $X2=0
+ $Y2=0
cc_1032 N_VPWR_c_1281_n N_A_1285_377#_c_1913_n 0.025977f $X=9.56 $Y=3.05 $X2=0
+ $Y2=0
cc_1033 N_VPWR_c_1282_n N_A_1285_377#_c_1913_n 0.0138793f $X=9.39 $Y=3.33 $X2=0
+ $Y2=0
cc_1034 N_VPWR_c_1283_n N_A_1285_377#_c_1913_n 0.0184897f $X=10.465 $Y=3.33
+ $X2=0 $Y2=0
cc_1035 N_VPWR_c_1292_n N_A_1285_377#_c_1913_n 0.00389376f $X=8.32 $Y=3.33 $X2=0
+ $Y2=0
cc_1036 N_VPWR_c_1297_n N_A_1285_377#_c_1913_n 0.0242244f $X=8.485 $Y=3.05 $X2=0
+ $Y2=0
cc_1037 N_VPWR_c_1270_n N_A_1285_377#_c_1913_n 0.0481175f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1038 N_VPWR_c_1276_n N_A_1285_377#_c_1926_n 0.0221136f $X=10.55 $Y=2.45 $X2=0
+ $Y2=0
cc_1039 N_VPWR_c_1292_n N_A_1285_377#_c_1914_n 0.0116773f $X=8.32 $Y=3.33 $X2=0
+ $Y2=0
cc_1040 N_VPWR_c_1297_n N_A_1285_377#_c_1914_n 0.00872136f $X=8.485 $Y=3.05
+ $X2=0 $Y2=0
cc_1041 N_VPWR_c_1270_n N_A_1285_377#_c_1914_n 0.00646299f $X=16.56 $Y=3.33
+ $X2=0 $Y2=0
cc_1042 N_VPWR_M1007_s N_A_1465_377#_c_1968_n 0.00843523f $X=8.34 $Y=1.96 $X2=0
+ $Y2=0
cc_1043 N_VPWR_c_1277_n N_X_c_1996_n 0.0386506f $X=14.54 $Y=1.985 $X2=0 $Y2=0
cc_1044 N_VPWR_c_1278_n N_X_c_1996_n 0.0563525f $X=15.49 $Y=2.305 $X2=0 $Y2=0
cc_1045 N_VPWR_c_1287_n N_X_c_1996_n 0.014552f $X=15.405 $Y=3.33 $X2=0 $Y2=0
cc_1046 N_VPWR_c_1270_n N_X_c_1996_n 0.0119791f $X=16.56 $Y=3.33 $X2=0 $Y2=0
cc_1047 N_VPWR_M1032_d N_X_c_1997_n 0.00275645f $X=15.34 $Y=1.84 $X2=0 $Y2=0
cc_1048 N_VPWR_c_1278_n N_X_c_1997_n 0.0184684f $X=15.49 $Y=2.305 $X2=0 $Y2=0
cc_1049 N_VPWR_c_1277_n N_X_c_1998_n 0.00711242f $X=14.54 $Y=1.985 $X2=0 $Y2=0
cc_1050 N_VPWR_c_1278_n N_X_c_1999_n 0.0322767f $X=15.49 $Y=2.305 $X2=0 $Y2=0
cc_1051 N_VPWR_c_1280_n N_X_c_1999_n 0.0323093f $X=16.49 $Y=2.305 $X2=0 $Y2=0
cc_1052 N_VPWR_c_1293_n N_X_c_1999_n 0.014552f $X=16.325 $Y=3.33 $X2=0 $Y2=0
cc_1053 N_VPWR_c_1270_n N_X_c_1999_n 0.0119791f $X=16.56 $Y=3.33 $X2=0 $Y2=0
cc_1054 N_VPWR_M1049_d N_X_c_2000_n 0.00432098f $X=16.29 $Y=1.84 $X2=0 $Y2=0
cc_1055 N_VPWR_c_1280_n N_X_c_2000_n 0.0268477f $X=16.49 $Y=2.305 $X2=0 $Y2=0
cc_1056 N_VPWR_c_1272_n N_VGND_c_2073_n 3.21545e-19 $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_1057 N_A_116_392#_c_1455_n N_A_296_392#_M1000_d 0.00448384f $X=2.525 $Y=2.055
+ $X2=-0.19 $Y2=-0.245
cc_1058 N_A_116_392#_c_1455_n N_A_296_392#_c_1515_n 0.0587823f $X=2.525 $Y=2.055
+ $X2=0 $Y2=0
cc_1059 N_A_116_392#_c_1451_n N_A_296_392#_c_1515_n 0.00774988f $X=4.02 $Y=1.685
+ $X2=0 $Y2=0
cc_1060 N_A_116_392#_c_1455_n N_A_296_392#_c_1516_n 0.00915303f $X=2.525
+ $Y=2.055 $X2=0 $Y2=0
cc_1061 N_A_116_392#_c_1456_n N_A_296_392#_c_1516_n 0.00144825f $X=2.61 $Y=1.97
+ $X2=0 $Y2=0
cc_1062 N_A_116_392#_c_1451_n N_A_296_392#_c_1516_n 0.025757f $X=4.02 $Y=1.685
+ $X2=0 $Y2=0
cc_1063 N_A_116_392#_c_1455_n N_A_296_392#_c_1517_n 0.0202766f $X=2.525 $Y=2.055
+ $X2=0 $Y2=0
cc_1064 N_A_116_392#_c_1455_n N_A_509_392#_M1003_s 0.00489304f $X=2.525 $Y=2.055
+ $X2=0 $Y2=0
cc_1065 N_A_116_392#_c_1451_n N_A_509_392#_c_1558_n 0.0275151f $X=4.02 $Y=1.685
+ $X2=0 $Y2=0
cc_1066 N_A_116_392#_c_1459_n N_A_509_392#_c_1558_n 0.0512738f $X=4.105 $Y=2.105
+ $X2=0 $Y2=0
cc_1067 N_A_116_392#_M1023_d N_A_509_392#_c_1559_n 0.00247267f $X=3.955 $Y=1.96
+ $X2=0 $Y2=0
cc_1068 N_A_116_392#_c_1459_n N_A_509_392#_c_1559_n 0.012787f $X=4.105 $Y=2.105
+ $X2=0 $Y2=0
cc_1069 N_A_116_392#_c_1459_n N_A_509_392#_c_1564_n 0.00151178f $X=4.105
+ $Y=2.105 $X2=0 $Y2=0
cc_1070 N_A_116_392#_c_1451_n N_A_509_392#_c_1556_n 0.0125064f $X=4.02 $Y=1.685
+ $X2=0 $Y2=0
cc_1071 N_A_116_392#_c_1459_n N_A_509_392#_c_1556_n 0.0653842f $X=4.105 $Y=2.105
+ $X2=0 $Y2=0
cc_1072 N_A_116_392#_c_1455_n N_A_299_126#_c_2324_n 0.00489672f $X=2.525
+ $Y=2.055 $X2=0 $Y2=0
cc_1073 N_A_116_392#_c_1451_n N_A_299_126#_c_2325_n 0.109901f $X=4.02 $Y=1.685
+ $X2=0 $Y2=0
cc_1074 N_A_116_392#_c_1452_n N_A_299_126#_c_2328_n 0.0145619f $X=2.695 $Y=1.685
+ $X2=0 $Y2=0
cc_1075 N_A_296_392#_c_1515_n N_A_509_392#_M1003_s 0.00738618f $X=2.99 $Y=2.395
+ $X2=0 $Y2=0
cc_1076 N_A_296_392#_M1003_d N_A_509_392#_c_1557_n 0.00224297f $X=3.005 $Y=1.96
+ $X2=0 $Y2=0
cc_1077 N_A_296_392#_c_1515_n N_A_509_392#_c_1557_n 0.00357384f $X=2.99 $Y=2.395
+ $X2=0 $Y2=0
cc_1078 N_A_296_392#_c_1524_n N_A_509_392#_c_1557_n 0.0164946f $X=3.145 $Y=2.395
+ $X2=0 $Y2=0
cc_1079 N_A_296_392#_c_1516_n N_A_509_392#_c_1558_n 0.00145482f $X=3.155
+ $Y=2.105 $X2=0 $Y2=0
cc_1080 N_A_296_392#_c_1515_n N_A_509_392#_c_1561_n 0.021143f $X=2.99 $Y=2.395
+ $X2=0 $Y2=0
cc_1081 N_A_509_392#_c_1550_n N_A_1191_121#_M1013_d 0.00270563f $X=11.975
+ $Y=1.02 $X2=0 $Y2=0
cc_1082 N_A_509_392#_c_1563_n N_A_1191_121#_M1019_s 0.00247227f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1083 N_A_509_392#_c_1563_n N_A_1191_121#_M1031_s 0.00243424f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1084 N_A_509_392#_c_1563_n N_A_1191_121#_c_1743_n 0.00759437f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1085 N_A_509_392#_c_1563_n N_A_1191_121#_c_1744_n 0.0182188f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1086 N_A_509_392#_c_1563_n N_A_1191_121#_c_1745_n 0.0291509f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1087 N_A_509_392#_c_1563_n N_A_1191_121#_c_1747_n 0.180826f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1088 N_A_509_392#_M1001_s N_A_1191_121#_c_1750_n 0.00251484f $X=11.61 $Y=1.96
+ $X2=0 $Y2=0
cc_1089 N_A_509_392#_c_1563_n N_A_1191_121#_c_1752_n 0.0242787f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1090 N_A_509_392#_c_1563_n N_A_1191_121#_c_1753_n 0.0312882f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1091 N_A_509_392#_c_1563_n N_A_1285_377#_M1019_d 0.00222287f $X=11.615
+ $Y=2.035 $X2=-0.19 $Y2=-0.245
cc_1092 N_A_509_392#_c_1563_n N_A_1285_377#_c_1915_n 0.00916663f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1093 N_A_509_392#_c_1563_n N_A_1285_377#_c_1913_n 0.00621187f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1094 N_A_509_392#_c_1563_n N_A_1285_377#_c_1926_n 0.00276748f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1095 N_A_509_392#_c_1563_n N_A_1465_377#_c_1968_n 0.0116025f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1096 N_A_509_392#_c_1563_n N_A_1465_377#_c_1970_n 0.00268168f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1097 N_A_509_392#_c_1551_n N_VGND_c_2077_n 0.0131469f $X=2.705 $Y=0.34 $X2=0
+ $Y2=0
cc_1098 N_A_509_392#_c_1547_n N_VGND_c_2078_n 0.00284916f $X=4.375 $Y=0.34 $X2=0
+ $Y2=0
cc_1099 N_A_509_392#_c_1545_n N_VGND_c_2093_n 0.0464419f $X=3.605 $Y=0.34 $X2=0
+ $Y2=0
cc_1100 N_A_509_392#_c_1547_n N_VGND_c_2093_n 0.0617583f $X=4.375 $Y=0.34 $X2=0
+ $Y2=0
cc_1101 N_A_509_392#_c_1551_n N_VGND_c_2093_n 0.0224527f $X=2.705 $Y=0.34 $X2=0
+ $Y2=0
cc_1102 N_A_509_392#_c_1552_n N_VGND_c_2093_n 0.0115893f $X=3.69 $Y=0.34 $X2=0
+ $Y2=0
cc_1103 N_A_509_392#_c_1545_n N_VGND_c_2100_n 0.0246622f $X=3.605 $Y=0.34 $X2=0
+ $Y2=0
cc_1104 N_A_509_392#_c_1547_n N_VGND_c_2100_n 0.0318225f $X=4.375 $Y=0.34 $X2=0
+ $Y2=0
cc_1105 N_A_509_392#_c_1551_n N_VGND_c_2100_n 0.0125544f $X=2.705 $Y=0.34 $X2=0
+ $Y2=0
cc_1106 N_A_509_392#_c_1552_n N_VGND_c_2100_n 0.00583135f $X=3.69 $Y=0.34 $X2=0
+ $Y2=0
cc_1107 N_A_509_392#_c_1545_n N_A_114_126#_c_2289_n 0.0211399f $X=3.605 $Y=0.34
+ $X2=0 $Y2=0
cc_1108 N_A_509_392#_M1004_d N_A_114_126#_c_2279_n 0.00868512f $X=2.56 $Y=0.31
+ $X2=0 $Y2=0
cc_1109 N_A_509_392#_c_1545_n N_A_114_126#_c_2279_n 0.00360515f $X=3.605 $Y=0.34
+ $X2=0 $Y2=0
cc_1110 N_A_509_392#_c_1551_n N_A_114_126#_c_2279_n 0.0246598f $X=2.705 $Y=0.34
+ $X2=0 $Y2=0
cc_1111 N_A_509_392#_c_1546_n N_A_299_126#_c_2325_n 0.0138021f $X=3.69 $Y=0.87
+ $X2=0 $Y2=0
cc_1112 N_A_509_392#_c_1556_n N_A_299_126#_c_2325_n 0.0136127f $X=4.547 $Y=1.92
+ $X2=0 $Y2=0
cc_1113 N_A_509_392#_c_1547_n N_A_299_126#_c_2326_n 0.0168109f $X=4.375 $Y=0.34
+ $X2=0 $Y2=0
cc_1114 N_A_509_392#_c_1548_n N_A_299_126#_c_2326_n 0.026002f $X=4.55 $Y=0.755
+ $X2=0 $Y2=0
cc_1115 N_A_509_392#_M1004_d N_A_299_126#_c_2328_n 0.00330374f $X=2.56 $Y=0.31
+ $X2=0 $Y2=0
cc_1116 N_A_1191_121#_c_1745_n N_A_1285_377#_M1019_d 8.76559e-19 $X=6.94 $Y=1.95
+ $X2=-0.19 $Y2=-0.245
cc_1117 N_A_1191_121#_c_1747_n N_A_1285_377#_M1033_s 0.00197722f $X=10.715
+ $Y=2.03 $X2=0 $Y2=0
cc_1118 N_A_1191_121#_c_1744_n N_A_1285_377#_c_1915_n 0.0469324f $X=6.125
+ $Y=2.74 $X2=0 $Y2=0
cc_1119 N_A_1191_121#_c_1745_n N_A_1285_377#_c_1915_n 0.0168414f $X=6.94 $Y=1.95
+ $X2=0 $Y2=0
cc_1120 N_A_1191_121#_c_1773_n N_A_1285_377#_c_1915_n 0.0347403f $X=7.025
+ $Y=2.57 $X2=0 $Y2=0
cc_1121 N_A_1191_121#_c_1773_n N_A_1285_377#_c_1911_n 0.0139345f $X=7.025
+ $Y=2.57 $X2=0 $Y2=0
cc_1122 N_A_1191_121#_c_1747_n N_A_1285_377#_c_1913_n 0.0153739f $X=10.715
+ $Y=2.03 $X2=0 $Y2=0
cc_1123 N_A_1191_121#_c_1747_n N_A_1285_377#_c_1926_n 0.0154682f $X=10.715
+ $Y=2.03 $X2=0 $Y2=0
cc_1124 N_A_1191_121#_M1045_d N_A_1285_377#_c_1914_n 0.00525997f $X=7.775
+ $Y=1.885 $X2=0 $Y2=0
cc_1125 N_A_1191_121#_c_1747_n N_A_1465_377#_M1005_s 0.0035622f $X=10.715
+ $Y=2.03 $X2=-0.19 $Y2=-0.245
cc_1126 N_A_1191_121#_c_1747_n N_A_1465_377#_M1007_d 0.00198204f $X=10.715
+ $Y=2.03 $X2=0 $Y2=0
cc_1127 N_A_1191_121#_M1045_d N_A_1465_377#_c_1968_n 0.00663155f $X=7.775
+ $Y=1.885 $X2=0 $Y2=0
cc_1128 N_A_1191_121#_c_1747_n N_A_1465_377#_c_1968_n 0.0860288f $X=10.715
+ $Y=2.03 $X2=0 $Y2=0
cc_1129 N_A_1191_121#_c_1747_n N_A_1465_377#_c_1970_n 0.0150487f $X=10.715
+ $Y=2.03 $X2=0 $Y2=0
cc_1130 N_A_1191_121#_c_1733_n N_VGND_c_2078_n 0.0075116f $X=6.06 $Y=1.025 $X2=0
+ $Y2=0
cc_1131 N_A_1191_121#_c_1734_n N_VGND_c_2078_n 0.0290212f $X=6.1 $Y=0.75 $X2=0
+ $Y2=0
cc_1132 N_A_1191_121#_c_1738_n N_VGND_c_2081_n 0.0460466f $X=10.8 $Y=1.945 $X2=0
+ $Y2=0
cc_1133 N_A_1191_121#_c_1739_n N_VGND_c_2081_n 0.0146661f $X=10.885 $Y=0.34
+ $X2=0 $Y2=0
cc_1134 N_A_1191_121#_c_1734_n N_VGND_c_2087_n 0.00553716f $X=6.1 $Y=0.75 $X2=0
+ $Y2=0
cc_1135 N_A_1191_121#_c_1739_n N_VGND_c_2090_n 0.0121867f $X=10.885 $Y=0.34
+ $X2=0 $Y2=0
cc_1136 N_A_1191_121#_c_1740_n N_VGND_c_2090_n 0.0591438f $X=11.65 $Y=0.34 $X2=0
+ $Y2=0
cc_1137 N_A_1191_121#_M1013_d N_VGND_c_2100_n 0.00246676f $X=11.43 $Y=0.37 $X2=0
+ $Y2=0
cc_1138 N_A_1191_121#_c_1734_n N_VGND_c_2100_n 0.00678664f $X=6.1 $Y=0.75 $X2=0
+ $Y2=0
cc_1139 N_A_1191_121#_c_1739_n N_VGND_c_2100_n 0.00660921f $X=10.885 $Y=0.34
+ $X2=0 $Y2=0
cc_1140 N_A_1191_121#_c_1740_n N_VGND_c_2100_n 0.0342794f $X=11.65 $Y=0.34 $X2=0
+ $Y2=0
cc_1141 N_A_1191_121#_c_1761_n N_A_1278_121#_M1002_s 0.00330483f $X=6.875
+ $Y=1.11 $X2=-0.19 $Y2=-0.245
cc_1142 N_A_1191_121#_c_1734_n N_A_1278_121#_c_2366_n 0.0104051f $X=6.1 $Y=0.75
+ $X2=0 $Y2=0
cc_1143 N_A_1191_121#_c_1761_n N_A_1278_121#_c_2366_n 0.0169041f $X=6.875
+ $Y=1.11 $X2=0 $Y2=0
cc_1144 N_A_1191_121#_c_1735_n N_A_1278_121#_c_2366_n 0.00652315f $X=7 $Y=0.765
+ $X2=0 $Y2=0
cc_1145 N_A_1191_121#_c_1761_n N_A_1278_121#_c_2367_n 0.00425327f $X=6.875
+ $Y=1.11 $X2=0 $Y2=0
cc_1146 N_A_1191_121#_c_1735_n N_A_1278_121#_c_2367_n 0.0196444f $X=7 $Y=0.765
+ $X2=0 $Y2=0
cc_1147 N_A_1191_121#_c_1737_n N_A_1278_121#_c_2367_n 0.0422737f $X=7.735
+ $Y=0.68 $X2=0 $Y2=0
cc_1148 N_A_1191_121#_c_1742_n N_A_1278_121#_c_2367_n 0.0185406f $X=7.86 $Y=0.68
+ $X2=0 $Y2=0
cc_1149 N_A_1191_121#_c_1742_n N_A_1278_121#_c_2371_n 0.0125333f $X=7.86 $Y=0.68
+ $X2=0 $Y2=0
cc_1150 N_A_1191_121#_c_1737_n N_A_1450_121#_M1006_d 0.00168086f $X=7.735
+ $Y=0.68 $X2=-0.19 $Y2=-0.245
cc_1151 N_A_1191_121#_M1040_s N_A_1450_121#_c_2419_n 0.00486971f $X=7.68
+ $Y=0.605 $X2=0 $Y2=0
cc_1152 N_A_1191_121#_c_1737_n N_A_1450_121#_c_2419_n 0.00498063f $X=7.735
+ $Y=0.68 $X2=0 $Y2=0
cc_1153 N_A_1191_121#_c_1742_n N_A_1450_121#_c_2419_n 0.0189683f $X=7.86 $Y=0.68
+ $X2=0 $Y2=0
cc_1154 N_A_1191_121#_c_1738_n N_A_1450_121#_c_2420_n 0.00207966f $X=10.8
+ $Y=1.945 $X2=0 $Y2=0
cc_1155 N_A_1191_121#_c_1737_n N_A_1450_121#_c_2422_n 0.0144331f $X=7.735
+ $Y=0.68 $X2=0 $Y2=0
cc_1156 N_A_1191_121#_c_1741_n N_A_1450_121#_c_2422_n 0.00998734f $X=7 $Y=1.145
+ $X2=0 $Y2=0
cc_1157 N_A_1191_121#_c_1742_n N_A_1450_121#_c_2423_n 3.61824e-19 $X=7.86
+ $Y=0.68 $X2=0 $Y2=0
cc_1158 N_A_1285_377#_c_1913_n N_A_1465_377#_M1007_d 0.0047939f $X=9.935 $Y=2.71
+ $X2=0 $Y2=0
cc_1159 N_A_1285_377#_c_1911_n N_A_1465_377#_c_1968_n 0.0107181f $X=7.98 $Y=2.99
+ $X2=0 $Y2=0
cc_1160 N_A_1285_377#_c_1913_n N_A_1465_377#_c_1968_n 0.0603383f $X=9.935
+ $Y=2.71 $X2=0 $Y2=0
cc_1161 N_A_1285_377#_c_1914_n N_A_1465_377#_c_1968_n 0.0129848f $X=8.065
+ $Y=2.71 $X2=0 $Y2=0
cc_1162 N_A_1285_377#_c_1911_n N_A_1465_377#_c_1970_n 0.0201386f $X=7.98 $Y=2.99
+ $X2=0 $Y2=0
cc_1163 N_A_1285_377#_c_1914_n N_A_1465_377#_c_1970_n 0.00476699f $X=8.065
+ $Y=2.71 $X2=0 $Y2=0
cc_1164 N_X_c_1990_n N_VGND_M1026_s 0.00176461f $X=15.925 $Y=1.045 $X2=0 $Y2=0
cc_1165 N_X_c_1993_n N_VGND_M1050_s 0.00338075f $X=16.445 $Y=1.045 $X2=0 $Y2=0
cc_1166 N_X_c_1989_n N_VGND_c_2082_n 0.0216048f $X=15.23 $Y=0.515 $X2=0 $Y2=0
cc_1167 N_X_c_1991_n N_VGND_c_2082_n 0.00752767f $X=15.315 $Y=1.045 $X2=0 $Y2=0
cc_1168 N_X_c_1989_n N_VGND_c_2083_n 0.0158413f $X=15.23 $Y=0.515 $X2=0 $Y2=0
cc_1169 N_X_c_1990_n N_VGND_c_2083_n 0.0152916f $X=15.925 $Y=1.045 $X2=0 $Y2=0
cc_1170 N_X_c_1992_n N_VGND_c_2083_n 0.0158413f $X=16.09 $Y=0.515 $X2=0 $Y2=0
cc_1171 N_X_c_1992_n N_VGND_c_2085_n 0.0164981f $X=16.09 $Y=0.515 $X2=0 $Y2=0
cc_1172 N_X_c_1993_n N_VGND_c_2085_n 0.023173f $X=16.445 $Y=1.045 $X2=0 $Y2=0
cc_1173 N_X_c_1989_n N_VGND_c_2094_n 0.0109942f $X=15.23 $Y=0.515 $X2=0 $Y2=0
cc_1174 N_X_c_1992_n N_VGND_c_2095_n 0.0109942f $X=16.09 $Y=0.515 $X2=0 $Y2=0
cc_1175 N_X_c_1989_n N_VGND_c_2100_n 0.00904371f $X=15.23 $Y=0.515 $X2=0 $Y2=0
cc_1176 N_X_c_1992_n N_VGND_c_2100_n 0.00904371f $X=16.09 $Y=0.515 $X2=0 $Y2=0
cc_1177 N_VGND_c_2075_n N_A_114_126#_M1025_s 0.00178571f $X=1.045 $Y=1.155
+ $X2=-0.19 $Y2=-0.245
cc_1178 N_VGND_c_2074_n N_A_114_126#_c_2274_n 0.0201555f $X=0.28 $Y=0.775 $X2=0
+ $Y2=0
cc_1179 N_VGND_c_2075_n N_A_114_126#_c_2274_n 0.0173292f $X=1.045 $Y=1.155 $X2=0
+ $Y2=0
cc_1180 N_VGND_c_2075_n N_A_114_126#_c_2275_n 0.00448545f $X=1.045 $Y=1.155
+ $X2=0 $Y2=0
cc_1181 N_VGND_c_2114_n N_A_114_126#_c_2275_n 0.022569f $X=1.17 $Y=0.805 $X2=0
+ $Y2=0
cc_1182 N_VGND_c_2077_n N_A_114_126#_c_2275_n 0.0154808f $X=2.145 $Y=0.365 $X2=0
+ $Y2=0
cc_1183 N_VGND_c_2092_n N_A_114_126#_c_2275_n 0.0550594f $X=1.98 $Y=0 $X2=0
+ $Y2=0
cc_1184 N_VGND_c_2100_n N_A_114_126#_c_2275_n 0.0350536f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1185 N_VGND_c_2074_n N_A_114_126#_c_2276_n 0.0162425f $X=0.28 $Y=0.775 $X2=0
+ $Y2=0
cc_1186 N_VGND_c_2092_n N_A_114_126#_c_2276_n 0.0207641f $X=1.98 $Y=0 $X2=0
+ $Y2=0
cc_1187 N_VGND_c_2100_n N_A_114_126#_c_2276_n 0.0126529f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1188 N_VGND_M1022_s N_A_114_126#_c_2278_n 0.0111424f $X=1.925 $Y=0.63 $X2=0
+ $Y2=0
cc_1189 N_VGND_c_2114_n N_A_114_126#_c_2278_n 0.0105495f $X=1.17 $Y=0.805 $X2=0
+ $Y2=0
cc_1190 N_VGND_c_2077_n N_A_114_126#_c_2278_n 0.0127545f $X=2.145 $Y=0.365 $X2=0
+ $Y2=0
cc_1191 N_VGND_c_2092_n N_A_114_126#_c_2278_n 0.00298933f $X=1.98 $Y=0 $X2=0
+ $Y2=0
cc_1192 N_VGND_c_2100_n N_A_114_126#_c_2278_n 0.00562944f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1193 N_VGND_M1022_s N_A_114_126#_c_2279_n 0.00425076f $X=1.925 $Y=0.63 $X2=0
+ $Y2=0
cc_1194 N_VGND_c_2077_n N_A_114_126#_c_2279_n 0.00511893f $X=2.145 $Y=0.365
+ $X2=0 $Y2=0
cc_1195 N_VGND_c_2100_n N_A_114_126#_c_2279_n 0.00983818f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1196 N_VGND_M1022_s N_A_299_126#_c_2324_n 0.00470132f $X=1.925 $Y=0.63 $X2=0
+ $Y2=0
cc_1197 N_VGND_c_2076_n N_A_299_126#_c_2327_n 0.0104027f $X=1.207 $Y=1.03 $X2=0
+ $Y2=0
cc_1198 N_VGND_c_2078_n N_A_1278_121#_c_2366_n 0.00470266f $X=5.54 $Y=0.515
+ $X2=0 $Y2=0
cc_1199 N_VGND_c_2086_n N_A_1278_121#_c_2367_n 0.0137091f $X=8.66 $Y=0 $X2=0
+ $Y2=0
cc_1200 N_VGND_c_2087_n N_A_1278_121#_c_2367_n 0.105357f $X=8.495 $Y=0 $X2=0
+ $Y2=0
cc_1201 N_VGND_c_2100_n N_A_1278_121#_c_2367_n 0.054907f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1202 N_VGND_c_2078_n N_A_1278_121#_c_2368_n 0.00581676f $X=5.54 $Y=0.515
+ $X2=0 $Y2=0
cc_1203 N_VGND_c_2087_n N_A_1278_121#_c_2368_n 0.0222946f $X=8.495 $Y=0 $X2=0
+ $Y2=0
cc_1204 N_VGND_c_2100_n N_A_1278_121#_c_2368_n 0.0112784f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1205 N_VGND_M1018_s N_A_1278_121#_c_2370_n 0.00797645f $X=8.515 $Y=0.18 $X2=0
+ $Y2=0
cc_1206 N_VGND_c_2086_n N_A_1278_121#_c_2370_n 0.0245264f $X=8.66 $Y=0 $X2=0
+ $Y2=0
cc_1207 N_VGND_c_2087_n N_A_1278_121#_c_2370_n 0.0034901f $X=8.495 $Y=0 $X2=0
+ $Y2=0
cc_1208 N_VGND_c_2088_n N_A_1278_121#_c_2370_n 0.0029521f $X=9.435 $Y=0 $X2=0
+ $Y2=0
cc_1209 N_VGND_c_2100_n N_A_1278_121#_c_2370_n 0.0115245f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1210 N_VGND_c_2079_n N_A_1278_121#_c_2372_n 0.0144673f $X=9.6 $Y=0.55 $X2=0
+ $Y2=0
cc_1211 N_VGND_c_2086_n N_A_1278_121#_c_2372_n 0.00282013f $X=8.66 $Y=0 $X2=0
+ $Y2=0
cc_1212 N_VGND_c_2088_n N_A_1278_121#_c_2372_n 0.0105866f $X=9.435 $Y=0 $X2=0
+ $Y2=0
cc_1213 N_VGND_c_2100_n N_A_1278_121#_c_2372_n 0.00888607f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1214 N_VGND_M1018_s N_A_1450_121#_c_2420_n 0.00419342f $X=8.515 $Y=0.18 $X2=0
+ $Y2=0
cc_1215 N_VGND_M1038_s N_A_1450_121#_c_2420_n 0.00176461f $X=9.46 $Y=0.37 $X2=0
+ $Y2=0
cc_1216 N_VGND_c_2079_n N_A_1450_121#_c_2420_n 0.0153337f $X=9.6 $Y=0.55 $X2=0
+ $Y2=0
cc_1217 N_VGND_c_2081_n N_A_1450_121#_c_2420_n 0.00464574f $X=10.46 $Y=0.515
+ $X2=0 $Y2=0
cc_1218 N_VGND_c_2079_n N_A_1450_121#_c_2421_n 0.0144673f $X=9.6 $Y=0.55 $X2=0
+ $Y2=0
cc_1219 N_VGND_c_2080_n N_A_1450_121#_c_2421_n 0.0109942f $X=10.295 $Y=0 $X2=0
+ $Y2=0
cc_1220 N_VGND_c_2081_n N_A_1450_121#_c_2421_n 0.0203066f $X=10.46 $Y=0.515
+ $X2=0 $Y2=0
cc_1221 N_VGND_c_2100_n N_A_1450_121#_c_2421_n 0.00904371f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1222 N_A_114_126#_c_2278_n N_A_299_126#_M1021_d 0.00316283f $X=2.14 $Y=0.875
+ $X2=-0.19 $Y2=-0.245
cc_1223 N_A_114_126#_c_2278_n N_A_299_126#_c_2324_n 0.0170749f $X=2.14 $Y=0.875
+ $X2=0 $Y2=0
cc_1224 N_A_114_126#_c_2279_n N_A_299_126#_c_2324_n 0.0289644f $X=3.05 $Y=0.842
+ $X2=0 $Y2=0
cc_1225 N_A_114_126#_c_2289_n N_A_299_126#_c_2325_n 0.0223181f $X=3.215 $Y=0.84
+ $X2=0 $Y2=0
cc_1226 N_A_114_126#_c_2279_n N_A_299_126#_c_2325_n 0.0155869f $X=3.05 $Y=0.842
+ $X2=0 $Y2=0
cc_1227 N_A_114_126#_c_2275_n N_A_299_126#_c_2327_n 8.50133e-19 $X=1.575
+ $Y=0.372 $X2=0 $Y2=0
cc_1228 N_A_114_126#_c_2278_n N_A_299_126#_c_2327_n 0.0138528f $X=2.14 $Y=0.875
+ $X2=0 $Y2=0
cc_1229 N_A_114_126#_c_2279_n N_A_299_126#_c_2328_n 0.0129027f $X=3.05 $Y=0.842
+ $X2=0 $Y2=0
cc_1230 N_A_1278_121#_c_2367_n N_A_1450_121#_c_2419_n 0.00484741f $X=8.155
+ $Y=0.34 $X2=0 $Y2=0
cc_1231 N_A_1278_121#_M1018_d N_A_1450_121#_c_2420_n 0.00176461f $X=9.03 $Y=0.37
+ $X2=0 $Y2=0
cc_1232 N_A_1278_121#_c_2370_n N_A_1450_121#_c_2420_n 0.0451131f $X=9.005
+ $Y=0.665 $X2=0 $Y2=0
cc_1233 N_A_1278_121#_c_2372_n N_A_1450_121#_c_2420_n 0.0146914f $X=9.17 $Y=0.55
+ $X2=0 $Y2=0
cc_1234 N_A_1278_121#_c_2371_n N_A_1450_121#_c_2423_n 0.0133492f $X=8.325
+ $Y=0.665 $X2=0 $Y2=0
