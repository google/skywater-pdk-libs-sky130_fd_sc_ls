* NGSPICE file created from sky130_fd_sc_ls__a21o_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_364_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.75e+11p pd=5.15e+06u as=6.38e+11p ps=5.45e+06u
M1001 VGND a_81_264# X VNB nshort w=740000u l=150000u
+  ad=4.541e+11p pd=4.09e+06u as=1.961e+11p ps=2.01e+06u
M1002 a_364_392# B1 a_81_264# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1003 VGND A2 a_452_136# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.93e+06u
M1004 a_81_264# B1 VGND VNB nshort w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1005 a_452_136# A1 a_81_264# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_364_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_81_264# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.08e+11p ps=2.79e+06u
.ends

