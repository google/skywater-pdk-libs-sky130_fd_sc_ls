* File: sky130_fd_sc_ls__dlrbn_1.spice
* Created: Wed Sep  2 11:03:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dlrbn_1.pex.spice"
.subckt sky130_fd_sc_ls__dlrbn_1  VNB VPB D GATE_N RESET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_D_M1008_g N_A_27_424#_M1008_s VNB NSHORT L=0.15 W=0.55
+ AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1006 N_A_231_74#_M1006_d N_GATE_N_M1006_g N_VGND_M1008_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_A_231_74#_M1014_g N_A_373_74#_M1014_s VNB NSHORT L=0.15
+ W=0.74 AD=0.215887 AS=0.2109 PD=1.42638 PS=2.05 NRD=30.804 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1002 A_608_74# N_A_27_424#_M1002_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.186713 PD=0.88 PS=1.23362 NRD=12.18 NRS=22.488 M=1 R=4.26667
+ SA=75000.9 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1003 N_A_686_74#_M1003_d N_A_231_74#_M1003_g A_608_74# VNB NSHORT L=0.15
+ W=0.64 AD=0.231547 AS=0.0768 PD=1.52755 PS=0.88 NRD=28.116 NRS=12.18 M=1
+ R=4.26667 SA=75001.3 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1012 A_841_118# N_A_373_74#_M1012_g N_A_686_74#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.151953 PD=0.66 PS=1.00245 NRD=18.564 NRS=57.132 M=1
+ R=2.8 SA=75002.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_889_92#_M1020_g A_841_118# VNB NSHORT L=0.15 W=0.42
+ AD=0.1533 AS=0.0504 PD=1.57 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8 SA=75002.5
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1015 A_1133_74# N_A_686_74#_M1015_g N_A_889_92#_M1015_s VNB NSHORT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_RESET_B_M1007_g A_1133_74# VNB NSHORT L=0.15 W=0.74
+ AD=0.1443 AS=0.0888 PD=1.13 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1017 N_Q_M1017_d N_A_889_92#_M1017_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1443 PD=2.05 PS=1.13 NRD=0 NRS=17.832 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_889_92#_M1010_g N_A_1437_112#_M1010_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.109083 AS=0.1925 PD=0.942248 PS=1.8 NRD=19.08 NRS=0 M=1
+ R=3.66667 SA=75000.3 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1019 N_Q_N_M1019_d N_A_1437_112#_M1019_g N_VGND_M1010_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.146767 PD=2.05 PS=1.26775 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_VPWR_M1016_d N_D_M1016_g N_A_27_424#_M1016_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2562 AS=0.2478 PD=1.45 PS=2.27 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75001 A=0.126 P=1.98 MULT=1
MM1018 N_A_231_74#_M1018_d N_GATE_N_M1018_g N_VPWR_M1016_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.2562 PD=2.27 PS=1.45 NRD=2.3443 NRS=75.0373 M=1 R=5.6
+ SA=75001 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_A_231_74#_M1009_g N_A_373_74#_M1009_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.230498 AS=0.383 PD=1.49739 PS=2.88 NRD=51.4367 NRS=23.443 M=1
+ R=5.6 SA=75000.3 SB=75002.2 A=0.126 P=1.98 MULT=1
MM1000 A_611_392# N_A_27_424#_M1000_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.274402 PD=1.27 PS=1.78261 NRD=15.7403 NRS=19.6803 M=1 R=6.66667
+ SA=75000.8 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1022 N_A_686_74#_M1022_d N_A_373_74#_M1022_g A_611_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.234366 AS=0.135 PD=1.9507 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75001.2 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1005 A_802_508# N_A_231_74#_M1005_g N_A_686_74#_M1022_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.11235 AS=0.0984338 PD=0.955 PS=0.819296 NRD=99.6623 NRS=46.886 M=1
+ R=2.8 SA=75001.6 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_889_92#_M1004_g A_802_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.130677 AS=0.11235 PD=1.10455 PS=0.955 NRD=4.6886 NRS=99.6623 M=1 R=2.8
+ SA=75002.3 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1021 N_A_889_92#_M1021_d N_A_686_74#_M1021_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.1736 AS=0.348473 PD=1.43 PS=2.94545 NRD=3.5066 NRS=8.7862 M=1
+ R=7.46667 SA=75001 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1023 N_VPWR_M1023_d N_RESET_B_M1023_g N_A_889_92#_M1021_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.2128 AS=0.1736 PD=1.5 PS=1.43 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1013 N_Q_M1013_d N_A_889_92#_M1013_g N_VPWR_M1023_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3248 AS=0.2128 PD=2.82 PS=1.5 NRD=4.3931 NRS=7.0329 M=1 R=7.46667
+ SA=75002 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_889_92#_M1011_g N_A_1437_112#_M1011_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1734 AS=0.231 PD=1.29429 PS=2.23 NRD=42.7884 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1001 N_Q_N_M1001_d N_A_1437_112#_M1001_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.2312 PD=2.83 PS=1.72571 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX24_noxref VNB VPB NWDIODE A=17.3933 P=22.02
c_79 VNB 0 5.58535e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__dlrbn_1.pxi.spice"
*
.ends
*
*
