* File: sky130_fd_sc_ls__o31ai_1.spice
* Created: Wed Sep  2 11:22:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o31ai_1.pex.spice"
.subckt sky130_fd_sc_ls__o31ai_1  VNB VPB A1 A2 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 N_A_114_74#_M1005_d N_A1_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_114_74#_M1005_d VNB NSHORT L=0.15 W=0.74
+ AD=0.3492 AS=0.1036 PD=1.7 PS=1.02 NRD=13.776 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1000 N_A_114_74#_M1000_d N_A3_M1000_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.74
+ AD=0.111 AS=0.3492 PD=1.04 PS=1.7 NRD=0 NRS=13.776 M=1 R=4.93333 SA=75001.6
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g N_A_114_74#_M1000_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2479 AS=0.111 PD=2.15 PS=1.04 NRD=8.1 NRS=3.24 M=1 R=4.93333 SA=75002.1
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1001 A_119_368# N_A1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1512 AS=0.3304 PD=1.39 PS=2.83 NRD=14.0658 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002 A=0.168 P=2.54 MULT=1
MM1007 A_203_368# N_A2_M1007_g A_119_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.2352
+ AS=0.1512 PD=1.54 PS=1.39 NRD=27.2451 NRS=14.0658 M=1 R=7.46667 SA=75000.6
+ SB=75001.6 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1004_d N_A3_M1004_g A_203_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.3864
+ AS=0.2352 PD=1.81 PS=1.54 NRD=1.7533 NRS=27.2451 M=1 R=7.46667 SA=75001.2
+ SB=75001.1 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1002_d N_B1_M1002_g N_Y_M1004_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.3864 PD=2.83 PS=1.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ls__o31ai_1.pxi.spice"
*
.ends
*
*
