* File: sky130_fd_sc_ls__sdfsbp_2.pex.spice
* Created: Wed Sep  2 11:27:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%A_27_74# 1 2 9 10 12 15 18 21 25 26 28 30
+ 31 33 39
c77 33 0 1.76481e-19 $X=1.94 $Y=1.975
r78 33 36 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.94 $Y=1.975 $X2=1.94
+ $Y2=2.055
r79 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=1.975 $X2=1.94 $Y2=1.975
r80 29 31 3.11956 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.465 $Y=2.055
+ $X2=0.275 $Y2=2.055
r81 28 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=2.055
+ $X2=1.94 $Y2=2.055
r82 28 29 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=1.775 $Y=2.055
+ $X2=0.465 $Y2=2.055
r83 26 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.065
+ $X2=0.98 $Y2=0.9
r84 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.98
+ $Y=1.065 $X2=0.98 $Y2=1.065
r85 23 30 0.565906 $w=3.3e-07 $l=1.8e-07 $layer=LI1_cond $X=0.445 $Y=1.065
+ $X2=0.265 $Y2=1.065
r86 23 25 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=0.445 $Y=1.065
+ $X2=0.98 $Y2=1.065
r87 19 31 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.275 $Y=2.14
+ $X2=0.275 $Y2=2.055
r88 19 21 9.85642 $w=3.78e-07 $l=3.25e-07 $layer=LI1_cond $X=0.275 $Y=2.14
+ $X2=0.275 $Y2=2.465
r89 18 31 3.40559 $w=2.75e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.17 $Y=1.97
+ $X2=0.275 $Y2=2.055
r90 17 30 6.17543 $w=2.65e-07 $l=2.07123e-07 $layer=LI1_cond $X=0.17 $Y=1.23
+ $X2=0.265 $Y2=1.065
r91 17 18 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.17 $Y=1.23
+ $X2=0.17 $Y2=1.97
r92 13 30 6.17543 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=0.9
+ $X2=0.265 $Y2=1.065
r93 13 15 10.2439 $w=3.58e-07 $l=3.2e-07 $layer=LI1_cond $X=0.265 $Y=0.9
+ $X2=0.265 $Y2=0.58
r94 10 34 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=2.015 $Y=2.245
+ $X2=1.94 $Y2=1.975
r95 10 12 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.015 $Y=2.245
+ $X2=2.015 $Y2=2.64
r96 9 39 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.07 $Y=0.58 $X2=1.07
+ $Y2=0.9
r97 2 21 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.155
+ $Y=2.32 $X2=0.3 $Y2=2.465
r98 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%SCE 3 6 7 9 11 12 14 17 20 23 24 25 27 34
+ 35 36
c84 34 0 1.76481e-19 $X=2.13 $Y=1.065
r85 34 36 46.8261 $w=5.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.22 $Y=1.065
+ $X2=2.22 $Y2=0.9
r86 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.13
+ $Y=1.065 $X2=2.13 $Y2=1.065
r87 29 30 4.49068 $w=3.22e-07 $l=3e-08 $layer=POLY_cond $X=0.495 $Y=1.635
+ $X2=0.525 $Y2=1.635
r88 27 35 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.13 $Y=1.295
+ $X2=2.13 $Y2=1.065
r89 26 27 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.13 $Y=1.4
+ $X2=2.13 $Y2=1.295
r90 24 32 15.7174 $w=3.22e-07 $l=1.05e-07 $layer=POLY_cond $X=0.92 $Y=1.635
+ $X2=1.025 $Y2=1.635
r91 24 30 59.1273 $w=3.22e-07 $l=3.95e-07 $layer=POLY_cond $X=0.92 $Y=1.635
+ $X2=0.525 $Y2=1.635
r92 23 25 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.92 $Y=1.6
+ $X2=1.085 $Y2=1.6
r93 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.92
+ $Y=1.635 $X2=0.92 $Y2=1.635
r94 20 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.965 $Y=1.485
+ $X2=2.13 $Y2=1.4
r95 20 25 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=1.965 $Y=1.485
+ $X2=1.085 $Y2=1.485
r96 17 36 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.4 $Y=0.58 $X2=2.4
+ $Y2=0.9
r97 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.025 $Y=2.245
+ $X2=1.025 $Y2=2.64
r98 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.025 $Y=2.155
+ $X2=1.025 $Y2=2.245
r99 10 32 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.025 $Y=1.8
+ $X2=1.025 $Y2=1.635
r100 10 11 137.992 $w=1.8e-07 $l=3.55e-07 $layer=POLY_cond $X=1.025 $Y=1.8
+ $X2=1.025 $Y2=2.155
r101 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.525 $Y=2.245
+ $X2=0.525 $Y2=2.64
r102 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.525 $Y=2.155
+ $X2=0.525 $Y2=2.245
r103 5 30 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.8
+ $X2=0.525 $Y2=1.635
r104 5 6 137.992 $w=1.8e-07 $l=3.55e-07 $layer=POLY_cond $X=0.525 $Y=1.8
+ $X2=0.525 $Y2=2.155
r105 1 29 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.47
+ $X2=0.495 $Y2=1.635
r106 1 3 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=0.495 $Y=1.47
+ $X2=0.495 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%D 1 2 3 5 8 11 12 13 17 19
r49 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.55 $Y=1.065
+ $X2=1.55 $Y2=1.23
r50 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.55 $Y=1.065
+ $X2=1.55 $Y2=0.9
r51 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=1.065 $X2=1.55 $Y2=1.065
r52 13 18 3.93517 $w=4.08e-07 $l=1.4e-07 $layer=LI1_cond $X=1.59 $Y=0.925
+ $X2=1.59 $Y2=1.065
r53 12 13 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.59 $Y=0.555
+ $X2=1.59 $Y2=0.925
r54 11 20 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.46 $Y=1.47
+ $X2=1.46 $Y2=1.23
r55 8 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.46 $Y=0.58 $X2=1.46
+ $Y2=0.9
r56 3 5 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.445 $Y=2.245
+ $X2=1.445 $Y2=2.64
r57 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.445 $Y=2.155 $X2=1.445
+ $Y2=2.245
r58 1 11 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.445 $Y=1.56 $X2=1.445
+ $Y2=1.47
r59 1 2 231.282 $w=1.8e-07 $l=5.95e-07 $layer=POLY_cond $X=1.445 $Y=1.56
+ $X2=1.445 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%SCD 2 3 5 6 7 10 13 15 16 17 20
r52 20 22 46.1517 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.925 $Y=1.115
+ $X2=2.925 $Y2=0.95
r53 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.97
+ $Y=1.115 $X2=2.97 $Y2=1.115
r54 17 21 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.12 $Y=1.285
+ $X2=2.97 $Y2=1.285
r55 15 16 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.79 $Y=1.81
+ $X2=2.79 $Y2=1.62
r56 13 16 52.1105 $w=4.2e-07 $l=2.1e-07 $layer=POLY_cond $X=2.925 $Y=1.41
+ $X2=2.925 $Y2=1.62
r57 12 20 5.95879 $w=4.2e-07 $l=4.5e-08 $layer=POLY_cond $X=2.925 $Y=1.16
+ $X2=2.925 $Y2=1.115
r58 12 13 33.1044 $w=4.2e-07 $l=2.5e-07 $layer=POLY_cond $X=2.925 $Y=1.16
+ $X2=2.925 $Y2=1.41
r59 10 22 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.79 $Y=0.58
+ $X2=2.79 $Y2=0.95
r60 6 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.715 $Y=1.885
+ $X2=2.79 $Y2=1.81
r61 6 7 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.715 $Y=1.885
+ $X2=2.525 $Y2=1.885
r62 3 5 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.435 $Y=2.245
+ $X2=2.435 $Y2=2.64
r63 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.435 $Y=2.155 $X2=2.435
+ $Y2=2.245
r64 1 7 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.435 $Y=1.96
+ $X2=2.525 $Y2=1.885
r65 1 2 75.7984 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=2.435 $Y=1.96
+ $X2=2.435 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%CLK 1 3 4 6 7
c34 4 0 9.27061e-20 $X=3.78 $Y=1.22
c35 1 0 1.34113e-19 $X=3.465 $Y=1.765
r36 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.83
+ $Y=1.385 $X2=3.83 $Y2=1.385
r37 7 11 7.78678 $w=3.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.08 $Y=1.365
+ $X2=3.83 $Y2=1.365
r38 4 10 40.5859 $w=4.46e-07 $l=2.07123e-07 $layer=POLY_cond $X=3.78 $Y=1.22
+ $X2=3.685 $Y2=1.385
r39 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.78 $Y=1.22 $X2=3.78
+ $Y2=0.74
r40 1 10 63.8213 $w=4.46e-07 $l=4.77493e-07 $layer=POLY_cond $X=3.465 $Y=1.765
+ $X2=3.685 $Y2=1.385
r41 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.465 $Y=1.765
+ $X2=3.465 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%A_871_74# 1 2 8 9 11 12 13 16 20 24 26 27
+ 28 31 32 34 37 40 44 46 47 48 49 52 53 59 60 63 64 67 68 69 71 72 73 75 77 80
+ 83 86 87 88 98
c272 87 0 1.69669e-19 $X=6.187 $Y=2.25
c273 83 0 1.33892e-19 $X=11.225 $Y=1.365
c274 80 0 7.75954e-20 $X=10.545 $Y=1.365
c275 73 0 1.56558e-19 $X=8.165 $Y=2.135
c276 59 0 1.02354e-19 $X=6.185 $Y=1.135
c277 47 0 9.27061e-20 $X=4.66 $Y=0.34
c278 46 0 1.10104e-19 $X=5.39 $Y=0.34
c279 37 0 1.21895e-19 $X=5.395 $Y=1.96
c280 9 0 3.32958e-20 $X=5.43 $Y=2.24
c281 8 0 6.21188e-20 $X=5.43 $Y=2.15
r282 84 98 46.1517 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=11.225 $Y=1.41
+ $X2=11.39 $Y2=1.41
r283 83 84 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=11.225
+ $Y=1.365 $X2=11.225 $Y2=1.365
r284 81 96 30.5693 $w=3.39e-07 $l=2.15e-07 $layer=POLY_cond $X=10.545 $Y=1.41
+ $X2=10.76 $Y2=1.41
r285 80 88 8.03587 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.545 $Y=1.365
+ $X2=10.38 $Y2=1.365
r286 80 83 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=10.545 $Y=1.365
+ $X2=11.225 $Y2=1.365
r287 80 81 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=10.545
+ $Y=1.365 $X2=10.545 $Y2=1.365
r288 77 88 118.412 $w=1.68e-07 $l=1.815e-06 $layer=LI1_cond $X=8.565 $Y=1.43
+ $X2=10.38 $Y2=1.43
r289 74 77 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.48 $Y=1.515
+ $X2=8.565 $Y2=1.43
r290 74 75 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=8.48 $Y=1.515
+ $X2=8.48 $Y2=2.05
r291 72 75 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.395 $Y=2.135
+ $X2=8.48 $Y2=2.05
r292 72 73 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=8.395 $Y=2.135
+ $X2=8.165 $Y2=2.135
r293 70 73 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.08 $Y=2.22
+ $X2=8.165 $Y2=2.135
r294 70 71 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=8.08 $Y=2.22
+ $X2=8.08 $Y2=2.905
r295 68 71 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.995 $Y=2.99
+ $X2=8.08 $Y2=2.905
r296 68 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.995 $Y=2.99
+ $X2=7.325 $Y2=2.99
r297 67 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.24 $Y=2.905
+ $X2=7.325 $Y2=2.99
r298 66 67 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.24 $Y=2.335
+ $X2=7.24 $Y2=2.905
r299 65 87 1.97946 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=6.305 $Y=2.25
+ $X2=6.187 $Y2=2.25
r300 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.155 $Y=2.25
+ $X2=7.24 $Y2=2.335
r301 64 65 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=7.155 $Y=2.25
+ $X2=6.305 $Y2=2.25
r302 62 87 4.45556 $w=2.02e-07 $l=9.97246e-08 $layer=LI1_cond $X=6.155 $Y=2.335
+ $X2=6.187 $Y2=2.25
r303 62 63 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.155 $Y=2.335
+ $X2=6.155 $Y2=2.905
r304 60 92 37.9199 $w=3.5e-07 $l=2.3e-07 $layer=POLY_cond $X=6.195 $Y=1.135
+ $X2=6.195 $Y2=1.365
r305 60 91 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.195 $Y=1.135
+ $X2=6.195 $Y2=0.97
r306 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.185
+ $Y=1.135 $X2=6.185 $Y2=1.135
r307 57 87 4.45556 $w=2.02e-07 $l=8.5e-08 $layer=LI1_cond $X=6.187 $Y=2.165
+ $X2=6.187 $Y2=2.25
r308 57 59 50.5113 $w=2.33e-07 $l=1.03e-06 $layer=LI1_cond $X=6.187 $Y=2.165
+ $X2=6.187 $Y2=1.135
r309 55 86 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=5.475 $Y=0.425
+ $X2=5.475 $Y2=1.29
r310 52 86 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.395 $Y=1.455
+ $X2=5.395 $Y2=1.29
r311 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.395
+ $Y=1.455 $X2=5.395 $Y2=1.455
r312 48 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.07 $Y=2.99
+ $X2=6.155 $Y2=2.905
r313 48 49 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=6.07 $Y=2.99
+ $X2=4.72 $Y2=2.99
r314 46 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.39 $Y=0.34
+ $X2=5.475 $Y2=0.425
r315 46 47 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.39 $Y=0.34
+ $X2=4.66 $Y2=0.34
r316 42 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.555 $Y=2.905
+ $X2=4.72 $Y2=2.99
r317 42 44 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=4.555 $Y=2.905
+ $X2=4.555 $Y2=2.725
r318 38 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.495 $Y=0.425
+ $X2=4.66 $Y2=0.34
r319 38 40 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.495 $Y=0.425
+ $X2=4.495 $Y2=0.505
r320 36 53 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.395 $Y=1.795
+ $X2=5.395 $Y2=1.455
r321 36 37 36.5727 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.395 $Y=1.795
+ $X2=5.395 $Y2=1.96
r322 35 53 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.395 $Y=1.44
+ $X2=5.395 $Y2=1.455
r323 32 34 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.76 $Y=2.2
+ $X2=11.76 $Y2=2.485
r324 31 32 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.76 $Y=2.11
+ $X2=11.76 $Y2=2.2
r325 30 31 190.468 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=11.76 $Y=1.62
+ $X2=11.76 $Y2=2.11
r326 28 30 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=11.67 $Y=1.545
+ $X2=11.76 $Y2=1.62
r327 28 98 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=11.67 $Y=1.545
+ $X2=11.39 $Y2=1.545
r328 27 96 10.5406 $w=4.2e-07 $l=7.5e-08 $layer=POLY_cond $X=10.835 $Y=1.41
+ $X2=10.76 $Y2=1.41
r329 26 84 5.95879 $w=4.2e-07 $l=4.5e-08 $layer=POLY_cond $X=11.18 $Y=1.41
+ $X2=11.225 $Y2=1.41
r330 26 27 45.6841 $w=4.2e-07 $l=3.45e-07 $layer=POLY_cond $X=11.18 $Y=1.41
+ $X2=10.835 $Y2=1.41
r331 22 96 21.8644 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=10.76 $Y=1.2
+ $X2=10.76 $Y2=1.41
r332 22 24 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=10.76 $Y=1.2
+ $X2=10.76 $Y2=0.69
r333 18 81 40.5221 $w=3.39e-07 $l=3.756e-07 $layer=POLY_cond $X=10.26 $Y=1.2
+ $X2=10.545 $Y2=1.41
r334 18 20 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=10.26 $Y=1.2
+ $X2=10.26 $Y2=0.69
r335 16 91 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=6.295 $Y=0.615
+ $X2=6.295 $Y2=0.97
r336 13 35 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.56 $Y=1.365
+ $X2=5.395 $Y2=1.44
r337 12 92 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.02 $Y=1.365
+ $X2=6.195 $Y2=1.365
r338 12 13 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=6.02 $Y=1.365
+ $X2=5.56 $Y2=1.365
r339 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.43 $Y=2.24 $X2=5.43
+ $Y2=2.525
r340 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.43 $Y=2.15 $X2=5.43
+ $Y2=2.24
r341 8 37 73.8548 $w=1.8e-07 $l=1.9e-07 $layer=POLY_cond $X=5.43 $Y=2.15
+ $X2=5.43 $Y2=1.96
r342 2 44 600 $w=1.7e-07 $l=9.73114e-07 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=1.84 $X2=4.555 $Y2=2.725
r343 1 40 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=4.355
+ $Y=0.37 $X2=4.495 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%A_1252_376# 1 2 7 9 10 12 14 17 19 22 24 28
+ 32 39 40 43 47
c91 47 0 1.02354e-19 $X=6.89 $Y=1.1
c92 24 0 1.50114e-19 $X=7.38 $Y=0.955
c93 22 0 1.15615e-19 $X=6.8 $Y=1.865
c94 7 0 7.37914e-20 $X=6.35 $Y=2.24
r95 39 40 10.3829 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=7.66 $Y=2.515
+ $X2=7.66 $Y2=2.295
r96 36 47 16.6207 $w=2.61e-07 $l=9e-08 $layer=POLY_cond $X=6.98 $Y=1.1 $X2=6.89
+ $Y2=1.1
r97 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.98
+ $Y=1.1 $X2=6.98 $Y2=1.1
r98 32 35 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=6.98 $Y=0.955
+ $X2=6.98 $Y2=1.1
r99 30 40 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.58 $Y=1.995 $X2=7.58
+ $Y2=2.295
r100 26 28 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=7.545 $Y=0.87
+ $X2=7.545 $Y2=0.58
r101 25 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.145 $Y=0.955
+ $X2=6.98 $Y2=0.955
r102 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.38 $Y=0.955
+ $X2=7.545 $Y2=0.87
r103 24 25 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=7.38 $Y=0.955
+ $X2=7.145 $Y2=0.955
r104 22 44 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.8 $Y=1.865 $X2=6.8
+ $Y2=1.955
r105 22 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.8 $Y=1.865
+ $X2=6.8 $Y2=1.7
r106 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.8
+ $Y=1.865 $X2=6.8 $Y2=1.865
r107 19 30 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.495 $Y=1.865
+ $X2=7.58 $Y2=1.995
r108 19 21 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=7.495 $Y=1.865
+ $X2=6.8 $Y2=1.865
r109 15 47 15.717 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.89 $Y=1.265
+ $X2=6.89 $Y2=1.1
r110 15 43 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.89 $Y=1.265
+ $X2=6.89 $Y2=1.7
r111 12 47 37.8582 $w=2.61e-07 $l=2.75409e-07 $layer=POLY_cond $X=6.685 $Y=0.935
+ $X2=6.89 $Y2=1.1
r112 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.685 $Y=0.935
+ $X2=6.685 $Y2=0.615
r113 11 17 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.44 $Y=1.955 $X2=6.35
+ $Y2=1.955
r114 10 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.635 $Y=1.955
+ $X2=6.8 $Y2=1.955
r115 10 11 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=6.635 $Y=1.955
+ $X2=6.44 $Y2=1.955
r116 7 17 112.932 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.35 $Y=2.24
+ $X2=6.35 $Y2=1.955
r117 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.35 $Y=2.24 $X2=6.35
+ $Y2=2.525
r118 2 39 600 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_PDIFF $count=1 $X=7.51
+ $Y=2.315 $X2=7.66 $Y2=2.515
r119 1 28 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=7.4
+ $Y=0.37 $X2=7.545 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%A_1069_81# 1 2 8 9 11 14 16 19 20 22 25 26
+ 29 30 32 35 37 38 40 43 44 48 49 50 51 53 55 56 59 60 62 66
c187 62 0 4.48044e-20 $X=7.51 $Y=1.295
c188 60 0 7.37914e-20 $X=5.72 $Y=2.295
c189 59 0 1.21895e-19 $X=5.705 $Y=2.515
c190 50 0 1.15615e-19 $X=6.645 $Y=1.48
c191 37 0 1.14148e-19 $X=9.365 $Y=1.16
c192 29 0 7.75954e-20 $X=9.815 $Y=1.955
c193 20 0 3.30716e-19 $X=9.365 $Y=2.045
c194 8 0 1.56558e-19 $X=7.435 $Y=2.15
r195 66 73 12.1213 $w=3.38e-07 $l=8.5e-08 $layer=POLY_cond $X=7.52 $Y=1.4
+ $X2=7.435 $Y2=1.4
r196 65 67 3.90344 $w=3.08e-07 $l=1.05e-07 $layer=LI1_cond $X=7.51 $Y=1.375
+ $X2=7.51 $Y2=1.48
r197 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.52
+ $Y=1.375 $X2=7.52 $Y2=1.375
r198 62 65 2.97405 $w=3.08e-07 $l=8e-08 $layer=LI1_cond $X=7.51 $Y=1.295
+ $X2=7.51 $Y2=1.375
r199 59 60 10.2717 $w=3.58e-07 $l=2.2e-07 $layer=LI1_cond $X=5.72 $Y=2.515
+ $X2=5.72 $Y2=2.295
r200 56 78 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=8.695 $Y=1.065
+ $X2=8.695 $Y2=1.16
r201 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.695
+ $Y=1.065 $X2=8.695 $Y2=1.065
r202 53 71 16.8321 $w=1.68e-07 $l=2.58e-07 $layer=LI1_cond $X=7.965 $Y=1.037
+ $X2=7.965 $Y2=1.295
r203 53 55 27.03 $w=2.73e-07 $l=6.45e-07 $layer=LI1_cond $X=8.05 $Y=1.037
+ $X2=8.695 $Y2=1.037
r204 52 62 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=7.665 $Y=1.295
+ $X2=7.51 $Y2=1.295
r205 51 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.88 $Y=1.295
+ $X2=7.965 $Y2=1.295
r206 51 52 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.88 $Y=1.295
+ $X2=7.665 $Y2=1.295
r207 49 67 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=7.355 $Y=1.48
+ $X2=7.51 $Y2=1.48
r208 49 50 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.355 $Y=1.48
+ $X2=6.645 $Y2=1.48
r209 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.56 $Y=1.395
+ $X2=6.645 $Y2=1.48
r210 47 48 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=6.56 $Y=0.8
+ $X2=6.56 $Y2=1.395
r211 44 46 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=0.635
+ $X2=5.985 $Y2=0.635
r212 43 47 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.475 $Y=0.635
+ $X2=6.56 $Y2=0.8
r213 43 46 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=6.475 $Y=0.635
+ $X2=5.985 $Y2=0.635
r214 41 44 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.815 $Y=0.8
+ $X2=5.9 $Y2=0.635
r215 41 60 97.5348 $w=1.68e-07 $l=1.495e-06 $layer=LI1_cond $X=5.815 $Y=0.8
+ $X2=5.815 $Y2=2.295
r216 37 39 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=9.365 $Y=1.16
+ $X2=9.365 $Y2=1.31
r217 37 38 31.303 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.365 $Y=1.16
+ $X2=9.365 $Y2=1.085
r218 33 40 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=9.83 $Y=1.235
+ $X2=9.815 $Y2=1.31
r219 33 35 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=9.83 $Y=1.235
+ $X2=9.83 $Y2=0.69
r220 30 32 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.815 $Y=2.045
+ $X2=9.815 $Y2=2.54
r221 29 30 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.815 $Y=1.955
+ $X2=9.815 $Y2=2.045
r222 28 40 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=9.815 $Y=1.385
+ $X2=9.815 $Y2=1.31
r223 28 29 221.565 $w=1.8e-07 $l=5.7e-07 $layer=POLY_cond $X=9.815 $Y=1.385
+ $X2=9.815 $Y2=1.955
r224 27 39 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.455 $Y=1.31
+ $X2=9.365 $Y2=1.31
r225 26 40 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.725 $Y=1.31
+ $X2=9.815 $Y2=1.31
r226 26 27 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.725 $Y=1.31
+ $X2=9.455 $Y2=1.31
r227 25 38 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=9.38 $Y=0.69
+ $X2=9.38 $Y2=1.085
r228 20 22 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.365 $Y=2.045
+ $X2=9.365 $Y2=2.54
r229 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.365 $Y=1.955
+ $X2=9.365 $Y2=2.045
r230 18 39 29.1532 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.365 $Y=1.385
+ $X2=9.365 $Y2=1.31
r231 18 19 221.565 $w=1.8e-07 $l=5.7e-07 $layer=POLY_cond $X=9.365 $Y=1.385
+ $X2=9.365 $Y2=1.955
r232 17 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.86 $Y=1.16
+ $X2=8.695 $Y2=1.16
r233 16 37 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.275 $Y=1.16
+ $X2=9.365 $Y2=1.16
r234 16 17 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=9.275 $Y=1.16
+ $X2=8.86 $Y2=1.16
r235 12 66 34.2249 $w=3.38e-07 $l=3.39411e-07 $layer=POLY_cond $X=7.76 $Y=1.16
+ $X2=7.52 $Y2=1.4
r236 12 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.76 $Y=1.16
+ $X2=7.76 $Y2=0.58
r237 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.435 $Y=2.24
+ $X2=7.435 $Y2=2.525
r238 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.435 $Y=2.15 $X2=7.435
+ $Y2=2.24
r239 7 73 17.4907 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=7.435 $Y=1.64
+ $X2=7.435 $Y2=1.4
r240 7 8 198.242 $w=1.8e-07 $l=5.1e-07 $layer=POLY_cond $X=7.435 $Y=1.64
+ $X2=7.435 $Y2=2.15
r241 2 59 600 $w=1.7e-07 $l=2.82843e-07 $layer=licon1_PDIFF $count=1 $X=5.505
+ $Y=2.315 $X2=5.705 $Y2=2.515
r242 1 46 182 $w=1.7e-07 $l=7.4619e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.405 $X2=5.985 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%SET_B 2 3 5 8 12 15 16 18 21 22 23 24 27 29
+ 32 33 35
c150 35 0 4.48044e-20 $X=8.06 $Y=1.715
c151 8 0 1.50114e-19 $X=8.15 $Y=0.58
r152 35 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.06 $Y=1.715
+ $X2=8.06 $Y2=1.88
r153 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.06 $Y=1.715
+ $X2=8.06 $Y2=1.55
r154 33 43 1.24963 $w=6.68e-07 $l=7e-08 $layer=LI1_cond $X=13.27 $Y=1.635
+ $X2=13.2 $Y2=1.635
r155 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.27
+ $Y=1.465 $X2=13.27 $Y2=1.465
r156 29 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=1.665
+ $X2=13.2 $Y2=1.665
r157 27 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.06
+ $Y=1.715 $X2=8.06 $Y2=1.715
r158 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=1.665
+ $X2=7.92 $Y2=1.665
r159 24 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=1.665
+ $X2=7.92 $Y2=1.665
r160 23 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.055 $Y=1.665
+ $X2=13.2 $Y2=1.665
r161 23 24 6.17573 $w=1.4e-07 $l=4.99e-06 $layer=MET1_cond $X=13.055 $Y=1.665
+ $X2=8.065 $Y2=1.665
r162 21 32 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=13.27 $Y=1.805
+ $X2=13.27 $Y2=1.465
r163 21 22 35.6818 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.27 $Y=1.805
+ $X2=13.27 $Y2=1.97
r164 20 32 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.27 $Y=1.3
+ $X2=13.27 $Y2=1.465
r165 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.25 $Y=2.465
+ $X2=13.25 $Y2=2.75
r166 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=13.25 $Y=2.375
+ $X2=13.25 $Y2=2.465
r167 15 22 157.427 $w=1.8e-07 $l=4.05e-07 $layer=POLY_cond $X=13.25 $Y=2.375
+ $X2=13.25 $Y2=1.97
r168 12 20 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=13.21 $Y=0.58
+ $X2=13.21 $Y2=1.3
r169 8 37 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=8.15 $Y=0.58
+ $X2=8.15 $Y2=1.55
r170 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.985 $Y=2.24
+ $X2=7.985 $Y2=2.525
r171 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.985 $Y=2.15 $X2=7.985
+ $Y2=2.24
r172 2 38 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=7.985 $Y=2.15
+ $X2=7.985 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%A_619_368# 1 2 9 11 13 15 17 18 19 20 21 22
+ 24 25 26 27 29 30 33 34 36 37 38 39 41 42 45 46 47 48 49 50 52 54 55 56 57 58
+ 60 63 66 67 71 74 78 85 86 89 91
c276 78 0 1.49424e-19 $X=11.885 $Y=1.065
c277 71 0 1.34113e-19 $X=4.555 $Y=1.515
c278 60 0 1.33892e-19 $X=12.205 $Y=1.065
c279 49 0 1.00509e-19 $X=12.28 $Y=3.065
c280 42 0 7.33293e-20 $X=11.16 $Y=1.97
c281 22 0 9.15331e-20 $X=5.27 $Y=0.9
c282 18 0 1.10104e-19 $X=5.195 $Y=0.975
c283 17 0 9.36703e-20 $X=4.85 $Y=3.075
r284 89 95 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=8.9 $Y=1.795
+ $X2=8.795 $Y2=1.795
r285 88 91 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=8.9 $Y=1.822
+ $X2=9.065 $Y2=1.822
r286 88 89 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.9
+ $Y=1.795 $X2=8.9 $Y2=1.795
r287 84 85 5.85433 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=1.965
+ $X2=3.545 $Y2=1.965
r288 82 84 7.24393 $w=3.48e-07 $l=2.2e-07 $layer=LI1_cond $X=3.24 $Y=1.965
+ $X2=3.46 $Y2=1.965
r289 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.885
+ $Y=1.065 $X2=11.885 $Y2=1.065
r290 76 78 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=11.885 $Y=1.7
+ $X2=11.885 $Y2=1.065
r291 74 76 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.72 $Y=1.785
+ $X2=11.885 $Y2=1.7
r292 74 91 173.214 $w=1.68e-07 $l=2.655e-06 $layer=LI1_cond $X=11.72 $Y=1.785
+ $X2=9.065 $Y2=1.785
r293 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.555
+ $Y=1.515 $X2=4.555 $Y2=1.515
r294 69 71 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.555 $Y=1.79
+ $X2=4.555 $Y2=1.515
r295 67 69 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.39 $Y=1.875
+ $X2=4.555 $Y2=1.79
r296 67 85 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=4.39 $Y=1.875
+ $X2=3.545 $Y2=1.875
r297 66 84 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.46 $Y=1.79 $X2=3.46
+ $Y2=1.965
r298 66 86 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.46 $Y=1.79
+ $X2=3.46 $Y2=1.01
r299 61 86 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=3.512 $Y=0.873
+ $X2=3.512 $Y2=1.01
r300 61 63 15.4218 $w=2.73e-07 $l=3.68e-07 $layer=LI1_cond $X=3.512 $Y=0.873
+ $X2=3.512 $Y2=0.505
r301 60 79 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=12.205 $Y=1.065
+ $X2=11.885 $Y2=1.065
r302 55 72 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=4.775 $Y=1.515
+ $X2=4.555 $Y2=1.515
r303 55 56 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.775 $Y=1.515
+ $X2=4.85 $Y2=1.515
r304 53 72 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=4.385 $Y=1.515
+ $X2=4.555 $Y2=1.515
r305 53 54 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=4.385 $Y=1.515
+ $X2=4.295 $Y2=1.557
r306 50 60 41.2111 $w=2.18e-07 $l=1.98997e-07 $layer=POLY_cond $X=12.43 $Y=0.9
+ $X2=12.355 $Y2=1.065
r307 50 52 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=12.43 $Y=0.9
+ $X2=12.43 $Y2=0.58
r308 48 60 41.2111 $w=2.18e-07 $l=1.98997e-07 $layer=POLY_cond $X=12.28 $Y=1.23
+ $X2=12.355 $Y2=1.065
r309 48 49 940.926 $w=1.5e-07 $l=1.835e-06 $layer=POLY_cond $X=12.28 $Y=1.23
+ $X2=12.28 $Y2=3.065
r310 46 49 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.205 $Y=3.14
+ $X2=12.28 $Y2=3.065
r311 46 47 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=12.205 $Y=3.14
+ $X2=11.31 $Y2=3.14
r312 45 47 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.235 $Y=3.065
+ $X2=11.31 $Y2=3.14
r313 44 45 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=11.235 $Y=2.045
+ $X2=11.235 $Y2=3.065
r314 43 58 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.79 $Y=1.97
+ $X2=10.715 $Y2=1.97
r315 42 44 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.16 $Y=1.97
+ $X2=11.235 $Y2=2.045
r316 42 43 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=11.16 $Y=1.97
+ $X2=10.79 $Y2=1.97
r317 39 58 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.715 $Y=2.045
+ $X2=10.715 $Y2=1.97
r318 39 41 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.715 $Y=2.045
+ $X2=10.715 $Y2=2.54
r319 37 58 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.64 $Y=1.97
+ $X2=10.715 $Y2=1.97
r320 37 38 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=10.64 $Y=1.97
+ $X2=10.34 $Y2=1.97
r321 34 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.265 $Y=2.045
+ $X2=10.34 $Y2=1.97
r322 34 36 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.265 $Y=2.045
+ $X2=10.265 $Y2=2.54
r323 32 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.795 $Y=1.96
+ $X2=8.795 $Y2=1.795
r324 32 33 571.734 $w=1.5e-07 $l=1.115e-06 $layer=POLY_cond $X=8.795 $Y=1.96
+ $X2=8.795 $Y2=3.075
r325 31 57 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.02 $Y=3.15 $X2=5.93
+ $Y2=3.15
r326 30 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.72 $Y=3.15
+ $X2=8.795 $Y2=3.075
r327 30 31 1384.47 $w=1.5e-07 $l=2.7e-06 $layer=POLY_cond $X=8.72 $Y=3.15
+ $X2=6.02 $Y2=3.15
r328 27 29 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.93 $Y=2.81
+ $X2=5.93 $Y2=2.525
r329 26 57 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.93 $Y=3.075
+ $X2=5.93 $Y2=3.15
r330 25 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.93 $Y=2.9 $X2=5.93
+ $Y2=2.81
r331 25 26 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=5.93 $Y=2.9
+ $X2=5.93 $Y2=3.075
r332 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.27 $Y=0.9 $X2=5.27
+ $Y2=0.615
r333 20 57 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.84 $Y=3.15 $X2=5.93
+ $Y2=3.15
r334 20 21 469.181 $w=1.5e-07 $l=9.15e-07 $layer=POLY_cond $X=5.84 $Y=3.15
+ $X2=4.925 $Y2=3.15
r335 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.195 $Y=0.975
+ $X2=5.27 $Y2=0.9
r336 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.195 $Y=0.975
+ $X2=4.925 $Y2=0.975
r337 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.85 $Y=3.075
+ $X2=4.925 $Y2=3.15
r338 16 56 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.85 $Y=1.68
+ $X2=4.85 $Y2=1.515
r339 16 17 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=4.85 $Y=1.68
+ $X2=4.85 $Y2=3.075
r340 15 56 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.85 $Y=1.35
+ $X2=4.85 $Y2=1.515
r341 14 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.85 $Y=1.05
+ $X2=4.925 $Y2=0.975
r342 14 15 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=4.85 $Y=1.05 $X2=4.85
+ $Y2=1.35
r343 11 54 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.295 $Y=1.765
+ $X2=4.295 $Y2=1.557
r344 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.295 $Y=1.765
+ $X2=4.295 $Y2=2.4
r345 7 54 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=4.28 $Y=1.35
+ $X2=4.295 $Y2=1.557
r346 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.28 $Y=1.35 $X2=4.28
+ $Y2=0.74
r347 2 82 600 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=1.84 $X2=3.24 $Y2=2.02
r348 1 63 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.42
+ $Y=0.37 $X2=3.565 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%A_2513_258# 1 2 8 9 11 14 18 19 22 23 25 26
+ 29 32 33 37
c103 8 0 1.21745e-19 $X=12.8 $Y=2.375
r104 35 37 5.22619 $w=4.28e-07 $l=1.95e-07 $layer=LI1_cond $X=14.035 $Y=2.695
+ $X2=14.23 $Y2=2.695
r105 32 37 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=14.23 $Y=2.48
+ $X2=14.23 $Y2=2.695
r106 31 33 3.70735 $w=2.5e-07 $l=2.26548e-07 $layer=LI1_cond $X=14.23 $Y=1.13
+ $X2=14.042 $Y2=1.045
r107 31 32 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=14.23 $Y=1.13
+ $X2=14.23 $Y2=2.48
r108 27 33 3.70735 $w=2.5e-07 $l=1.43332e-07 $layer=LI1_cond $X=13.935 $Y=0.96
+ $X2=14.042 $Y2=1.045
r109 27 29 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=13.935 $Y=0.96
+ $X2=13.935 $Y2=0.58
r110 25 33 2.76166 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=13.77 $Y=1.045
+ $X2=14.042 $Y2=1.045
r111 25 26 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=13.77 $Y=1.045
+ $X2=12.895 $Y2=1.045
r112 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.73
+ $Y=1.455 $X2=12.73 $Y2=1.455
r113 20 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.73 $Y=1.13
+ $X2=12.895 $Y2=1.045
r114 20 22 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=12.73 $Y=1.13
+ $X2=12.73 $Y2=1.455
r115 18 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=12.73 $Y=1.795
+ $X2=12.73 $Y2=1.455
r116 18 19 39.9504 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.73 $Y=1.795
+ $X2=12.73 $Y2=1.96
r117 17 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.73 $Y=1.29
+ $X2=12.73 $Y2=1.455
r118 14 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=12.82 $Y=0.58
+ $X2=12.82 $Y2=1.29
r119 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.8 $Y=2.465
+ $X2=12.8 $Y2=2.75
r120 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.8 $Y=2.375 $X2=12.8
+ $Y2=2.465
r121 8 19 161.315 $w=1.8e-07 $l=4.15e-07 $layer=POLY_cond $X=12.8 $Y=2.375
+ $X2=12.8 $Y2=1.96
r122 2 35 600 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=1 $X=13.89
+ $Y=2.47 $X2=14.035 $Y2=2.695
r123 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=13.795
+ $Y=0.37 $X2=13.935 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%A_2067_74# 1 2 3 4 5 18 20 22 23 24 26 29
+ 32 33 35 36 40 43 44 46 47 50 51 53 56 59 61 63 64 65 68 70 71 72 74 75 80 84
+ 88 90 92 93 96 104 105
c240 104 0 1.95075e-19 $X=12.105 $Y=2.125
c241 70 0 1.00509e-19 $X=11.82 $Y=2.125
r242 106 107 2.86159 $w=5.68e-07 $l=8.5e-08 $layer=LI1_cond $X=12.105 $Y=2.225
+ $X2=12.105 $Y2=2.31
r243 104 106 2.09838 $w=5.68e-07 $l=1e-07 $layer=LI1_cond $X=12.105 $Y=2.125
+ $X2=12.105 $Y2=2.225
r244 104 105 8.28231 $w=5.68e-07 $l=8.5e-08 $layer=LI1_cond $X=12.105 $Y=2.125
+ $X2=12.105 $Y2=2.04
r245 96 98 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=10.545 $Y=0.81
+ $X2=10.545 $Y2=0.945
r246 93 111 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=13.81 $Y=1.465
+ $X2=13.81 $Y2=2.145
r247 92 93 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=13.81
+ $Y=1.465 $X2=13.81 $Y2=1.465
r248 90 111 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=13.81
+ $Y=2.145 $X2=13.81 $Y2=2.145
r249 90 92 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=13.81 $Y=2.14
+ $X2=13.81 $Y2=1.465
r250 86 90 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.475 $Y=2.225
+ $X2=13.81 $Y2=2.225
r251 86 88 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=13.475 $Y=2.31
+ $X2=13.475 $Y2=2.75
r252 85 106 7.98728 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=12.39 $Y=2.225
+ $X2=12.105 $Y2=2.225
r253 84 86 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=13.31 $Y=2.225
+ $X2=13.475 $Y2=2.225
r254 84 85 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=13.31 $Y=2.225
+ $X2=12.39 $Y2=2.225
r255 82 105 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=12.305 $Y=0.73
+ $X2=12.305 $Y2=2.04
r256 80 107 5.04194 $w=3.98e-07 $l=1.75e-07 $layer=LI1_cond $X=12.02 $Y=2.485
+ $X2=12.02 $Y2=2.31
r257 75 102 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=11.465 $Y=0.565
+ $X2=11.465 $Y2=0.945
r258 75 77 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=11.55 $Y=0.565
+ $X2=12.215 $Y2=0.565
r259 74 82 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.22 $Y=0.565
+ $X2=12.305 $Y2=0.73
r260 74 77 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=12.22 $Y=0.565
+ $X2=12.215 $Y2=0.565
r261 73 98 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.71 $Y=0.945
+ $X2=10.545 $Y2=0.945
r262 72 102 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.38 $Y=0.945
+ $X2=11.465 $Y2=0.945
r263 72 73 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.38 $Y=0.945
+ $X2=10.71 $Y2=0.945
r264 70 104 7.98728 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=11.82 $Y=2.125
+ $X2=12.105 $Y2=2.125
r265 70 71 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=11.82 $Y=2.125
+ $X2=10.575 $Y2=2.125
r266 66 71 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.45 $Y=2.21
+ $X2=10.575 $Y2=2.125
r267 66 68 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=10.45 $Y=2.21
+ $X2=10.45 $Y2=2.46
r268 60 111 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=13.81 $Y=2.16
+ $X2=13.81 $Y2=2.145
r269 58 93 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=13.81 $Y=1.45
+ $X2=13.81 $Y2=1.465
r270 58 59 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=13.81 $Y=1.45
+ $X2=13.81 $Y2=1.375
r271 54 65 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=16.27 $Y=1.3
+ $X2=16.255 $Y2=1.375
r272 54 56 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=16.27 $Y=1.3
+ $X2=16.27 $Y2=0.79
r273 51 53 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=16.255 $Y=1.765
+ $X2=16.255 $Y2=2.34
r274 50 51 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=16.255 $Y=1.675
+ $X2=16.255 $Y2=1.765
r275 49 65 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=16.255 $Y=1.45
+ $X2=16.255 $Y2=1.375
r276 49 50 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=16.255 $Y=1.45
+ $X2=16.255 $Y2=1.675
r277 48 64 13.2179 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=15.335 $Y=1.375
+ $X2=15.245 $Y2=1.375
r278 47 65 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=16.165 $Y=1.375
+ $X2=16.255 $Y2=1.375
r279 47 48 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=16.165 $Y=1.375
+ $X2=15.335 $Y2=1.375
r280 44 46 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=15.245 $Y=1.765
+ $X2=15.245 $Y2=2.4
r281 43 44 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=15.245 $Y=1.675
+ $X2=15.245 $Y2=1.765
r282 42 64 10.9219 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=15.245 $Y=1.45
+ $X2=15.245 $Y2=1.375
r283 42 43 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=15.245 $Y=1.45
+ $X2=15.245 $Y2=1.675
r284 38 64 10.9219 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=15.23 $Y=1.3
+ $X2=15.245 $Y2=1.375
r285 38 40 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=15.23 $Y=1.3
+ $X2=15.23 $Y2=0.74
r286 37 63 13.2179 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=14.885 $Y=1.375
+ $X2=14.795 $Y2=1.375
r287 36 64 13.2179 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=15.155 $Y=1.375
+ $X2=15.245 $Y2=1.375
r288 36 37 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=15.155 $Y=1.375
+ $X2=14.885 $Y2=1.375
r289 33 35 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=14.795 $Y=1.765
+ $X2=14.795 $Y2=2.4
r290 32 33 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=14.795 $Y=1.675
+ $X2=14.795 $Y2=1.765
r291 31 63 10.9219 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=14.795 $Y=1.45
+ $X2=14.795 $Y2=1.375
r292 31 32 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=14.795 $Y=1.45
+ $X2=14.795 $Y2=1.675
r293 27 63 10.9219 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=14.78 $Y=1.3
+ $X2=14.795 $Y2=1.375
r294 27 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=14.78 $Y=1.3
+ $X2=14.78 $Y2=0.74
r295 24 61 64.3434 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=14.26 $Y=2.395
+ $X2=14.26 $Y2=2.235
r296 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=14.26 $Y=2.395
+ $X2=14.26 $Y2=2.68
r297 23 60 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=13.975 $Y=2.235
+ $X2=13.81 $Y2=2.16
r298 22 61 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=14.17 $Y=2.235
+ $X2=14.26 $Y2=2.235
r299 22 23 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=14.17 $Y=2.235
+ $X2=13.975 $Y2=2.235
r300 21 59 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.975 $Y=1.375
+ $X2=13.81 $Y2=1.375
r301 20 63 13.2179 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=14.705 $Y=1.375
+ $X2=14.795 $Y2=1.375
r302 20 21 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=14.705 $Y=1.375
+ $X2=13.975 $Y2=1.375
r303 16 59 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=13.72 $Y=1.3
+ $X2=13.81 $Y2=1.375
r304 16 18 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=13.72 $Y=1.3
+ $X2=13.72 $Y2=0.58
r305 5 88 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=13.325
+ $Y=2.54 $X2=13.475 $Y2=2.75
r306 4 80 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=11.835
+ $Y=2.275 $X2=11.985 $Y2=2.485
r307 3 68 600 $w=1.7e-07 $l=4.08167e-07 $layer=licon1_PDIFF $count=1 $X=10.34
+ $Y=2.12 $X2=10.49 $Y2=2.46
r308 2 77 91 $w=1.7e-07 $l=8.46906e-07 $layer=licon1_NDIFF $count=2 $X=11.46
+ $Y=0.37 $X2=12.215 $Y2=0.565
r309 1 96 182 $w=1.7e-07 $l=5.3479e-07 $layer=licon1_NDIFF $count=1 $X=10.335
+ $Y=0.37 $X2=10.545 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%A_3177_368# 1 2 7 9 12 14 16 19 23 27 33 36
+ 40
c69 7 0 1.00299e-19 $X=16.805 $Y=1.765
r70 40 41 1.2359 $w=3.9e-07 $l=1e-08 $layer=POLY_cond $X=17.255 $Y=1.532
+ $X2=17.265 $Y2=1.532
r71 39 40 51.9077 $w=3.9e-07 $l=4.2e-07 $layer=POLY_cond $X=16.835 $Y=1.532
+ $X2=17.255 $Y2=1.532
r72 38 39 3.70769 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=16.805 $Y=1.532
+ $X2=16.835 $Y2=1.532
r73 34 38 10.5051 $w=3.9e-07 $l=8.5e-08 $layer=POLY_cond $X=16.72 $Y=1.532
+ $X2=16.805 $Y2=1.532
r74 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.72
+ $Y=1.465 $X2=16.72 $Y2=1.465
r75 31 36 1.47678 $w=3.3e-07 $l=1.78e-07 $layer=LI1_cond $X=16.22 $Y=1.465
+ $X2=16.042 $Y2=1.465
r76 31 33 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=16.22 $Y=1.465
+ $X2=16.72 $Y2=1.465
r77 27 29 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=16.03 $Y=1.985
+ $X2=16.03 $Y2=2.695
r78 25 36 5.00808 $w=3.42e-07 $l=1.70895e-07 $layer=LI1_cond $X=16.03 $Y=1.63
+ $X2=16.042 $Y2=1.465
r79 25 27 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=16.03 $Y=1.63
+ $X2=16.03 $Y2=1.985
r80 21 36 5.00808 $w=3.42e-07 $l=1.65e-07 $layer=LI1_cond $X=16.042 $Y=1.3
+ $X2=16.042 $Y2=1.465
r81 21 23 22.2373 $w=3.53e-07 $l=6.85e-07 $layer=LI1_cond $X=16.042 $Y=1.3
+ $X2=16.042 $Y2=0.615
r82 17 41 25.2441 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=17.265 $Y=1.3
+ $X2=17.265 $Y2=1.532
r83 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=17.265 $Y=1.3
+ $X2=17.265 $Y2=0.74
r84 14 40 25.2441 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=17.255 $Y=1.765
+ $X2=17.255 $Y2=1.532
r85 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=17.255 $Y=1.765
+ $X2=17.255 $Y2=2.4
r86 10 39 25.2441 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=16.835 $Y=1.3
+ $X2=16.835 $Y2=1.532
r87 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=16.835 $Y=1.3
+ $X2=16.835 $Y2=0.74
r88 7 38 25.2441 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=16.805 $Y=1.765
+ $X2=16.805 $Y2=1.532
r89 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=16.805 $Y=1.765
+ $X2=16.805 $Y2=2.4
r90 2 29 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=15.885
+ $Y=1.84 $X2=16.03 $Y2=2.695
r91 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=15.885
+ $Y=1.84 $X2=16.03 $Y2=1.985
r92 1 23 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=15.91
+ $Y=0.47 $X2=16.055 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%VPWR 1 2 3 4 5 6 7 8 9 10 11 36 40 46 48 52
+ 56 60 64 70 76 80 82 87 88 90 91 93 94 96 97 98 100 105 113 137 141 147 150
+ 155 161 163 168 171 175
c200 161 0 9.36703e-20 $X=4.22 $Y=3.032
c201 52 0 6.75068e-20 $X=8.5 $Y=2.57
r202 174 175 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.52 $Y=3.33
+ $X2=17.52 $Y2=3.33
r203 171 172 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.56 $Y=3.33
+ $X2=16.56 $Y2=3.33
r204 168 169 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r205 164 169 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r206 164 166 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r207 163 166 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r208 163 164 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r209 159 161 10.8262 $w=7.63e-07 $l=1.4e-07 $layer=LI1_cond $X=4.08 $Y=3.032
+ $X2=4.22 $Y2=3.032
r210 159 160 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r211 157 159 0.390875 $w=7.63e-07 $l=2.5e-08 $layer=LI1_cond $X=4.055 $Y=3.032
+ $X2=4.08 $Y2=3.032
r212 154 160 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r213 153 157 7.11393 $w=7.63e-07 $l=4.55e-07 $layer=LI1_cond $X=3.6 $Y=3.032
+ $X2=4.055 $Y2=3.032
r214 153 155 9.80992 $w=7.63e-07 $l=7.5e-08 $layer=LI1_cond $X=3.6 $Y=3.032
+ $X2=3.525 $Y2=3.032
r215 153 154 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r216 151 154 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r217 150 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r218 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r219 145 175 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.04 $Y=3.33
+ $X2=17.52 $Y2=3.33
r220 145 172 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.04 $Y=3.33
+ $X2=16.56 $Y2=3.33
r221 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=3.33
+ $X2=17.04 $Y2=3.33
r222 142 171 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.665 $Y=3.33
+ $X2=16.54 $Y2=3.33
r223 142 144 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=16.665 $Y=3.33
+ $X2=17.04 $Y2=3.33
r224 141 174 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=17.395 $Y=3.33
+ $X2=17.577 $Y2=3.33
r225 141 144 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=17.395 $Y=3.33
+ $X2=17.04 $Y2=3.33
r226 140 172 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.08 $Y=3.33
+ $X2=16.56 $Y2=3.33
r227 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.08 $Y=3.33
+ $X2=16.08 $Y2=3.33
r228 137 171 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.415 $Y=3.33
+ $X2=16.54 $Y2=3.33
r229 137 139 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=16.415 $Y=3.33
+ $X2=16.08 $Y2=3.33
r230 136 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=16.08 $Y2=3.33
r231 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r232 133 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=15.12 $Y2=3.33
r233 132 133 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r234 130 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=14.16 $Y2=3.33
r235 129 132 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=13.2 $Y=3.33
+ $X2=14.16 $Y2=3.33
r236 129 130 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r237 127 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r238 126 127 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=12.72
+ $Y=3.33 $X2=12.72 $Y2=3.33
r239 124 127 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=12.72 $Y2=3.33
r240 123 126 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=9.84 $Y=3.33
+ $X2=12.72 $Y2=3.33
r241 123 124 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r242 121 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r243 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r244 118 168 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.665 $Y=3.33
+ $X2=8.5 $Y2=3.33
r245 118 120 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=8.665 $Y=3.33
+ $X2=9.36 $Y2=3.33
r246 117 166 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r247 117 160 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r248 116 161 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=4.22 $Y2=3.33
r249 116 117 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r250 113 163 12.2593 $w=1.7e-07 $l=2.87e-07 $layer=LI1_cond $X=6.41 $Y=3.33
+ $X2=6.697 $Y2=3.33
r251 113 116 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=6.41 $Y=3.33
+ $X2=4.56 $Y2=3.33
r252 112 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r253 111 112 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r254 109 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r255 109 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r256 108 111 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r257 108 109 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r258 106 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=0.8 $Y2=3.33
r259 106 108 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=1.2 $Y2=3.33
r260 105 150 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.495 $Y=3.33
+ $X2=2.67 $Y2=3.33
r261 105 111 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.495 $Y=3.33
+ $X2=2.16 $Y2=3.33
r262 103 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r263 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r264 100 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.8 $Y2=3.33
r265 100 102 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r266 98 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r267 98 169 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r268 96 135 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=15.305 $Y=3.33
+ $X2=15.12 $Y2=3.33
r269 96 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.305 $Y=3.33
+ $X2=15.47 $Y2=3.33
r270 95 139 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=15.635 $Y=3.33
+ $X2=16.08 $Y2=3.33
r271 95 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.635 $Y=3.33
+ $X2=15.47 $Y2=3.33
r272 93 132 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=14.485 $Y=3.33
+ $X2=14.16 $Y2=3.33
r273 93 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.485 $Y=3.33
+ $X2=14.57 $Y2=3.33
r274 92 135 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=14.655 $Y=3.33
+ $X2=15.12 $Y2=3.33
r275 92 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.655 $Y=3.33
+ $X2=14.57 $Y2=3.33
r276 90 126 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=12.94 $Y=3.33
+ $X2=12.72 $Y2=3.33
r277 90 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.94 $Y=3.33
+ $X2=13.025 $Y2=3.33
r278 89 129 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=13.11 $Y=3.33
+ $X2=13.2 $Y2=3.33
r279 89 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.11 $Y=3.33
+ $X2=13.025 $Y2=3.33
r280 87 120 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=9.425 $Y=3.33
+ $X2=9.36 $Y2=3.33
r281 87 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.425 $Y=3.33
+ $X2=9.55 $Y2=3.33
r282 86 123 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.675 $Y=3.33
+ $X2=9.84 $Y2=3.33
r283 86 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.675 $Y=3.33
+ $X2=9.55 $Y2=3.33
r284 82 85 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=17.52 $Y=1.985
+ $X2=17.52 $Y2=2.815
r285 80 174 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=17.52 $Y=3.245
+ $X2=17.577 $Y2=3.33
r286 80 85 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=17.52 $Y=3.245
+ $X2=17.52 $Y2=2.815
r287 76 79 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=16.54 $Y=1.985
+ $X2=16.54 $Y2=2.815
r288 74 171 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.54 $Y=3.245
+ $X2=16.54 $Y2=3.33
r289 74 79 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=16.54 $Y=3.245
+ $X2=16.54 $Y2=2.815
r290 70 73 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=15.47 $Y=1.985
+ $X2=15.47 $Y2=2.815
r291 68 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.47 $Y=3.245
+ $X2=15.47 $Y2=3.33
r292 68 73 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=15.47 $Y=3.245
+ $X2=15.47 $Y2=2.815
r293 64 67 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=14.57 $Y=1.985
+ $X2=14.57 $Y2=2.815
r294 62 94 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.57 $Y=3.245
+ $X2=14.57 $Y2=3.33
r295 62 67 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=14.57 $Y=3.245
+ $X2=14.57 $Y2=2.815
r296 58 91 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.025 $Y=3.245
+ $X2=13.025 $Y2=3.33
r297 58 60 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=13.025 $Y=3.245
+ $X2=13.025 $Y2=2.75
r298 54 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.55 $Y=3.245
+ $X2=9.55 $Y2=3.33
r299 54 56 23.9708 $w=2.48e-07 $l=5.2e-07 $layer=LI1_cond $X=9.55 $Y=3.245
+ $X2=9.55 $Y2=2.725
r300 50 168 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.5 $Y=3.245
+ $X2=8.5 $Y2=3.33
r301 50 52 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=8.5 $Y=3.245
+ $X2=8.5 $Y2=2.57
r302 49 163 12.2593 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=6.985 $Y=3.33
+ $X2=6.697 $Y2=3.33
r303 48 168 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.335 $Y=3.33
+ $X2=8.5 $Y2=3.33
r304 48 49 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=8.335 $Y=3.33
+ $X2=6.985 $Y2=3.33
r305 44 163 2.42056 $w=5.75e-07 $l=8.5e-08 $layer=LI1_cond $X=6.697 $Y=3.245
+ $X2=6.697 $Y2=3.33
r306 44 46 13.6249 $w=5.73e-07 $l=6.55e-07 $layer=LI1_cond $X=6.697 $Y=3.245
+ $X2=6.697 $Y2=2.59
r307 43 150 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=2.67 $Y2=3.33
r308 43 155 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=3.525 $Y2=3.33
r309 38 150 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=3.245
+ $X2=2.67 $Y2=3.33
r310 38 40 14.1586 $w=3.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.67 $Y=3.245
+ $X2=2.67 $Y2=2.815
r311 34 147 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=3.245
+ $X2=0.8 $Y2=3.33
r312 34 36 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.8 $Y=3.245
+ $X2=0.8 $Y2=2.475
r313 11 85 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=17.33
+ $Y=1.84 $X2=17.48 $Y2=2.815
r314 11 82 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=17.33
+ $Y=1.84 $X2=17.48 $Y2=1.985
r315 10 79 600 $w=1.7e-07 $l=1.09287e-06 $layer=licon1_PDIFF $count=1 $X=16.33
+ $Y=1.84 $X2=16.58 $Y2=2.815
r316 10 76 300 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_PDIFF $count=2 $X=16.33
+ $Y=1.84 $X2=16.58 $Y2=1.985
r317 9 73 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=15.32
+ $Y=1.84 $X2=15.47 $Y2=2.815
r318 9 70 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=15.32
+ $Y=1.84 $X2=15.47 $Y2=1.985
r319 8 67 400 $w=1.7e-07 $l=4.47325e-07 $layer=licon1_PDIFF $count=1 $X=14.335
+ $Y=2.47 $X2=14.57 $Y2=2.815
r320 8 64 400 $w=1.7e-07 $l=5.90931e-07 $layer=licon1_PDIFF $count=1 $X=14.335
+ $Y=2.47 $X2=14.57 $Y2=1.985
r321 7 60 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=12.875
+ $Y=2.54 $X2=13.025 $Y2=2.75
r322 6 56 600 $w=1.7e-07 $l=6.75851e-07 $layer=licon1_PDIFF $count=1 $X=9.44
+ $Y=2.12 $X2=9.59 $Y2=2.725
r323 5 52 600 $w=1.7e-07 $l=5.52992e-07 $layer=licon1_PDIFF $count=1 $X=8.06
+ $Y=2.315 $X2=8.5 $Y2=2.57
r324 4 46 600 $w=1.7e-07 $l=3.87137e-07 $layer=licon1_PDIFF $count=1 $X=6.425
+ $Y=2.315 $X2=6.695 $Y2=2.59
r325 3 157 300 $w=1.7e-07 $l=1.2053e-06 $layer=licon1_PDIFF $count=2 $X=3.54
+ $Y=1.84 $X2=4.055 $Y2=2.815
r326 2 40 600 $w=1.7e-07 $l=5.69408e-07 $layer=licon1_PDIFF $count=1 $X=2.51
+ $Y=2.32 $X2=2.67 $Y2=2.815
r327 1 36 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=2.32 $X2=0.8 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%A_304_464# 1 2 3 4 15 18 19 21 26 28 30 31
+ 36 39 40
c113 40 0 9.15331e-20 $X=5.13 $Y=2.13
c114 21 0 9.54145e-20 $X=4.89 $Y=2.215
r115 39 42 7.47549 $w=4.78e-07 $l=3e-07 $layer=LI1_cond $X=5.13 $Y=2.215
+ $X2=5.13 $Y2=2.515
r116 39 40 7.40287 $w=4.78e-07 $l=8.5e-08 $layer=LI1_cond $X=5.13 $Y=2.215
+ $X2=5.13 $Y2=2.13
r117 38 40 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=4.975 $Y=0.845
+ $X2=4.975 $Y2=2.13
r118 36 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.055 $Y=0.68
+ $X2=5.055 $Y2=0.845
r119 31 33 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.8 $Y=2.215
+ $X2=3.8 $Y2=2.395
r120 28 29 18.4636 $w=2.61e-07 $l=3.95e-07 $layer=LI1_cond $X=2.155 $Y=0.565
+ $X2=2.55 $Y2=0.565
r121 22 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.885 $Y=2.215
+ $X2=3.8 $Y2=2.215
r122 21 39 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=4.89 $Y=2.215
+ $X2=5.13 $Y2=2.215
r123 21 22 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=4.89 $Y=2.215
+ $X2=3.885 $Y2=2.215
r124 20 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=2.395
+ $X2=2.55 $Y2=2.395
r125 19 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.715 $Y=2.395
+ $X2=3.8 $Y2=2.395
r126 19 20 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=3.715 $Y=2.395
+ $X2=2.635 $Y2=2.395
r127 18 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=2.31
+ $X2=2.55 $Y2=2.395
r128 17 29 3.24614 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=0.73
+ $X2=2.55 $Y2=0.565
r129 17 18 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=2.55 $Y=0.73
+ $X2=2.55 $Y2=2.31
r130 16 26 6.39056 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=1.955 $Y=2.395
+ $X2=1.73 $Y2=2.395
r131 15 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=2.395
+ $X2=2.55 $Y2=2.395
r132 15 16 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.465 $Y=2.395
+ $X2=1.955 $Y2=2.395
r133 4 42 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=5.06
+ $Y=2.315 $X2=5.205 $Y2=2.515
r134 3 26 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=1.52
+ $Y=2.32 $X2=1.73 $Y2=2.465
r135 2 36 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=4.91
+ $Y=0.405 $X2=5.055 $Y2=0.68
r136 1 28 182 $w=1.7e-07 $l=7.10845e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.37 $X2=2.155 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%A_1789_424# 1 2 3 12 14 15 16 17 20 23
c54 17 0 1.20006e-19 $X=10.125 $Y=2.99
c55 14 0 1.43203e-19 $X=10 $Y=2.3
r56 18 20 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=10.94 $Y=2.905
+ $X2=10.94 $Y2=2.465
r57 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.775 $Y=2.99
+ $X2=10.94 $Y2=2.905
r58 16 17 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=10.775 $Y=2.99
+ $X2=10.125 $Y2=2.99
r59 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10 $Y=2.905
+ $X2=10.125 $Y2=2.99
r60 14 25 2.97632 $w=2.5e-07 $l=1e-07 $layer=LI1_cond $X=10 $Y=2.3 $X2=10
+ $Y2=2.2
r61 14 15 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=10 $Y=2.3 $X2=10
+ $Y2=2.905
r62 13 23 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.255 $Y=2.215
+ $X2=9.09 $Y2=2.215
r63 12 25 4.16685 $w=1.7e-07 $l=1.32288e-07 $layer=LI1_cond $X=9.875 $Y=2.215
+ $X2=10 $Y2=2.2
r64 12 13 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=9.875 $Y=2.215
+ $X2=9.255 $Y2=2.215
r65 3 20 300 $w=1.7e-07 $l=4.13249e-07 $layer=licon1_PDIFF $count=2 $X=10.79
+ $Y=2.12 $X2=10.94 $Y2=2.465
r66 2 25 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=9.89
+ $Y=2.12 $X2=10.04 $Y2=2.265
r67 1 23 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=8.945
+ $Y=2.12 $X2=9.09 $Y2=2.295
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%A_2277_455# 1 2 9 11 12 15
r32 13 15 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=12.575 $Y=2.885
+ $X2=12.575 $Y2=2.75
r33 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.41 $Y=2.97
+ $X2=12.575 $Y2=2.885
r34 11 12 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=12.41 $Y=2.97
+ $X2=11.62 $Y2=2.97
r35 7 12 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=11.492 $Y=2.885
+ $X2=11.62 $Y2=2.97
r36 7 9 15.1399 $w=2.53e-07 $l=3.35e-07 $layer=LI1_cond $X=11.492 $Y=2.885
+ $X2=11.492 $Y2=2.55
r37 2 15 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=12.43
+ $Y=2.54 $X2=12.575 $Y2=2.75
r38 1 9 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=11.385
+ $Y=2.275 $X2=11.53 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%Q_N 1 2 9 13 14 15 22 30
r28 20 30 2.30489 $w=3.83e-07 $l=7.7e-08 $layer=LI1_cond $X=15.042 $Y=1.218
+ $X2=15.042 $Y2=1.295
r29 15 32 4.63829 $w=3.83e-07 $l=1.11e-07 $layer=LI1_cond $X=15.042 $Y=1.299
+ $X2=15.042 $Y2=1.41
r30 15 30 0.119734 $w=3.83e-07 $l=4e-09 $layer=LI1_cond $X=15.042 $Y=1.299
+ $X2=15.042 $Y2=1.295
r31 15 20 0.119734 $w=3.83e-07 $l=4e-09 $layer=LI1_cond $X=15.042 $Y=1.214
+ $X2=15.042 $Y2=1.218
r32 14 15 8.65081 $w=3.83e-07 $l=2.89e-07 $layer=LI1_cond $X=15.042 $Y=0.925
+ $X2=15.042 $Y2=1.214
r33 13 14 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=15.042 $Y=0.555
+ $X2=15.042 $Y2=0.925
r34 13 22 1.19734 $w=3.83e-07 $l=4e-08 $layer=LI1_cond $X=15.042 $Y=0.555
+ $X2=15.042 $Y2=0.515
r35 9 11 37.5109 $w=2.53e-07 $l=8.3e-07 $layer=LI1_cond $X=14.977 $Y=1.985
+ $X2=14.977 $Y2=2.815
r36 9 32 25.9865 $w=2.53e-07 $l=5.75e-07 $layer=LI1_cond $X=14.977 $Y=1.985
+ $X2=14.977 $Y2=1.41
r37 2 11 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=14.87
+ $Y=1.84 $X2=15.02 $Y2=2.815
r38 2 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=14.87
+ $Y=1.84 $X2=15.02 $Y2=1.985
r39 1 22 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=14.855
+ $Y=0.37 $X2=15.015 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%Q 1 2 9 14 15 16 17 28
c30 15 0 1.00299e-19 $X=17.045 $Y=1.82
r31 21 28 1.18634 $w=3.38e-07 $l=3.5e-08 $layer=LI1_cond $X=17.055 $Y=0.96
+ $X2=17.055 $Y2=0.925
r32 17 30 7.79401 $w=3.38e-07 $l=1.45e-07 $layer=LI1_cond $X=17.055 $Y=0.985
+ $X2=17.055 $Y2=1.13
r33 17 21 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=17.055 $Y=0.985
+ $X2=17.055 $Y2=0.96
r34 17 28 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=17.055 $Y=0.9
+ $X2=17.055 $Y2=0.925
r35 16 17 13.0497 $w=3.38e-07 $l=3.85e-07 $layer=LI1_cond $X=17.055 $Y=0.515
+ $X2=17.055 $Y2=0.9
r36 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=17.14 $Y=1.82
+ $X2=17.14 $Y2=1.13
r37 14 15 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=17.045 $Y=1.985
+ $X2=17.045 $Y2=1.82
r38 7 14 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=17.045 $Y=2
+ $X2=17.045 $Y2=1.985
r39 7 9 26.09 $w=3.58e-07 $l=8.15e-07 $layer=LI1_cond $X=17.045 $Y=2 $X2=17.045
+ $Y2=2.815
r40 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=16.88
+ $Y=1.84 $X2=17.03 $Y2=1.985
r41 2 9 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=16.88
+ $Y=1.84 $X2=17.03 $Y2=2.815
r42 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=16.91
+ $Y=0.37 $X2=17.05 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%VGND 1 2 3 4 5 6 7 8 9 10 11 36 40 44 48 52
+ 56 60 64 68 72 74 76 79 80 82 83 85 86 88 89 91 92 93 95 107 111 116 137 141
+ 147 150 153 156 159 163
r183 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.52 $Y=0
+ $X2=17.52 $Y2=0
r184 159 160 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.56 $Y=0
+ $X2=16.56 $Y2=0
r185 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r186 153 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r187 150 151 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r188 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r189 145 163 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.04 $Y=0
+ $X2=17.52 $Y2=0
r190 145 160 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.04 $Y=0
+ $X2=16.56 $Y2=0
r191 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=0
+ $X2=17.04 $Y2=0
r192 142 159 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.705 $Y=0
+ $X2=16.58 $Y2=0
r193 142 144 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=16.705 $Y=0
+ $X2=17.04 $Y2=0
r194 141 162 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=17.395 $Y=0
+ $X2=17.577 $Y2=0
r195 141 144 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=17.395 $Y=0
+ $X2=17.04 $Y2=0
r196 140 160 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.08 $Y=0
+ $X2=16.56 $Y2=0
r197 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.08 $Y=0
+ $X2=16.08 $Y2=0
r198 137 159 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.455 $Y=0
+ $X2=16.58 $Y2=0
r199 137 139 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=16.455 $Y=0
+ $X2=16.08 $Y2=0
r200 136 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=16.08 $Y2=0
r201 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r202 133 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=15.12 $Y2=0
r203 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r204 130 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=14.16 $Y2=0
r205 129 130 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r206 127 130 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=13.2 $Y2=0
r207 126 129 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=9.84 $Y=0
+ $X2=13.2 $Y2=0
r208 126 127 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r209 124 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r210 123 124 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r211 121 156 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.53 $Y=0
+ $X2=8.365 $Y2=0
r212 121 123 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=8.53 $Y=0
+ $X2=9.36 $Y2=0
r213 120 157 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.4 $Y2=0
r214 120 154 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=6.96 $Y2=0
r215 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r216 117 153 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=7.15 $Y=0
+ $X2=6.982 $Y2=0
r217 117 119 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=7.15 $Y=0
+ $X2=7.92 $Y2=0
r218 116 156 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.2 $Y=0
+ $X2=8.365 $Y2=0
r219 116 119 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=8.2 $Y=0 $X2=7.92
+ $Y2=0
r220 115 154 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r221 115 151 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=4.08 $Y2=0
r222 114 115 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r223 112 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.16 $Y=0
+ $X2=3.995 $Y2=0
r224 112 114 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=4.16 $Y=0
+ $X2=6.48 $Y2=0
r225 111 153 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=6.815 $Y=0
+ $X2=6.982 $Y2=0
r226 111 114 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.815 $Y=0
+ $X2=6.48 $Y2=0
r227 110 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=4.08 $Y2=0
r228 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r229 107 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.83 $Y=0
+ $X2=3.995 $Y2=0
r230 107 109 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=3.6
+ $Y2=0
r231 106 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r232 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r233 103 106 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=2.64 $Y2=0
r234 103 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=0.72 $Y2=0
r235 102 105 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0
+ $X2=2.64 $Y2=0
r236 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r237 100 147 9.89127 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=1.02 $Y=0
+ $X2=0.817 $Y2=0
r238 100 102 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=1.2
+ $Y2=0
r239 98 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r240 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r241 95 147 9.89127 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.817 $Y2=0
r242 95 97 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r243 93 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r244 93 157 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r245 91 135 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=15.405 $Y=0
+ $X2=15.12 $Y2=0
r246 91 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.405 $Y=0
+ $X2=15.53 $Y2=0
r247 90 139 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=15.655 $Y=0
+ $X2=16.08 $Y2=0
r248 90 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.655 $Y=0
+ $X2=15.53 $Y2=0
r249 88 132 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=14.35 $Y=0
+ $X2=14.16 $Y2=0
r250 88 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.35 $Y=0
+ $X2=14.515 $Y2=0
r251 87 135 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=14.68 $Y=0
+ $X2=15.12 $Y2=0
r252 87 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.68 $Y=0
+ $X2=14.515 $Y2=0
r253 85 129 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=13.26 $Y=0 $X2=13.2
+ $Y2=0
r254 85 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.26 $Y=0
+ $X2=13.425 $Y2=0
r255 84 132 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=13.59 $Y=0
+ $X2=14.16 $Y2=0
r256 84 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.59 $Y=0
+ $X2=13.425 $Y2=0
r257 82 123 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=9.45 $Y=0 $X2=9.36
+ $Y2=0
r258 82 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.45 $Y=0 $X2=9.615
+ $Y2=0
r259 81 126 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=9.78 $Y=0 $X2=9.84
+ $Y2=0
r260 81 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.78 $Y=0 $X2=9.615
+ $Y2=0
r261 79 105 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.84 $Y=0 $X2=2.64
+ $Y2=0
r262 79 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.84 $Y=0 $X2=3.005
+ $Y2=0
r263 78 109 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.17 $Y=0 $X2=3.6
+ $Y2=0
r264 78 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=0 $X2=3.005
+ $Y2=0
r265 74 162 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=17.52 $Y=0.085
+ $X2=17.577 $Y2=0
r266 74 76 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=17.52 $Y=0.085
+ $X2=17.52 $Y2=0.515
r267 70 159 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.58 $Y=0.085
+ $X2=16.58 $Y2=0
r268 70 72 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=16.58 $Y=0.085
+ $X2=16.58 $Y2=0.515
r269 66 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.53 $Y=0.085
+ $X2=15.53 $Y2=0
r270 66 68 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=15.53 $Y=0.085
+ $X2=15.53 $Y2=0.515
r271 62 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.515 $Y=0.085
+ $X2=14.515 $Y2=0
r272 62 64 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=14.515 $Y=0.085
+ $X2=14.515 $Y2=0.625
r273 58 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.425 $Y=0.085
+ $X2=13.425 $Y2=0
r274 58 60 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=13.425 $Y=0.085
+ $X2=13.425 $Y2=0.57
r275 54 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.615 $Y=0.085
+ $X2=9.615 $Y2=0
r276 54 56 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=9.615 $Y=0.085
+ $X2=9.615 $Y2=0.59
r277 50 156 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.365 $Y=0.085
+ $X2=8.365 $Y2=0
r278 50 52 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.365 $Y=0.085
+ $X2=8.365 $Y2=0.515
r279 46 153 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=6.982 $Y=0.085
+ $X2=6.982 $Y2=0
r280 46 48 15.4806 $w=3.33e-07 $l=4.5e-07 $layer=LI1_cond $X=6.982 $Y=0.085
+ $X2=6.982 $Y2=0.535
r281 42 150 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=0.085
+ $X2=3.995 $Y2=0
r282 42 44 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=3.995 $Y=0.085
+ $X2=3.995 $Y2=0.505
r283 38 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.005 $Y=0.085
+ $X2=3.005 $Y2=0
r284 38 40 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.005 $Y=0.085
+ $X2=3.005 $Y2=0.565
r285 34 147 1.50354 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.817 $Y=0.085
+ $X2=0.817 $Y2=0
r286 34 36 12.2358 $w=4.03e-07 $l=4.3e-07 $layer=LI1_cond $X=0.817 $Y=0.085
+ $X2=0.817 $Y2=0.515
r287 11 76 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=17.34
+ $Y=0.37 $X2=17.48 $Y2=0.515
r288 10 72 91 $w=1.7e-07 $l=2.96648e-07 $layer=licon1_NDIFF $count=2 $X=16.345
+ $Y=0.47 $X2=16.62 $Y2=0.515
r289 9 68 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=15.305
+ $Y=0.37 $X2=15.49 $Y2=0.515
r290 8 64 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=14.37
+ $Y=0.37 $X2=14.515 $Y2=0.625
r291 7 60 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=13.285
+ $Y=0.37 $X2=13.425 $Y2=0.57
r292 6 56 182 $w=1.7e-07 $l=2.89137e-07 $layer=licon1_NDIFF $count=1 $X=9.455
+ $Y=0.37 $X2=9.615 $Y2=0.59
r293 5 52 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.225
+ $Y=0.37 $X2=8.365 $Y2=0.515
r294 4 48 182 $w=1.7e-07 $l=1.94422e-07 $layer=licon1_NDIFF $count=1 $X=6.76
+ $Y=0.405 $X2=6.9 $Y2=0.535
r295 3 44 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=3.855
+ $Y=0.37 $X2=3.995 $Y2=0.505
r296 2 40 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.37 $X2=3.005 $Y2=0.565
r297 1 36 182 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.815 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFSBP_2%A_1794_74# 1 2 3 12 14 15 19 20 21 22
c47 15 0 1.14148e-19 $X=9.28 $Y=1.09
r48 22 25 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=11.045 $Y=0.34
+ $X2=11.045 $Y2=0.52
r49 20 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.88 $Y=0.34
+ $X2=11.045 $Y2=0.34
r50 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.88 $Y=0.34
+ $X2=10.21 $Y2=0.34
r51 17 19 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=10.085 $Y=1.005
+ $X2=10.085 $Y2=0.515
r52 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.085 $Y=0.425
+ $X2=10.21 $Y2=0.34
r53 16 19 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=10.085 $Y=0.425
+ $X2=10.085 $Y2=0.515
r54 14 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.96 $Y=1.09
+ $X2=10.085 $Y2=1.005
r55 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.96 $Y=1.09
+ $X2=9.28 $Y2=1.09
r56 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.155 $Y=1.005
+ $X2=9.28 $Y2=1.09
r57 10 12 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=9.155 $Y=1.005
+ $X2=9.155 $Y2=0.515
r58 3 25 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=10.835
+ $Y=0.37 $X2=11.045 $Y2=0.52
r59 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.905
+ $Y=0.37 $X2=10.045 $Y2=0.515
r60 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=8.97
+ $Y=0.37 $X2=9.115 $Y2=0.515
.ends

