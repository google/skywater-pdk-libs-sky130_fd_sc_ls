* File: sky130_fd_sc_ls__clkbuf_8.pex.spice
* Created: Fri Aug 28 13:09:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__CLKBUF_8%A 1 3 6 10 12 14 15 16 23 24
r52 24 25 1.28533 $w=3.75e-07 $l=1e-08 $layer=POLY_cond $X=0.995 $Y=1.557
+ $X2=1.005 $Y2=1.557
r53 22 24 8.35467 $w=3.75e-07 $l=6.5e-08 $layer=POLY_cond $X=0.93 $Y=1.557
+ $X2=0.995 $Y2=1.557
r54 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.93
+ $Y=1.515 $X2=0.93 $Y2=1.515
r55 20 22 46.9147 $w=3.75e-07 $l=3.65e-07 $layer=POLY_cond $X=0.565 $Y=1.557
+ $X2=0.93 $Y2=1.557
r56 19 20 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=0.55 $Y=1.557
+ $X2=0.565 $Y2=1.557
r57 16 23 5.62821 $w=4.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.93 $Y2=1.565
r58 15 16 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.72 $Y2=1.565
r59 12 25 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=1.557
r60 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r61 8 24 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.557
r62 8 10 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.58
r63 4 20 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.565 $Y=1.35
+ $X2=0.565 $Y2=1.557
r64 4 6 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=0.565 $Y=1.35 $X2=0.565
+ $Y2=0.58
r65 1 19 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.55 $Y=1.765
+ $X2=0.55 $Y2=1.557
r66 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.55 $Y=1.765
+ $X2=0.55 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__CLKBUF_8%A_125_368# 1 2 9 12 13 15 17 20 22 24 26 27
+ 29 32 35 36 38 41 44 45 47 50 53 54 56 59 62 63 65 68 71 72 74 77 81 83 85 87
+ 88 89 92 98 103 122
r217 121 122 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.77 $Y=1.355
+ $X2=4.785 $Y2=1.355
r218 120 121 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=4.355 $Y=1.355
+ $X2=4.77 $Y2=1.355
r219 117 118 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=3.855 $Y=1.355
+ $X2=4.305 $Y2=1.355
r220 116 117 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=3.805 $Y=1.355
+ $X2=3.855 $Y2=1.355
r221 115 116 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=3.425 $Y=1.355
+ $X2=3.805 $Y2=1.355
r222 114 115 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.355 $Y=1.355
+ $X2=3.425 $Y2=1.355
r223 113 114 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.995 $Y=1.355
+ $X2=3.355 $Y2=1.355
r224 112 113 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.905 $Y=1.355
+ $X2=2.995 $Y2=1.355
r225 111 112 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.565 $Y=1.355
+ $X2=2.905 $Y2=1.355
r226 110 111 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=2.455 $Y=1.355
+ $X2=2.565 $Y2=1.355
r227 109 110 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=2.005 $Y=1.355
+ $X2=2.455 $Y2=1.355
r228 108 109 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.995 $Y=1.355
+ $X2=2.005 $Y2=1.355
r229 104 106 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.54 $Y=1.355
+ $X2=1.555 $Y2=1.355
r230 99 120 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=4.35 $Y=1.355
+ $X2=4.355 $Y2=1.355
r231 99 118 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=4.35 $Y=1.355
+ $X2=4.305 $Y2=1.355
r232 98 99 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=4.35
+ $Y=1.355 $X2=4.35 $Y2=1.355
r233 96 108 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=1.63 $Y=1.355
+ $X2=1.995 $Y2=1.355
r234 96 106 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.63 $Y=1.355
+ $X2=1.555 $Y2=1.355
r235 95 98 94.9892 $w=3.28e-07 $l=2.72e-06 $layer=LI1_cond $X=1.63 $Y=1.355
+ $X2=4.35 $Y2=1.355
r236 95 96 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=1.63
+ $Y=1.355 $X2=1.63 $Y2=1.355
r237 93 103 3.70735 $w=2.5e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.445 $Y=1.355
+ $X2=1.36 $Y2=1.25
r238 93 95 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.445 $Y=1.355
+ $X2=1.63 $Y2=1.355
r239 91 103 2.76166 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=1.36 $Y=1.52
+ $X2=1.36 $Y2=1.25
r240 91 92 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.36 $Y=1.52
+ $X2=1.36 $Y2=1.95
r241 90 102 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=2.035
+ $X2=0.78 $Y2=2.035
r242 89 92 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.275 $Y=2.035
+ $X2=1.36 $Y2=1.95
r243 89 90 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.275 $Y=2.035
+ $X2=0.945 $Y2=2.035
r244 87 103 3.70735 $w=2.5e-07 $l=2.23495e-07 $layer=LI1_cond $X=1.275 $Y=1.065
+ $X2=1.36 $Y2=1.25
r245 87 88 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.275 $Y=1.065
+ $X2=0.945 $Y2=1.065
r246 83 102 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=2.12
+ $X2=0.78 $Y2=2.035
r247 83 85 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.78 $Y=2.12
+ $X2=0.78 $Y2=2.815
r248 79 88 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=0.98
+ $X2=0.945 $Y2=1.065
r249 79 81 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=0.78 $Y=0.98 $X2=0.78
+ $Y2=0.58
r250 75 122 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.785 $Y=1.19
+ $X2=4.785 $Y2=1.355
r251 75 77 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.785 $Y=1.19
+ $X2=4.785 $Y2=0.58
r252 72 74 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.77 $Y=1.765
+ $X2=4.77 $Y2=2.4
r253 71 72 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.77 $Y=1.675
+ $X2=4.77 $Y2=1.765
r254 70 121 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.52
+ $X2=4.77 $Y2=1.355
r255 70 71 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=4.77 $Y=1.52
+ $X2=4.77 $Y2=1.675
r256 66 120 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.19
+ $X2=4.355 $Y2=1.355
r257 66 68 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.355 $Y=1.19
+ $X2=4.355 $Y2=0.58
r258 63 65 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.305 $Y=1.765
+ $X2=4.305 $Y2=2.4
r259 62 63 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.305 $Y=1.675
+ $X2=4.305 $Y2=1.765
r260 61 118 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.52
+ $X2=4.305 $Y2=1.355
r261 61 62 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=4.305 $Y=1.52
+ $X2=4.305 $Y2=1.675
r262 57 117 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.19
+ $X2=3.855 $Y2=1.355
r263 57 59 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.855 $Y=1.19
+ $X2=3.855 $Y2=0.58
r264 54 56 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.805 $Y=1.765
+ $X2=3.805 $Y2=2.4
r265 53 54 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.805 $Y=1.675
+ $X2=3.805 $Y2=1.765
r266 52 116 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.805 $Y=1.52
+ $X2=3.805 $Y2=1.355
r267 52 53 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=3.805 $Y=1.52
+ $X2=3.805 $Y2=1.675
r268 48 115 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.425 $Y=1.19
+ $X2=3.425 $Y2=1.355
r269 48 50 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.425 $Y=1.19
+ $X2=3.425 $Y2=0.58
r270 45 47 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.355 $Y=1.765
+ $X2=3.355 $Y2=2.4
r271 44 45 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.355 $Y=1.675
+ $X2=3.355 $Y2=1.765
r272 43 114 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.52
+ $X2=3.355 $Y2=1.355
r273 43 44 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=3.355 $Y=1.52
+ $X2=3.355 $Y2=1.675
r274 39 113 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.995 $Y=1.19
+ $X2=2.995 $Y2=1.355
r275 39 41 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.995 $Y=1.19
+ $X2=2.995 $Y2=0.58
r276 36 38 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.905 $Y=1.765
+ $X2=2.905 $Y2=2.4
r277 35 36 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.905 $Y=1.675
+ $X2=2.905 $Y2=1.765
r278 34 112 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.905 $Y=1.52
+ $X2=2.905 $Y2=1.355
r279 34 35 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=2.905 $Y=1.52
+ $X2=2.905 $Y2=1.675
r280 30 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.565 $Y=1.19
+ $X2=2.565 $Y2=1.355
r281 30 32 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.565 $Y=1.19
+ $X2=2.565 $Y2=0.58
r282 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.455 $Y=1.765
+ $X2=2.455 $Y2=2.4
r283 26 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.455 $Y=1.675
+ $X2=2.455 $Y2=1.765
r284 25 110 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.455 $Y=1.52
+ $X2=2.455 $Y2=1.355
r285 25 26 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=2.455 $Y=1.52
+ $X2=2.455 $Y2=1.675
r286 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.005 $Y=1.765
+ $X2=2.005 $Y2=2.4
r287 18 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.995 $Y=1.19
+ $X2=1.995 $Y2=1.355
r288 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.995 $Y=1.19
+ $X2=1.995 $Y2=0.58
r289 17 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.005 $Y=1.675
+ $X2=2.005 $Y2=1.765
r290 16 109 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.005 $Y=1.52
+ $X2=2.005 $Y2=1.355
r291 16 17 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=2.005 $Y=1.52
+ $X2=2.005 $Y2=1.675
r292 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.555 $Y=1.765
+ $X2=1.555 $Y2=2.4
r293 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.555 $Y=1.675
+ $X2=1.555 $Y2=1.765
r294 11 106 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.555 $Y=1.52
+ $X2=1.555 $Y2=1.355
r295 11 12 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=1.555 $Y=1.52
+ $X2=1.555 $Y2=1.675
r296 7 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.54 $Y=1.19
+ $X2=1.54 $Y2=1.355
r297 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.54 $Y=1.19 $X2=1.54
+ $Y2=0.58
r298 2 102 400 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_PDIFF $count=1 $X=0.625
+ $Y=1.84 $X2=0.78 $Y2=2.115
r299 2 85 400 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=0.625
+ $Y=1.84 $X2=0.78 $Y2=2.815
r300 1 81 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__CLKBUF_8%VPWR 1 2 3 4 5 6 19 21 27 31 35 39 43 47 49
+ 53 55 60 65 70 79 82 85 88 92
r85 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r86 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r87 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r88 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r89 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r90 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r91 74 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r92 74 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r93 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r94 71 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.195 $Y=3.33
+ $X2=4.03 $Y2=3.33
r95 71 73 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.195 $Y=3.33
+ $X2=4.56 $Y2=3.33
r96 70 91 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=4.83 $Y=3.33
+ $X2=5.055 $Y2=3.33
r97 70 73 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.83 $Y=3.33 $X2=4.56
+ $Y2=3.33
r98 69 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r99 69 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r100 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r101 66 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=3.33
+ $X2=3.13 $Y2=3.33
r102 66 68 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.215 $Y=3.33
+ $X2=3.6 $Y2=3.33
r103 65 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.865 $Y=3.33
+ $X2=4.03 $Y2=3.33
r104 65 68 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.865 $Y=3.33
+ $X2=3.6 $Y2=3.33
r105 64 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r106 64 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r108 61 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.28 $Y2=3.33
r109 61 63 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.68 $Y2=3.33
r110 60 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=2.23 $Y2=3.33
r111 60 63 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=1.68 $Y2=3.33
r112 59 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r113 59 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r114 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r115 56 76 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r116 56 58 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r117 55 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.28 $Y2=3.33
r118 55 58 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=0.72 $Y2=3.33
r119 53 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r120 53 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r121 49 52 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=4.995 $Y=2.115
+ $X2=4.995 $Y2=2.815
r122 47 91 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.995 $Y=3.245
+ $X2=5.055 $Y2=3.33
r123 47 52 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.995 $Y=3.245
+ $X2=4.995 $Y2=2.815
r124 43 46 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=4.03 $Y=2.115
+ $X2=4.03 $Y2=2.815
r125 41 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.03 $Y=3.245
+ $X2=4.03 $Y2=3.33
r126 41 46 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.03 $Y=3.245
+ $X2=4.03 $Y2=2.815
r127 37 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=3.245
+ $X2=3.13 $Y2=3.33
r128 37 39 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=3.13 $Y=3.245
+ $X2=3.13 $Y2=2.195
r129 36 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.23 $Y2=3.33
r130 35 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=3.33
+ $X2=3.13 $Y2=3.33
r131 35 36 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.045 $Y=3.33
+ $X2=2.395 $Y2=3.33
r132 31 34 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.23 $Y=2.115
+ $X2=2.23 $Y2=2.815
r133 29 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=3.33
r134 29 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=2.815
r135 25 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=3.245
+ $X2=1.28 $Y2=3.33
r136 25 27 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.28 $Y=3.245
+ $X2=1.28 $Y2=2.455
r137 21 24 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115
+ $X2=0.28 $Y2=2.815
r138 19 76 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r139 19 24 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r140 6 52 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.845
+ $Y=1.84 $X2=4.995 $Y2=2.815
r141 6 49 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=4.845
+ $Y=1.84 $X2=4.995 $Y2=2.115
r142 5 46 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.88
+ $Y=1.84 $X2=4.03 $Y2=2.815
r143 5 43 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.88
+ $Y=1.84 $X2=4.03 $Y2=2.115
r144 4 39 300 $w=1.7e-07 $l=4.23409e-07 $layer=licon1_PDIFF $count=2 $X=2.98
+ $Y=1.84 $X2=3.13 $Y2=2.195
r145 3 34 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.84 $X2=2.23 $Y2=2.815
r146 3 31 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.84 $X2=2.23 $Y2=2.115
r147 2 27 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.84 $X2=1.28 $Y2=2.455
r148 1 24 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r149 1 21 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__CLKBUF_8%X 1 2 3 4 5 6 7 8 27 31 35 36 37 38 41 47
+ 49 51 55 61 63 65 69 75 79 80 81 82 84 86 87 95 97
c154 84 0 1.31725e-19 $X=4.795 $Y=0.935
r155 92 95 0.64744 $w=4.43e-07 $l=2.5e-08 $layer=LI1_cond $X=4.932 $Y=1.69
+ $X2=4.932 $Y2=1.665
r156 87 92 7.04599 $w=1.68e-07 $l=1.08e-07 $layer=LI1_cond $X=5.04 $Y=1.775
+ $X2=4.932 $Y2=1.775
r157 87 95 0.776928 $w=4.43e-07 $l=3e-08 $layer=LI1_cond $X=4.932 $Y=1.635
+ $X2=4.932 $Y2=1.665
r158 87 91 6.03414 $w=4.43e-07 $l=2.33e-07 $layer=LI1_cond $X=4.932 $Y=1.635
+ $X2=4.932 $Y2=1.402
r159 86 91 2.77104 $w=4.43e-07 $l=1.07e-07 $layer=LI1_cond $X=4.932 $Y=1.295
+ $X2=4.932 $Y2=1.402
r160 86 97 7.56636 $w=4.43e-07 $l=1.15e-07 $layer=LI1_cond $X=4.932 $Y=1.295
+ $X2=4.932 $Y2=1.18
r161 83 84 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.57 $Y=0.935
+ $X2=4.795 $Y2=0.935
r162 77 84 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.795 $Y=1.02
+ $X2=4.795 $Y2=0.935
r163 77 97 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.795 $Y=1.02
+ $X2=4.795 $Y2=1.18
r164 73 83 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.57 $Y=0.85
+ $X2=4.57 $Y2=0.935
r165 73 75 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.57 $Y=0.85
+ $X2=4.57 $Y2=0.58
r166 69 71 36.7895 $w=2.58e-07 $l=8.3e-07 $layer=LI1_cond $X=4.515 $Y=1.985
+ $X2=4.515 $Y2=2.815
r167 67 92 27.2053 $w=1.68e-07 $l=4.17e-07 $layer=LI1_cond $X=4.515 $Y=1.775
+ $X2=4.932 $Y2=1.775
r168 67 69 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=4.515 $Y=1.86
+ $X2=4.515 $Y2=1.985
r169 66 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=0.935
+ $X2=3.64 $Y2=0.935
r170 65 83 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.485 $Y=0.935
+ $X2=4.57 $Y2=0.935
r171 65 66 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.485 $Y=0.935
+ $X2=3.725 $Y2=0.935
r172 64 81 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=3.68 $Y=1.775
+ $X2=3.547 $Y2=1.775
r173 63 67 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.385 $Y=1.775
+ $X2=4.515 $Y2=1.775
r174 63 64 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=4.385 $Y=1.775
+ $X2=3.68 $Y2=1.775
r175 59 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=0.85
+ $X2=3.64 $Y2=0.935
r176 59 61 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.64 $Y=0.85
+ $X2=3.64 $Y2=0.58
r177 55 57 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=3.547 $Y=1.985
+ $X2=3.547 $Y2=2.815
r178 53 81 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.547 $Y=1.86
+ $X2=3.547 $Y2=1.775
r179 53 55 5.43605 $w=2.63e-07 $l=1.25e-07 $layer=LI1_cond $X=3.547 $Y=1.86
+ $X2=3.547 $Y2=1.985
r180 52 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.865 $Y=0.935
+ $X2=2.74 $Y2=0.935
r181 51 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.555 $Y=0.935
+ $X2=3.64 $Y2=0.935
r182 51 52 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.555 $Y=0.935
+ $X2=2.865 $Y2=0.935
r183 50 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.845 $Y=1.775
+ $X2=2.715 $Y2=1.775
r184 49 81 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=3.415 $Y=1.775
+ $X2=3.547 $Y2=1.775
r185 49 50 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.415 $Y=1.775
+ $X2=2.845 $Y2=1.775
r186 45 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=0.85
+ $X2=2.74 $Y2=0.935
r187 45 47 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=2.74 $Y=0.85
+ $X2=2.74 $Y2=0.58
r188 41 43 36.7895 $w=2.58e-07 $l=8.3e-07 $layer=LI1_cond $X=2.715 $Y=1.985
+ $X2=2.715 $Y2=2.815
r189 39 79 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=1.86
+ $X2=2.715 $Y2=1.775
r190 39 41 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=2.715 $Y=1.86
+ $X2=2.715 $Y2=1.985
r191 37 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.615 $Y=0.935
+ $X2=2.74 $Y2=0.935
r192 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.615 $Y=0.935
+ $X2=1.945 $Y2=0.935
r193 35 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.585 $Y=1.775
+ $X2=2.715 $Y2=1.775
r194 35 36 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.585 $Y=1.775
+ $X2=1.88 $Y2=1.775
r195 31 33 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=1.747 $Y=1.985
+ $X2=1.747 $Y2=2.815
r196 29 36 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=1.747 $Y=1.86
+ $X2=1.88 $Y2=1.775
r197 29 31 5.43605 $w=2.63e-07 $l=1.25e-07 $layer=LI1_cond $X=1.747 $Y=1.86
+ $X2=1.747 $Y2=1.985
r198 25 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.78 $Y=0.85
+ $X2=1.945 $Y2=0.935
r199 25 27 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=1.78 $Y=0.85
+ $X2=1.78 $Y2=0.58
r200 8 71 400 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=4.38
+ $Y=1.84 $X2=4.535 $Y2=2.815
r201 8 69 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=4.38
+ $Y=1.84 $X2=4.535 $Y2=1.985
r202 7 57 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.43
+ $Y=1.84 $X2=3.58 $Y2=2.815
r203 7 55 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.43
+ $Y=1.84 $X2=3.58 $Y2=1.985
r204 6 43 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=1.84 $X2=2.68 $Y2=2.815
r205 6 41 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=1.84 $X2=2.68 $Y2=1.985
r206 5 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.63
+ $Y=1.84 $X2=1.78 $Y2=2.815
r207 5 31 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.63
+ $Y=1.84 $X2=1.78 $Y2=1.985
r208 4 75 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.37 $X2=4.57 $Y2=0.58
r209 3 61 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.5
+ $Y=0.37 $X2=3.64 $Y2=0.58
r210 2 47 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.64
+ $Y=0.37 $X2=2.78 $Y2=0.58
r211 1 27 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=1.615
+ $Y=0.37 $X2=1.78 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__CLKBUF_8%VGND 1 2 3 4 5 6 19 21 25 27 31 33 37 41 43
+ 45 47 49 54 59 68 71 74 77 81
c85 81 0 1.31725e-19 $X=5.04 $Y=0
r86 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r87 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r88 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r89 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r90 69 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r91 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r92 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r93 63 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r94 63 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r95 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r96 60 77 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=4.305 $Y=0 $X2=4.105
+ $Y2=0
r97 60 62 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.305 $Y=0 $X2=4.56
+ $Y2=0
r98 59 80 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5.057
+ $Y2=0
r99 59 62 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=4.56
+ $Y2=0
r100 58 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r101 58 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r102 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r103 55 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.21
+ $Y2=0
r104 55 57 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.6
+ $Y2=0
r105 54 77 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=3.905 $Y=0 $X2=4.105
+ $Y2=0
r106 54 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.905 $Y=0 $X2=3.6
+ $Y2=0
r107 53 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r108 53 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r109 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r110 50 65 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r111 50 52 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r112 49 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.28
+ $Y2=0
r113 49 52 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=0.72 $Y2=0
r114 47 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r115 47 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r116 43 80 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5 $Y=0.085
+ $X2=5.057 $Y2=0
r117 43 45 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.515
r118 39 77 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=0.085
+ $X2=4.105 $Y2=0
r119 39 41 12.3888 $w=3.98e-07 $l=4.3e-07 $layer=LI1_cond $X=4.105 $Y=0.085
+ $X2=4.105 $Y2=0.515
r120 35 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0
r121 35 37 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0.515
r122 34 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.28
+ $Y2=0
r123 33 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.21
+ $Y2=0
r124 33 34 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.045 $Y=0 $X2=2.445
+ $Y2=0
r125 29 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0
r126 29 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0.515
r127 28 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.28
+ $Y2=0
r128 27 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.28
+ $Y2=0
r129 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=0
+ $X2=1.445 $Y2=0
r130 23 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0
r131 23 25 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0.58
r132 19 65 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r133 19 21 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.58
r134 6 45 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.37 $X2=5 $Y2=0.515
r135 5 41 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=3.93
+ $Y=0.37 $X2=4.105 $Y2=0.515
r136 4 37 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.07
+ $Y=0.37 $X2=3.21 $Y2=0.515
r137 3 31 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.37 $X2=2.28 $Y2=0.515
r138 2 25 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.58
r139 1 21 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

