* File: sky130_fd_sc_ls__o32a_2.spice
* Created: Fri Aug 28 13:54:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o32a_2.pex.spice"
.subckt sky130_fd_sc_ls__o32a_2  VNB VPB A1 A2 A3 B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1007 N_X_M1007_d N_A_83_264#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.3404 PD=1.02 PS=2.4 NRD=0 NRS=14.184 M=1 R=4.93333 SA=75000.4
+ SB=75003.8 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1007_d N_A_83_264#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.8
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1005 N_A_349_74#_M1005_d N_A1_M1005_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.4
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g N_A_349_74#_M1005_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1003 N_A_349_74#_M1003_d N_A3_M1003_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1554 PD=1.09 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.4
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1002 N_A_83_264#_M1002_d N_B2_M1002_g N_A_349_74#_M1003_d VNB NSHORT L=0.15
+ W=0.74 AD=0.33855 AS=0.1295 PD=1.655 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75002.9 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1006 N_A_349_74#_M1006_d N_B1_M1006_g N_A_83_264#_M1002_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2627 AS=0.33855 PD=2.19 PS=1.655 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.9 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1008 N_X_M1008_d N_A_83_264#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1009 N_X_M1008_d N_A_83_264#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.307366 PD=1.42 PS=1.76453 NRD=1.7533 NRS=23.3051 M=1 R=7.46667
+ SA=75000.7 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1001 A_346_368# N_A1_M1001_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.274434 PD=1.27 PS=1.57547 NRD=15.7403 NRS=27.0678 M=1 R=6.66667
+ SA=75001.4 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1011 A_430_368# N_A2_M1011_g A_346_368# VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.135 PD=1.39 PS=1.27 NRD=27.5603 NRS=15.7403 M=1 R=6.66667 SA=75001.8
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1004 N_A_83_264#_M1004_d N_A3_M1004_g A_430_368# VPB PHIGHVT L=0.15 W=1
+ AD=0.21 AS=0.195 PD=1.42 PS=1.39 NRD=13.7703 NRS=27.5603 M=1 R=6.66667
+ SA=75002.3 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1000 A_652_368# N_B2_M1000_g N_A_83_264#_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.21 AS=0.21 PD=1.42 PS=1.42 NRD=30.5153 NRS=13.7703 M=1 R=6.66667
+ SA=75002.9 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1012_d N_B1_M1012_g A_652_368# VPB PHIGHVT L=0.15 W=1 AD=0.295
+ AS=0.21 PD=2.59 PS=1.42 NRD=1.9503 NRS=30.5153 M=1 R=6.66667 SA=75003.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ls__o32a_2.pxi.spice"
*
.ends
*
*
