# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ls__o2bb2ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__o2bb2ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.480000 1.630000 ;
        RECT 0.125000 1.630000 0.355000 2.415000 ;
        RECT 0.125000 2.415000 0.820000 2.450000 ;
        RECT 0.125000 2.450000 2.335000 2.585000 ;
        RECT 0.650000 2.585000 2.335000 2.620000 ;
        RECT 1.965000 1.350000 2.335000 1.680000 ;
        RECT 2.165000 1.680000 2.335000 2.450000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.375000 1.445000 1.795000 1.780000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.695000 1.350000 4.025000 1.720000 ;
        RECT 3.695000 1.720000 5.495000 1.780000 ;
        RECT 3.695000 1.780000 5.095000 1.890000 ;
        RECT 4.925000 1.350000 5.495000 1.720000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.345000 1.180000 4.675000 1.550000 ;
    END
  END B2
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 5.760000 0.245000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 5.950000 3.520000 ;
    END
  END VPB
  PIN Y
    ANTENNADIFFAREA  0.896000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.000000 0.595000 3.290000 1.130000 ;
        RECT 3.005000 1.130000 3.290000 2.060000 ;
        RECT 3.005000 2.060000 4.695000 2.230000 ;
        RECT 3.005000 2.230000 3.290000 2.980000 ;
        RECT 4.465000 2.230000 4.695000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  2.755000 0.445000 3.245000 ;
      RECT 0.145000  0.085000 0.475000 1.030000 ;
      RECT 0.645000  0.255000 1.910000 0.425000 ;
      RECT 0.645000  0.425000 0.975000 0.935000 ;
      RECT 0.650000  1.105000 2.675000 1.180000 ;
      RECT 0.650000  1.180000 1.405000 1.275000 ;
      RECT 0.650000  1.275000 0.980000 1.950000 ;
      RECT 0.650000  1.950000 1.995000 2.245000 ;
      RECT 1.155000  0.605000 1.405000 1.010000 ;
      RECT 1.155000  1.010000 2.675000 1.105000 ;
      RECT 1.185000  2.790000 1.515000 3.245000 ;
      RECT 1.580000  0.425000 1.910000 0.825000 ;
      RECT 1.720000  2.245000 1.995000 2.280000 ;
      RECT 2.080000  0.085000 2.340000 0.825000 ;
      RECT 2.505000  1.180000 2.675000 1.300000 ;
      RECT 2.505000  1.300000 2.835000 1.630000 ;
      RECT 2.505000  1.820000 2.835000 3.245000 ;
      RECT 2.570000  0.255000 3.790000 0.425000 ;
      RECT 2.570000  0.425000 2.820000 0.825000 ;
      RECT 3.460000  0.425000 3.790000 0.840000 ;
      RECT 3.460000  0.840000 5.645000 1.010000 ;
      RECT 3.460000  1.010000 3.790000 1.130000 ;
      RECT 3.460000  2.400000 3.790000 3.245000 ;
      RECT 3.960000  0.085000 4.290000 0.670000 ;
      RECT 3.965000  2.400000 4.295000 2.905000 ;
      RECT 3.965000  2.905000 5.195000 3.075000 ;
      RECT 4.470000  0.350000 4.690000 0.770000 ;
      RECT 4.470000  0.770000 5.645000 0.840000 ;
      RECT 4.865000  2.060000 5.195000 2.905000 ;
      RECT 4.870000  0.085000 5.215000 0.600000 ;
      RECT 5.315000  1.010000 5.645000 1.130000 ;
      RECT 5.395000  0.350000 5.645000 0.770000 ;
      RECT 5.395000  1.950000 5.645000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_ls__o2bb2ai_2
END LIBRARY
