* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 a_1320_119# a_1034_392# a_1234_119# VNB nshort w=420000u l=150000u
+  ad=9.87e+10p pd=1.31e+06u as=1.176e+11p ps=1.4e+06u
M1001 VGND a_1997_272# a_1972_74# VNB nshort w=420000u l=150000u
+  ad=1.59428e+12p pd=1.37e+07u as=8.82e+10p ps=1.26e+06u
M1002 a_1972_74# a_835_98# a_1745_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=4.687e+11p ps=3.25e+06u
M1003 a_1745_74# a_1034_392# a_1367_93# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1004 Q a_2399_424# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 a_312_81# a_27_88# a_225_81# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.499e+11p ps=2.87e+06u
M1006 a_300_464# D a_312_81# VNB nshort w=420000u l=150000u
+  ad=3.738e+11p pd=3.46e+06u as=0p ps=0u
M1007 VGND RESET_B a_1397_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 VPWR a_1367_93# a_1343_461# VPB phighvt w=420000u l=150000u
+  ad=2.19608e+12p pd=1.864e+07u as=1.134e+11p ps=1.38e+06u
M1009 a_1234_119# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.765e+11p pd=3.02e+06u as=0p ps=0u
M1010 a_2399_424# a_1745_74# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1011 a_300_464# D a_216_464# VPB phighvt w=640000u l=150000u
+  ad=9.687e+11p pd=6.63e+06u as=1.728e+11p ps=1.82e+06u
M1012 a_225_81# SCD a_545_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1013 a_1367_93# a_1234_119# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1014 a_1993_508# a_1034_392# a_1745_74# VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=4.42975e+11p ps=3.64e+06u
M1015 Q a_2399_424# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1016 a_1997_272# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1017 a_216_464# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1745_74# a_835_98# a_1367_93# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1397_119# a_1367_93# a_1320_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR SCE a_27_88# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1021 a_1997_272# a_1745_74# a_2135_74# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1022 a_535_464# a_27_88# a_300_464# VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1023 VPWR a_1745_74# a_1997_272# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_545_81# SCE a_300_464# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_2399_424# a_1745_74# VGND VNB nshort w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1026 VPWR SCD a_535_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR CLK a_835_98# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1028 VGND CLK a_835_98# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.619e+11p ps=2.38e+06u
M1029 a_1343_461# a_835_98# a_1234_119# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1034_392# a_835_98# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1031 a_1367_93# a_1234_119# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1034_392# a_835_98# VGND VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1033 VGND SCE a_27_88# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1034 VPWR a_1997_272# a_1993_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1234_119# a_835_98# a_300_464# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_2135_74# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND RESET_B a_225_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_300_464# RESET_B VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1234_119# a_1034_392# a_300_464# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
