* NGSPICE file created from sky130_fd_sc_ls__dlrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
M1000 VGND a_230_74# a_363_82# VNB nshort w=740000u l=150000u
+  ad=1.8561e+12p pd=1.54e+07u as=2.109e+11p ps=2.05e+06u
M1001 a_773_124# a_230_74# a_641_80# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.692e+11p ps=2.3e+06u
M1002 a_569_80# a_27_112# VGND VNB nshort w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1003 VPWR a_821_98# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=2.8212e+12p pd=2.104e+07u as=3.36e+11p ps=2.84e+06u
M1004 VGND a_821_98# a_1449_368# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1005 VPWR RESET_B a_821_98# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.92e+11p ps=2.94e+06u
M1006 VGND RESET_B a_1049_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1007 Q_N a_1449_368# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1008 VPWR a_821_98# a_1449_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1009 a_230_74# GATE VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1010 a_641_80# a_230_74# a_566_392# VPB phighvt w=1e+06u l=150000u
+  ad=3.328e+11p pd=2.77e+06u as=2.7e+11p ps=2.54e+06u
M1011 Q_N a_1449_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1012 VGND D a_27_112# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1013 a_1049_74# a_641_80# a_821_98# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1014 VGND a_1449_368# Q_N VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_230_74# GATE VPWR VPB phighvt w=840000u l=150000u
+  ad=2.898e+11p pd=2.37e+06u as=0p ps=0u
M1016 a_566_392# a_27_112# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_821_98# a_773_124# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_1449_368# Q_N VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR D a_27_112# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1020 a_757_508# a_363_82# a_641_80# VPB phighvt w=420000u l=150000u
+  ad=2.121e+11p pd=1.85e+06u as=0p ps=0u
M1021 VPWR a_821_98# a_757_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_641_80# a_363_82# a_569_80# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q a_821_98# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1024 VGND a_821_98# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_230_74# a_363_82# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1026 Q a_821_98# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_821_98# a_641_80# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

