# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__o311a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.105000 1.470000 8.035000 1.800000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.525000 1.220000 8.535000 1.300000 ;
        RECT 6.525000 1.300000 6.935000 1.550000 ;
        RECT 6.765000 1.130000 8.535000 1.220000 ;
        RECT 8.205000 1.300000 8.535000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.870000 1.420000 6.200000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.220000 4.165000 1.265000 ;
        RECT 2.505000 1.265000 2.910000 1.550000 ;
        RECT 2.740000 1.095000 4.165000 1.220000 ;
        RECT 3.995000 1.265000 4.165000 1.470000 ;
        RECT 3.995000 1.470000 5.360000 1.640000 ;
        RECT 4.925000 1.640000 5.360000 1.800000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.435000 3.825000 1.780000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.345400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.140000 0.945000 1.310000 ;
        RECT 0.125000 1.310000 0.355000 1.480000 ;
        RECT 0.125000 1.480000 0.895000 1.650000 ;
        RECT 0.565000 1.650000 0.895000 1.720000 ;
        RECT 0.565000 1.720000 1.895000 1.890000 ;
        RECT 0.565000 1.890000 0.895000 2.980000 ;
        RECT 0.615000 0.350000 0.945000 0.880000 ;
        RECT 0.615000 0.880000 2.070000 1.050000 ;
        RECT 0.615000 1.050000 0.945000 1.140000 ;
        RECT 1.565000 1.890000 1.895000 2.980000 ;
        RECT 1.740000 0.350000 2.070000 0.880000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.970000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 1.065000  2.060000 1.395000 3.245000 ;
      RECT 1.115000  0.085000 1.570000 0.680000 ;
      RECT 1.255000  1.220000 2.265000 1.550000 ;
      RECT 2.095000  1.550000 2.265000 1.720000 ;
      RECT 2.095000  1.720000 2.985000 1.890000 ;
      RECT 2.150000  2.060000 2.480000 3.245000 ;
      RECT 2.240000  0.085000 2.570000 1.050000 ;
      RECT 2.655000  1.890000 2.985000 1.950000 ;
      RECT 2.655000  1.950000 4.420000 1.970000 ;
      RECT 2.655000  1.970000 6.100000 2.120000 ;
      RECT 2.655000  2.120000 2.985000 2.980000 ;
      RECT 2.800000  0.255000 5.595000 0.425000 ;
      RECT 2.800000  0.425000 3.130000 0.925000 ;
      RECT 3.225000  2.290000 3.920000 3.245000 ;
      RECT 3.300000  0.595000 5.095000 0.765000 ;
      RECT 3.300000  0.765000 4.075000 0.925000 ;
      RECT 4.090000  1.940000 4.420000 1.950000 ;
      RECT 4.090000  2.120000 6.100000 2.140000 ;
      RECT 4.090000  2.140000 4.420000 2.980000 ;
      RECT 4.335000  0.935000 4.585000 1.130000 ;
      RECT 4.335000  1.130000 5.700000 1.300000 ;
      RECT 4.590000  2.310000 4.920000 2.370000 ;
      RECT 4.590000  2.370000 7.575000 2.395000 ;
      RECT 4.590000  2.395000 6.550000 2.540000 ;
      RECT 4.590000  2.540000 4.920000 3.245000 ;
      RECT 4.765000  0.765000 5.095000 0.960000 ;
      RECT 5.150000  2.710000 6.550000 2.905000 ;
      RECT 5.150000  2.905000 8.525000 2.960000 ;
      RECT 5.265000  0.425000 5.595000 0.790000 ;
      RECT 5.265000  0.790000 8.525000 0.960000 ;
      RECT 5.530000  1.300000 5.700000 1.950000 ;
      RECT 5.530000  1.950000 6.100000 1.970000 ;
      RECT 5.750000  2.140000 6.100000 2.200000 ;
      RECT 5.765000  0.085000 6.095000 0.620000 ;
      RECT 6.220000  2.960000 8.525000 3.075000 ;
      RECT 6.265000  0.370000 6.595000 0.790000 ;
      RECT 6.265000  0.960000 6.595000 1.050000 ;
      RECT 6.380000  1.970000 7.575000 2.370000 ;
      RECT 6.720000  2.565000 8.025000 2.735000 ;
      RECT 6.765000  0.085000 7.095000 0.620000 ;
      RECT 7.265000  0.350000 7.595000 0.790000 ;
      RECT 7.765000  0.085000 8.095000 0.620000 ;
      RECT 7.775000  1.970000 8.025000 2.565000 ;
      RECT 8.195000  1.970000 8.525000 2.905000 ;
      RECT 8.275000  0.350000 8.525000 0.790000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_ls__o311a_4
