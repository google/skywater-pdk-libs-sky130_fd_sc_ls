* NGSPICE file created from sky130_fd_sc_ls__or4_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__or4_1 A B C D VGND VNB VPB VPWR X
M1000 a_133_392# D a_44_392# VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=2.95e+11p ps=2.59e+06u
M1001 VGND C a_44_392# VNB nshort w=550000u l=150000u
+  ad=7.822e+11p pd=6.34e+06u as=3.96e+11p ps=3.64e+06u
M1002 a_44_392# D VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A a_44_392# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_44_392# B VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_331_392# VPB phighvt w=1e+06u l=150000u
+  ad=5.718e+11p pd=3.32e+06u as=4.2e+11p ps=2.84e+06u
M1006 X a_44_392# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1007 a_217_392# C a_133_392# VPB phighvt w=1e+06u l=150000u
+  ad=4.2e+11p pd=2.84e+06u as=0p ps=0u
M1008 X a_44_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1009 a_331_392# B a_217_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

