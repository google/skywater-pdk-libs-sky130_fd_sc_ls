* File: sky130_fd_sc_ls__mux2i_4.pex.spice
* Created: Fri Aug 28 13:30:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__MUX2I_4%A1 3 5 7 10 12 14 17 19 21 22 24 27 29 30 31
+ 46 47
c85 46 0 4.70544e-20 $X=1.72 $Y=1.515
r86 47 48 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=1.855 $Y=1.557
+ $X2=1.87 $Y2=1.557
r87 45 47 17.5865 $w=3.7e-07 $l=1.35e-07 $layer=POLY_cond $X=1.72 $Y=1.557
+ $X2=1.855 $Y2=1.557
r88 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.72
+ $Y=1.515 $X2=1.72 $Y2=1.515
r89 43 45 41.0351 $w=3.7e-07 $l=3.15e-07 $layer=POLY_cond $X=1.405 $Y=1.557
+ $X2=1.72 $Y2=1.557
r90 42 43 6.51351 $w=3.7e-07 $l=5e-08 $layer=POLY_cond $X=1.355 $Y=1.557
+ $X2=1.405 $Y2=1.557
r91 41 42 52.1081 $w=3.7e-07 $l=4e-07 $layer=POLY_cond $X=0.955 $Y=1.557
+ $X2=1.355 $Y2=1.557
r92 40 41 3.90811 $w=3.7e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.557
+ $X2=0.955 $Y2=1.557
r93 38 40 29.3108 $w=3.7e-07 $l=2.25e-07 $layer=POLY_cond $X=0.7 $Y=1.557
+ $X2=0.925 $Y2=1.557
r94 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.7
+ $Y=1.515 $X2=0.7 $Y2=1.515
r95 36 38 25.4027 $w=3.7e-07 $l=1.95e-07 $layer=POLY_cond $X=0.505 $Y=1.557
+ $X2=0.7 $Y2=1.557
r96 35 36 1.3027 $w=3.7e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.505 $Y2=1.557
r97 31 46 1.07204 $w=4.28e-07 $l=4e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.72
+ $Y2=1.565
r98 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r99 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r100 29 39 0.53602 $w=4.28e-07 $l=2e-08 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.7
+ $Y2=1.565
r101 25 48 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.87 $Y=1.35
+ $X2=1.87 $Y2=1.557
r102 25 27 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.87 $Y=1.35
+ $X2=1.87 $Y2=0.795
r103 22 47 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.557
r104 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r105 19 43 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.557
r106 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r107 15 42 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.355 $Y=1.35
+ $X2=1.355 $Y2=1.557
r108 15 17 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.355 $Y=1.35
+ $X2=1.355 $Y2=0.795
r109 12 41 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.557
r110 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r111 8 40 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=1.557
r112 8 10 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=0.795
r113 5 36 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.557
r114 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r115 1 35 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r116 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_4%A0 3 5 7 10 12 14 17 19 21 22 23 26 29 30 32
+ 33 34 35
c86 5 0 1.11086e-19 $X=2.315 $Y=1.765
r87 48 49 3.9187 $w=3.69e-07 $l=3e-08 $layer=POLY_cond $X=3.275 $Y=1.557
+ $X2=3.305 $Y2=1.557
r88 46 48 26.7778 $w=3.69e-07 $l=2.05e-07 $layer=POLY_cond $X=3.07 $Y=1.557
+ $X2=3.275 $Y2=1.557
r89 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.515 $X2=3.07 $Y2=1.515
r90 44 46 34.6152 $w=3.69e-07 $l=2.65e-07 $layer=POLY_cond $X=2.805 $Y=1.557
+ $X2=3.07 $Y2=1.557
r91 43 44 0.653117 $w=3.69e-07 $l=5e-09 $layer=POLY_cond $X=2.8 $Y=1.557
+ $X2=2.805 $Y2=1.557
r92 42 47 10.37 $w=4e-07 $l=3.4e-07 $layer=LI1_cond $X=2.73 $Y=1.565 $X2=3.07
+ $Y2=1.565
r93 41 43 9.14363 $w=3.69e-07 $l=7e-08 $layer=POLY_cond $X=2.73 $Y=1.557 $X2=2.8
+ $Y2=1.557
r94 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.73
+ $Y=1.515 $X2=2.73 $Y2=1.515
r95 39 41 54.2087 $w=3.69e-07 $l=4.15e-07 $layer=POLY_cond $X=2.315 $Y=1.557
+ $X2=2.73 $Y2=1.557
r96 38 39 1.95935 $w=3.69e-07 $l=1.5e-08 $layer=POLY_cond $X=2.3 $Y=1.557
+ $X2=2.315 $Y2=1.557
r97 35 47 1.525 $w=4e-07 $l=5e-08 $layer=LI1_cond $X=3.12 $Y=1.565 $X2=3.07
+ $Y2=1.565
r98 34 42 2.745 $w=4e-07 $l=9e-08 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.73
+ $Y2=1.565
r99 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.805 $Y=1.765
+ $X2=3.805 $Y2=2.4
r100 29 30 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.805 $Y=1.675
+ $X2=3.805 $Y2=1.765
r101 28 33 18.8402 $w=1.65e-07 $l=9.40744e-08 $layer=POLY_cond $X=3.805 $Y=1.5
+ $X2=3.762 $Y2=1.425
r102 28 29 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.805 $Y=1.5
+ $X2=3.805 $Y2=1.675
r103 24 33 18.8402 $w=1.65e-07 $l=9.94987e-08 $layer=POLY_cond $X=3.705 $Y=1.35
+ $X2=3.762 $Y2=1.425
r104 24 26 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.705 $Y=1.35
+ $X2=3.705 $Y2=0.795
r105 23 49 29.2437 $w=3.69e-07 $l=1.71184e-07 $layer=POLY_cond $X=3.395 $Y=1.425
+ $X2=3.305 $Y2=1.557
r106 22 33 6.66866 $w=1.5e-07 $l=1.32e-07 $layer=POLY_cond $X=3.63 $Y=1.425
+ $X2=3.762 $Y2=1.425
r107 22 23 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=3.63 $Y=1.425
+ $X2=3.395 $Y2=1.425
r108 19 49 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.305 $Y=1.765
+ $X2=3.305 $Y2=1.557
r109 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.305 $Y=1.765
+ $X2=3.305 $Y2=2.4
r110 15 48 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.275 $Y=1.35
+ $X2=3.275 $Y2=1.557
r111 15 17 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.275 $Y=1.35
+ $X2=3.275 $Y2=0.795
r112 12 44 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.805 $Y=1.765
+ $X2=2.805 $Y2=1.557
r113 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.805 $Y=1.765
+ $X2=2.805 $Y2=2.4
r114 8 43 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.8 $Y=1.35 $X2=2.8
+ $Y2=1.557
r115 8 10 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.8 $Y=1.35 $X2=2.8
+ $Y2=0.795
r116 5 39 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.315 $Y=1.765
+ $X2=2.315 $Y2=1.557
r117 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.315 $Y=1.765
+ $X2=2.315 $Y2=2.4
r118 1 38 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.3 $Y=1.35 $X2=2.3
+ $Y2=1.557
r119 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.3 $Y=1.35 $X2=2.3
+ $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_4%A_1030_268# 1 2 7 9 10 12 13 15 16 18 19 21
+ 24 26 28 31 33 38 42 44 48 51 55 58 59
c127 33 0 9.92943e-20 $X=6.67 $Y=1.505
r128 65 66 43.6405 $w=3.7e-07 $l=3.35e-07 $layer=POLY_cond $X=6.335 $Y=1.552
+ $X2=6.67 $Y2=1.552
r129 64 65 25.4027 $w=3.7e-07 $l=1.95e-07 $layer=POLY_cond $X=6.14 $Y=1.552
+ $X2=6.335 $Y2=1.552
r130 63 64 51.4568 $w=3.7e-07 $l=3.95e-07 $layer=POLY_cond $X=5.745 $Y=1.552
+ $X2=6.14 $Y2=1.552
r131 62 63 7.16487 $w=3.7e-07 $l=5.5e-08 $layer=POLY_cond $X=5.69 $Y=1.552
+ $X2=5.745 $Y2=1.552
r132 55 68 11.7243 $w=3.7e-07 $l=9e-08 $layer=POLY_cond $X=6.675 $Y=1.552
+ $X2=6.765 $Y2=1.552
r133 55 66 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=6.675 $Y=1.552
+ $X2=6.67 $Y2=1.552
r134 51 59 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=9.74 $Y=1.71 $X2=9.74
+ $Y2=1.01
r135 46 59 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.66 $Y=0.845
+ $X2=9.66 $Y2=1.01
r136 46 48 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=9.66 $Y=0.845
+ $X2=9.66 $Y2=0.555
r137 45 58 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.455 $Y=1.795
+ $X2=9.32 $Y2=1.795
r138 44 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.655 $Y=1.795
+ $X2=9.74 $Y2=1.71
r139 44 45 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=9.655 $Y=1.795
+ $X2=9.455 $Y2=1.795
r140 40 58 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.32 $Y=1.88
+ $X2=9.32 $Y2=1.795
r141 40 42 4.48172 $w=2.68e-07 $l=1.05e-07 $layer=LI1_cond $X=9.32 $Y=1.88
+ $X2=9.32 $Y2=1.985
r142 39 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=1.795
+ $X2=6.755 $Y2=1.795
r143 38 58 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.185 $Y=1.795
+ $X2=9.32 $Y2=1.795
r144 38 39 152.989 $w=1.68e-07 $l=2.345e-06 $layer=LI1_cond $X=9.185 $Y=1.795
+ $X2=6.84 $Y2=1.795
r145 36 62 48.8514 $w=3.7e-07 $l=3.75e-07 $layer=POLY_cond $X=5.315 $Y=1.552
+ $X2=5.69 $Y2=1.552
r146 36 60 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.315 $Y=1.552
+ $X2=5.24 $Y2=1.552
r147 35 36 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.315
+ $Y=1.505 $X2=5.315 $Y2=1.505
r148 33 56 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.755 $Y=1.505
+ $X2=6.755 $Y2=1.795
r149 33 55 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.675
+ $Y=1.505 $X2=6.675 $Y2=1.505
r150 33 35 47.32 $w=3.28e-07 $l=1.355e-06 $layer=LI1_cond $X=6.67 $Y=1.505
+ $X2=5.315 $Y2=1.505
r151 29 68 23.9667 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=6.765 $Y=1.34
+ $X2=6.765 $Y2=1.552
r152 29 31 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.765 $Y=1.34
+ $X2=6.765 $Y2=0.78
r153 26 66 23.9667 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=6.67 $Y=1.765
+ $X2=6.67 $Y2=1.552
r154 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.67 $Y=1.765
+ $X2=6.67 $Y2=2.4
r155 22 65 23.9667 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=6.335 $Y=1.34
+ $X2=6.335 $Y2=1.552
r156 22 24 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.335 $Y=1.34
+ $X2=6.335 $Y2=0.78
r157 19 64 23.9667 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=6.14 $Y=1.765
+ $X2=6.14 $Y2=1.552
r158 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.14 $Y=1.765
+ $X2=6.14 $Y2=2.4
r159 16 63 23.9667 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=5.745 $Y=1.34
+ $X2=5.745 $Y2=1.552
r160 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.745 $Y=1.34
+ $X2=5.745 $Y2=0.86
r161 13 62 23.9667 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=5.69 $Y=1.765
+ $X2=5.69 $Y2=1.552
r162 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.69 $Y=1.765
+ $X2=5.69 $Y2=2.4
r163 10 36 23.9667 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=5.315 $Y=1.34
+ $X2=5.315 $Y2=1.552
r164 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.315 $Y=1.34
+ $X2=5.315 $Y2=0.86
r165 7 60 23.9667 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=5.24 $Y=1.765
+ $X2=5.24 $Y2=1.552
r166 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.24 $Y=1.765
+ $X2=5.24 $Y2=2.4
r167 2 42 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=9.2
+ $Y=1.84 $X2=9.35 $Y2=1.985
r168 1 48 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=9.45
+ $Y=0.41 $X2=9.66 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_4%S 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 35 36 37 38 65
c108 28 0 1.15153e-19 $X=9.375 $Y=1.26
c109 1 0 9.92943e-20 $X=7.17 $Y=1.765
r110 65 66 24.8454 $w=3.88e-07 $l=2e-07 $layer=POLY_cond $X=9.375 $Y=1.512
+ $X2=9.575 $Y2=1.512
r111 63 65 11.1804 $w=3.88e-07 $l=9e-08 $layer=POLY_cond $X=9.285 $Y=1.512
+ $X2=9.375 $Y2=1.512
r112 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.285
+ $Y=1.425 $X2=9.285 $Y2=1.425
r113 61 63 19.8763 $w=3.88e-07 $l=1.6e-07 $layer=POLY_cond $X=9.125 $Y=1.512
+ $X2=9.285 $Y2=1.512
r114 60 61 31.0567 $w=3.88e-07 $l=2.5e-07 $layer=POLY_cond $X=8.875 $Y=1.512
+ $X2=9.125 $Y2=1.512
r115 59 60 31.6778 $w=3.88e-07 $l=2.55e-07 $layer=POLY_cond $X=8.62 $Y=1.512
+ $X2=8.875 $Y2=1.512
r116 57 59 1.8634 $w=3.88e-07 $l=1.5e-08 $layer=POLY_cond $X=8.605 $Y=1.512
+ $X2=8.62 $Y2=1.512
r117 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.605
+ $Y=1.425 $X2=8.605 $Y2=1.425
r118 55 57 19.8763 $w=3.88e-07 $l=1.6e-07 $layer=POLY_cond $X=8.445 $Y=1.512
+ $X2=8.605 $Y2=1.512
r119 53 55 22.3608 $w=3.88e-07 $l=1.8e-07 $layer=POLY_cond $X=8.265 $Y=1.512
+ $X2=8.445 $Y2=1.512
r120 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.265
+ $Y=1.425 $X2=8.265 $Y2=1.425
r121 51 53 11.8015 $w=3.88e-07 $l=9.5e-08 $layer=POLY_cond $X=8.17 $Y=1.512
+ $X2=8.265 $Y2=1.512
r122 50 51 47.8273 $w=3.88e-07 $l=3.85e-07 $layer=POLY_cond $X=7.785 $Y=1.512
+ $X2=8.17 $Y2=1.512
r123 49 50 20.4974 $w=3.88e-07 $l=1.65e-07 $layer=POLY_cond $X=7.62 $Y=1.512
+ $X2=7.785 $Y2=1.512
r124 47 49 4.34794 $w=3.88e-07 $l=3.5e-08 $layer=POLY_cond $X=7.585 $Y=1.512
+ $X2=7.62 $Y2=1.512
r125 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.585
+ $Y=1.425 $X2=7.585 $Y2=1.425
r126 45 47 28.5722 $w=3.88e-07 $l=2.3e-07 $layer=POLY_cond $X=7.355 $Y=1.512
+ $X2=7.585 $Y2=1.512
r127 44 45 22.982 $w=3.88e-07 $l=1.85e-07 $layer=POLY_cond $X=7.17 $Y=1.512
+ $X2=7.355 $Y2=1.512
r128 38 64 2.40092 $w=3.58e-07 $l=7.5e-08 $layer=LI1_cond $X=9.36 $Y=1.36
+ $X2=9.285 $Y2=1.36
r129 37 64 12.965 $w=3.58e-07 $l=4.05e-07 $layer=LI1_cond $X=8.88 $Y=1.36
+ $X2=9.285 $Y2=1.36
r130 37 58 8.80338 $w=3.58e-07 $l=2.75e-07 $layer=LI1_cond $X=8.88 $Y=1.36
+ $X2=8.605 $Y2=1.36
r131 36 58 6.56252 $w=3.58e-07 $l=2.05e-07 $layer=LI1_cond $X=8.4 $Y=1.36
+ $X2=8.605 $Y2=1.36
r132 36 54 4.32166 $w=3.58e-07 $l=1.35e-07 $layer=LI1_cond $X=8.4 $Y=1.36
+ $X2=8.265 $Y2=1.36
r133 35 54 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=7.92 $Y=1.36
+ $X2=8.265 $Y2=1.36
r134 35 48 10.7241 $w=3.58e-07 $l=3.35e-07 $layer=LI1_cond $X=7.92 $Y=1.36
+ $X2=7.585 $Y2=1.36
r135 34 48 4.64178 $w=3.58e-07 $l=1.45e-07 $layer=LI1_cond $X=7.44 $Y=1.36
+ $X2=7.585 $Y2=1.36
r136 31 66 25.1189 $w=1.5e-07 $l=2.53e-07 $layer=POLY_cond $X=9.575 $Y=1.765
+ $X2=9.575 $Y2=1.512
r137 31 33 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.575 $Y=1.765
+ $X2=9.575 $Y2=2.26
r138 28 65 25.1189 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=9.375 $Y=1.26
+ $X2=9.375 $Y2=1.512
r139 28 30 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.375 $Y=1.26
+ $X2=9.375 $Y2=0.78
r140 25 61 25.1189 $w=1.5e-07 $l=2.53e-07 $layer=POLY_cond $X=9.125 $Y=1.765
+ $X2=9.125 $Y2=1.512
r141 25 27 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.125 $Y=1.765
+ $X2=9.125 $Y2=2.26
r142 22 60 25.1189 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=8.875 $Y=1.26
+ $X2=8.875 $Y2=1.512
r143 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.875 $Y=1.26
+ $X2=8.875 $Y2=0.78
r144 19 59 25.1189 $w=1.5e-07 $l=2.53e-07 $layer=POLY_cond $X=8.62 $Y=1.765
+ $X2=8.62 $Y2=1.512
r145 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.62 $Y=1.765
+ $X2=8.62 $Y2=2.4
r146 16 55 25.1189 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=8.445 $Y=1.26
+ $X2=8.445 $Y2=1.512
r147 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.445 $Y=1.26
+ $X2=8.445 $Y2=0.78
r148 13 51 25.1189 $w=1.5e-07 $l=2.53e-07 $layer=POLY_cond $X=8.17 $Y=1.765
+ $X2=8.17 $Y2=1.512
r149 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.17 $Y=1.765
+ $X2=8.17 $Y2=2.4
r150 10 50 25.1189 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=7.785 $Y=1.26
+ $X2=7.785 $Y2=1.512
r151 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.785 $Y=1.26
+ $X2=7.785 $Y2=0.78
r152 7 49 25.1189 $w=1.5e-07 $l=2.53e-07 $layer=POLY_cond $X=7.62 $Y=1.765
+ $X2=7.62 $Y2=1.512
r153 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.62 $Y=1.765
+ $X2=7.62 $Y2=2.4
r154 4 45 25.1189 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=7.355 $Y=1.26
+ $X2=7.355 $Y2=1.512
r155 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.355 $Y=1.26
+ $X2=7.355 $Y2=0.78
r156 1 44 25.1189 $w=1.5e-07 $l=2.53e-07 $layer=POLY_cond $X=7.17 $Y=1.765
+ $X2=7.17 $Y2=1.512
r157 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.17 $Y=1.765
+ $X2=7.17 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_4%Y 1 2 3 4 5 6 7 8 9 10 33 35 37 39 40 41 45
+ 49 51 53 59 61 63 67 69 70 73 75 77 78 79 86 91
c129 77 0 6.40318e-20 $X=2.08 $Y=2.035
r130 91 92 1.37742 $w=6.2e-07 $l=7e-08 $layer=LI1_cond $X=3.865 $Y=1.965
+ $X2=3.865 $Y2=2.035
r131 86 91 5.90323 $w=6.2e-07 $l=3e-07 $layer=LI1_cond $X=3.865 $Y=1.665
+ $X2=3.865 $Y2=1.965
r132 79 82 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.08 $Y=2.035
+ $X2=3.08 $Y2=2.23
r133 70 86 9.50836 $w=6.2e-07 $l=1.83712e-07 $layer=LI1_cond $X=4 $Y=1.55
+ $X2=3.865 $Y2=1.665
r134 69 85 4.20453 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=4 $Y=1.18 $X2=4
+ $Y2=1.057
r135 69 70 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4 $Y=1.18 $X2=4
+ $Y2=1.55
r136 68 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=2.035
+ $X2=3.08 $Y2=2.035
r137 67 92 8.52869 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=3.485 $Y=2.035
+ $X2=3.865 $Y2=2.035
r138 67 68 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.485 $Y=2.035
+ $X2=3.245 $Y2=2.035
r139 64 78 7.45506 $w=2.07e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=1.057
+ $X2=2.085 $Y2=1.057
r140 64 66 36.9252 $w=2.43e-07 $l=7.85e-07 $layer=LI1_cond $X=2.25 $Y=1.057
+ $X2=3.035 $Y2=1.057
r141 63 85 2.90557 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=3.915 $Y=1.057
+ $X2=4 $Y2=1.057
r142 63 66 41.3939 $w=2.43e-07 $l=8.8e-07 $layer=LI1_cond $X=3.915 $Y=1.057
+ $X2=3.035 $Y2=1.057
r143 62 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=2.035
+ $X2=2.08 $Y2=2.035
r144 61 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=2.035
+ $X2=3.08 $Y2=2.035
r145 61 62 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.915 $Y=2.035
+ $X2=2.245 $Y2=2.035
r146 57 78 0.261258 $w=3.3e-07 $l=1.22e-07 $layer=LI1_cond $X=2.085 $Y=0.935
+ $X2=2.085 $Y2=1.057
r147 57 59 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.085 $Y=0.935
+ $X2=2.085 $Y2=0.68
r148 54 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=2.035
+ $X2=1.18 $Y2=2.035
r149 53 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.915 $Y=2.035
+ $X2=2.08 $Y2=2.035
r150 53 54 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.915 $Y=2.035
+ $X2=1.265 $Y2=2.035
r151 52 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=1.095
+ $X2=1.14 $Y2=1.095
r152 51 78 7.45506 $w=2.07e-07 $l=1.83016e-07 $layer=LI1_cond $X=1.92 $Y=1.095
+ $X2=2.085 $Y2=1.057
r153 51 52 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.92 $Y=1.095
+ $X2=1.225 $Y2=1.095
r154 47 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=2.12
+ $X2=1.18 $Y2=2.035
r155 47 49 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.18 $Y=2.12
+ $X2=1.18 $Y2=2.57
r156 43 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=1.01
+ $X2=1.14 $Y2=1.095
r157 43 45 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.14 $Y=1.01
+ $X2=1.14 $Y2=0.82
r158 42 72 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=0.365 $Y=2.035
+ $X2=0.24 $Y2=1.97
r159 41 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=2.035
+ $X2=1.18 $Y2=2.035
r160 41 42 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.095 $Y=2.035
+ $X2=0.365 $Y2=2.035
r161 39 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=1.095
+ $X2=1.14 $Y2=1.095
r162 39 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.055 $Y=1.095
+ $X2=0.365 $Y2=1.095
r163 35 72 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=0.24 $Y=2.12 $X2=0.24
+ $Y2=1.97
r164 35 37 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=0.24 $Y=2.12
+ $X2=0.24 $Y2=2.4
r165 31 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.365 $Y2=1.095
r166 31 33 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=0.57
r167 10 91 300 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=2 $X=3.88
+ $Y=1.84 $X2=4.08 $Y2=1.965
r168 9 82 600 $w=1.7e-07 $l=4.79687e-07 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.84 $X2=3.08 $Y2=2.23
r169 8 77 300 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.035
r170 7 75 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.035
r171 7 49 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.57
r172 6 72 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r173 6 37 300 $w=1.7e-07 $l=6.28331e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.4
r174 5 85 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.78
+ $Y=0.425 $X2=3.92 $Y2=1.02
r175 4 66 182 $w=1.7e-07 $l=6.70242e-07 $layer=licon1_NDIFF $count=1 $X=2.875
+ $Y=0.425 $X2=3.035 $Y2=1.02
r176 3 59 91 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=2 $X=1.945
+ $Y=0.425 $X2=2.085 $Y2=0.68
r177 2 45 182 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.425 $X2=1.14 $Y2=0.82
r178 1 33 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.425 $X2=0.28 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_4%A_116_368# 1 2 3 4 15 17 18 21 25 27 29 32
r65 31 32 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=5.465 $Y=2.902
+ $X2=5.3 $Y2=2.902
r66 25 31 0.233829 $w=3.43e-07 $l=7e-09 $layer=LI1_cond $X=5.472 $Y=2.902
+ $X2=5.465 $Y2=2.902
r67 25 27 30.331 $w=3.43e-07 $l=9.08e-07 $layer=LI1_cond $X=5.472 $Y=2.902
+ $X2=6.38 $Y2=2.902
r68 24 29 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.715 $Y=2.99
+ $X2=1.59 $Y2=2.99
r69 24 32 233.888 $w=1.68e-07 $l=3.585e-06 $layer=LI1_cond $X=1.715 $Y=2.99
+ $X2=5.3 $Y2=2.99
r70 19 29 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=2.905
+ $X2=1.59 $Y2=2.99
r71 19 21 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=1.59 $Y=2.905
+ $X2=1.59 $Y2=2.455
r72 17 29 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.465 $Y=2.99
+ $X2=1.59 $Y2=2.99
r73 17 18 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.465 $Y=2.99
+ $X2=0.895 $Y2=2.99
r74 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.73 $Y=2.905
+ $X2=0.895 $Y2=2.99
r75 13 15 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.73 $Y=2.905
+ $X2=0.73 $Y2=2.415
r76 4 27 600 $w=1.7e-07 $l=1.05428e-06 $layer=licon1_PDIFF $count=1 $X=6.215
+ $Y=1.84 $X2=6.38 $Y2=2.815
r77 3 31 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.315
+ $Y=1.84 $X2=5.465 $Y2=2.815
r78 2 21 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.455
r79 1 15 300 $w=1.7e-07 $l=6.45659e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_4%A_478_368# 1 2 3 4 13 15 17 21 26 31 35 40
+ 42
r73 35 37 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.045 $Y=2.475
+ $X2=5.045 $Y2=2.65
r74 31 33 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.58 $Y=2.455
+ $X2=3.58 $Y2=2.65
r75 26 28 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.58 $Y=2.455
+ $X2=2.58 $Y2=2.65
r76 22 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.56 $Y=2.475
+ $X2=7.395 $Y2=2.475
r77 21 42 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.23 $Y=2.475
+ $X2=8.395 $Y2=2.475
r78 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.23 $Y=2.475
+ $X2=7.56 $Y2=2.475
r79 18 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.13 $Y=2.475
+ $X2=5.045 $Y2=2.475
r80 17 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.23 $Y=2.475
+ $X2=7.395 $Y2=2.475
r81 17 18 137.005 $w=1.68e-07 $l=2.1e-06 $layer=LI1_cond $X=7.23 $Y=2.475
+ $X2=5.13 $Y2=2.475
r82 16 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=2.65
+ $X2=3.58 $Y2=2.65
r83 15 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=2.65
+ $X2=5.045 $Y2=2.65
r84 15 16 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=4.96 $Y=2.65
+ $X2=3.745 $Y2=2.65
r85 14 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=2.65
+ $X2=2.58 $Y2=2.65
r86 13 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=2.65
+ $X2=3.58 $Y2=2.65
r87 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=2.65
+ $X2=2.745 $Y2=2.65
r88 4 42 300 $w=1.7e-07 $l=7.06028e-07 $layer=licon1_PDIFF $count=2 $X=8.245
+ $Y=1.84 $X2=8.395 $Y2=2.475
r89 3 40 300 $w=1.7e-07 $l=7.06028e-07 $layer=licon1_PDIFF $count=2 $X=7.245
+ $Y=1.84 $X2=7.395 $Y2=2.475
r90 2 31 600 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=1 $X=3.38
+ $Y=1.84 $X2=3.58 $Y2=2.455
r91 1 26 600 $w=1.7e-07 $l=7.03616e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.84 $X2=2.58 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_4%VPWR 1 2 3 4 5 6 19 23 27 31 33 36 37 39 43
+ 46 48 56 61 66 72 75 78 82
r130 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r131 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r132 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r133 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r134 70 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r135 70 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r136 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r137 67 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.01 $Y=3.33
+ $X2=8.885 $Y2=3.33
r138 67 69 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=9.01 $Y=3.33
+ $X2=9.36 $Y2=3.33
r139 66 81 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=9.635 $Y=3.33
+ $X2=9.857 $Y2=3.33
r140 66 69 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.635 $Y=3.33
+ $X2=9.36 $Y2=3.33
r141 65 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r142 65 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r143 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r144 62 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.06 $Y=3.33
+ $X2=7.895 $Y2=3.33
r145 62 64 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=8.06 $Y=3.33
+ $X2=8.4 $Y2=3.33
r146 61 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.76 $Y=3.33
+ $X2=8.885 $Y2=3.33
r147 61 64 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.76 $Y=3.33
+ $X2=8.4 $Y2=3.33
r148 60 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r149 60 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r150 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r151 57 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.06 $Y=3.33
+ $X2=6.895 $Y2=3.33
r152 57 59 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.06 $Y=3.33
+ $X2=7.44 $Y2=3.33
r153 56 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.73 $Y=3.33
+ $X2=7.895 $Y2=3.33
r154 56 59 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.73 $Y=3.33
+ $X2=7.44 $Y2=3.33
r155 55 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r156 54 55 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r157 50 54 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=6.48 $Y2=3.33
r158 50 51 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r159 48 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.73 $Y=3.33
+ $X2=6.895 $Y2=3.33
r160 48 54 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.73 $Y=3.33
+ $X2=6.48 $Y2=3.33
r161 46 55 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.48 $Y2=3.33
r162 46 51 1.33793 $w=4.9e-07 $l=4.8e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=0.24 $Y2=3.33
r163 42 43 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.915 $Y=2.03
+ $X2=6.08 $Y2=2.03
r164 37 81 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.8 $Y=3.245
+ $X2=9.857 $Y2=3.33
r165 37 39 36.6686 $w=3.28e-07 $l=1.05e-06 $layer=LI1_cond $X=9.8 $Y=3.245
+ $X2=9.8 $Y2=2.195
r166 34 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=3.245
+ $X2=8.885 $Y2=3.33
r167 34 36 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=8.885 $Y=3.245
+ $X2=8.885 $Y2=2.555
r168 33 45 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=2.22
+ $X2=8.885 $Y2=2.135
r169 33 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=8.885 $Y=2.22
+ $X2=8.885 $Y2=2.555
r170 29 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.895 $Y=3.245
+ $X2=7.895 $Y2=3.33
r171 29 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.895 $Y=3.245
+ $X2=7.895 $Y2=2.815
r172 25 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.895 $Y=3.245
+ $X2=6.895 $Y2=3.33
r173 25 27 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.895 $Y=3.245
+ $X2=6.895 $Y2=2.815
r174 23 45 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.76 $Y=2.135
+ $X2=8.885 $Y2=2.135
r175 23 43 174.845 $w=1.68e-07 $l=2.68e-06 $layer=LI1_cond $X=8.76 $Y=2.135
+ $X2=6.08 $Y2=2.135
r176 19 42 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=5.89 $Y=2.03
+ $X2=5.915 $Y2=2.03
r177 19 21 26.5365 $w=3.78e-07 $l=8.75e-07 $layer=LI1_cond $X=5.89 $Y=2.03
+ $X2=5.015 $Y2=2.03
r178 6 39 300 $w=1.7e-07 $l=4.23409e-07 $layer=licon1_PDIFF $count=2 $X=9.65
+ $Y=1.84 $X2=9.8 $Y2=2.195
r179 5 45 600 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=8.695
+ $Y=1.84 $X2=8.845 $Y2=2.135
r180 5 36 600 $w=1.7e-07 $l=7.86432e-07 $layer=licon1_PDIFF $count=1 $X=8.695
+ $Y=1.84 $X2=8.845 $Y2=2.555
r181 4 31 600 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=7.695
+ $Y=1.84 $X2=7.895 $Y2=2.815
r182 3 27 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.84 $X2=6.895 $Y2=2.815
r183 2 42 600 $w=1.7e-07 $l=2.54165e-07 $layer=licon1_PDIFF $count=1 $X=5.765
+ $Y=1.84 $X2=5.915 $Y2=2.03
r184 1 21 300 $w=1.7e-07 $l=5.96825e-07 $layer=licon1_PDIFF $count=2 $X=4.495
+ $Y=1.84 $X2=5.015 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_4%A_114_85# 1 2 3 4 15 17 18 21 23 26 28 29 31
+ 35 37 38 39 41
c109 35 0 1.15153e-19 $X=8.66 $Y=0.555
r110 43 44 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=7.57 $Y=0.665
+ $X2=7.57 $Y2=0.925
r111 41 43 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=7.57 $Y=0.555
+ $X2=7.57 $Y2=0.665
r112 38 39 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.355 $Y=0.705
+ $X2=5.525 $Y2=0.705
r113 33 35 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=8.66 $Y=0.84
+ $X2=8.66 $Y2=0.555
r114 32 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.735 $Y=0.925
+ $X2=7.57 $Y2=0.925
r115 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.495 $Y=0.925
+ $X2=8.66 $Y2=0.84
r116 31 32 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=8.495 $Y=0.925
+ $X2=7.735 $Y2=0.925
r117 29 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.405 $Y=0.665
+ $X2=7.57 $Y2=0.665
r118 29 39 122.652 $w=1.68e-07 $l=1.88e-06 $layer=LI1_cond $X=7.405 $Y=0.665
+ $X2=5.525 $Y2=0.665
r119 28 38 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.765 $Y=0.745
+ $X2=5.355 $Y2=0.745
r120 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.68 $Y=0.66
+ $X2=4.765 $Y2=0.745
r121 25 26 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.68 $Y=0.425
+ $X2=4.68 $Y2=0.66
r122 24 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=0.34
+ $X2=1.57 $Y2=0.34
r123 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.595 $Y=0.34
+ $X2=4.68 $Y2=0.425
r124 23 24 186.588 $w=1.68e-07 $l=2.86e-06 $layer=LI1_cond $X=4.595 $Y=0.34
+ $X2=1.735 $Y2=0.34
r125 19 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.425
+ $X2=1.57 $Y2=0.34
r126 19 21 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.57 $Y=0.425
+ $X2=1.57 $Y2=0.675
r127 17 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=0.34
+ $X2=1.57 $Y2=0.34
r128 17 18 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.405 $Y=0.34
+ $X2=0.875 $Y2=0.34
r129 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.71 $Y=0.425
+ $X2=0.875 $Y2=0.34
r130 13 15 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.71 $Y=0.425
+ $X2=0.71 $Y2=0.675
r131 4 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.52
+ $Y=0.41 $X2=8.66 $Y2=0.555
r132 3 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.43
+ $Y=0.41 $X2=7.57 $Y2=0.555
r133 2 21 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.425 $X2=1.57 $Y2=0.675
r134 1 15 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.425 $X2=0.71 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_4%A_475_85# 1 2 3 4 13 20 22 26 27
r44 26 27 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.55 $Y=1.045
+ $X2=6.385 $Y2=1.045
r45 24 27 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=5.53 $Y=1.085
+ $X2=6.385 $Y2=1.085
r46 22 24 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=4.425 $Y=1.085
+ $X2=5.53 $Y2=1.085
r47 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.34 $Y=1
+ $X2=4.425 $Y2=1.085
r48 19 20 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.34 $Y=0.765
+ $X2=4.34 $Y2=1
r49 15 18 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=2.585 $Y=0.68
+ $X2=3.49 $Y2=0.68
r50 13 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.255 $Y=0.68
+ $X2=4.34 $Y2=0.765
r51 13 18 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=4.255 $Y=0.68
+ $X2=3.49 $Y2=0.68
r52 4 26 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=6.41
+ $Y=0.41 $X2=6.55 $Y2=1.005
r53 3 24 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.39
+ $Y=0.49 $X2=5.53 $Y2=1.085
r54 2 18 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=3.35
+ $Y=0.425 $X2=3.49 $Y2=0.68
r55 1 15 182 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_NDIFF $count=1 $X=2.375
+ $Y=0.425 $X2=2.585 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__MUX2I_4%VGND 1 2 3 4 5 18 20 22 26 30 33 34 35 37 45
+ 55 56 59 63 70 76
r95 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r96 71 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r97 70 73 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.06 $Y=0 $X2=7.06
+ $Y2=0.325
r98 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r99 64 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r100 63 66 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.04 $Y=0 $X2=6.04
+ $Y2=0.325
r101 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r102 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r103 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r104 53 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=7.92
+ $Y2=0
r105 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r106 50 76 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.325 $Y=0 $X2=8.115
+ $Y2=0
r107 50 52 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=8.325 $Y=0
+ $X2=8.88 $Y2=0
r108 49 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r109 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r110 46 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.185 $Y=0 $X2=5.06
+ $Y2=0
r111 46 48 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.185 $Y=0
+ $X2=5.52 $Y2=0
r112 45 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.875 $Y=0 $X2=6.04
+ $Y2=0
r113 45 48 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.875 $Y=0
+ $X2=5.52 $Y2=0
r114 43 44 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r115 40 44 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=4.56
+ $Y2=0
r116 39 43 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=4.56
+ $Y2=0
r117 39 40 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r118 37 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.935 $Y=0 $X2=5.06
+ $Y2=0
r119 37 43 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.935 $Y=0
+ $X2=4.56 $Y2=0
r120 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r121 35 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r122 35 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r123 33 52 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.995 $Y=0
+ $X2=8.88 $Y2=0
r124 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.995 $Y=0 $X2=9.16
+ $Y2=0
r125 32 55 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=9.325 $Y=0
+ $X2=9.84 $Y2=0
r126 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.325 $Y=0 $X2=9.16
+ $Y2=0
r127 28 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.16 $Y=0.085
+ $X2=9.16 $Y2=0
r128 28 30 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=9.16 $Y=0.085
+ $X2=9.16 $Y2=0.555
r129 24 76 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.115 $Y=0.085
+ $X2=8.115 $Y2=0
r130 24 26 12.8964 $w=4.18e-07 $l=4.7e-07 $layer=LI1_cond $X=8.115 $Y=0.085
+ $X2=8.115 $Y2=0.555
r131 23 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.225 $Y=0 $X2=7.06
+ $Y2=0
r132 22 76 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=7.905 $Y=0 $X2=8.115
+ $Y2=0
r133 22 23 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.905 $Y=0
+ $X2=7.225 $Y2=0
r134 21 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.205 $Y=0 $X2=6.04
+ $Y2=0
r135 20 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.895 $Y=0 $X2=7.06
+ $Y2=0
r136 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.895 $Y=0 $X2=6.205
+ $Y2=0
r137 16 59 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.06 $Y=0.085
+ $X2=5.06 $Y2=0
r138 16 18 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=5.06 $Y=0.085
+ $X2=5.06 $Y2=0.325
r139 5 30 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=8.95
+ $Y=0.41 $X2=9.16 $Y2=0.555
r140 4 26 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=7.86
+ $Y=0.41 $X2=8.115 $Y2=0.555
r141 3 73 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=6.84
+ $Y=0.41 $X2=7.06 $Y2=0.325
r142 2 66 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=5.82
+ $Y=0.49 $X2=6.04 $Y2=0.325
r143 1 18 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.875
+ $Y=0.18 $X2=5.02 $Y2=0.325
.ends

