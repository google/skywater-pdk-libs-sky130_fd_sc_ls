* File: sky130_fd_sc_ls__and3_2.pxi.spice
* Created: Wed Sep  2 10:54:51 2020
* 
x_PM_SKY130_FD_SC_LS__AND3_2%A N_A_c_56_n N_A_c_57_n N_A_c_63_n N_A_M1000_g
+ N_A_c_58_n N_A_M1006_g A A A N_A_c_61_n PM_SKY130_FD_SC_LS__AND3_2%A
x_PM_SKY130_FD_SC_LS__AND3_2%B N_B_c_92_n N_B_M1008_g N_B_c_93_n N_B_M1005_g B B
+ PM_SKY130_FD_SC_LS__AND3_2%B
x_PM_SKY130_FD_SC_LS__AND3_2%C N_C_c_125_n N_C_M1003_g N_C_c_126_n N_C_M1002_g C
+ PM_SKY130_FD_SC_LS__AND3_2%C
x_PM_SKY130_FD_SC_LS__AND3_2%A_41_384# N_A_41_384#_M1006_s N_A_41_384#_M1000_s
+ N_A_41_384#_M1008_d N_A_41_384#_M1007_g N_A_41_384#_c_163_n
+ N_A_41_384#_M1001_g N_A_41_384#_M1009_g N_A_41_384#_c_164_n
+ N_A_41_384#_M1004_g N_A_41_384#_c_159_n N_A_41_384#_c_174_n
+ N_A_41_384#_c_191_n N_A_41_384#_c_166_n N_A_41_384#_c_160_n
+ N_A_41_384#_c_167_n N_A_41_384#_c_168_n N_A_41_384#_c_161_n
+ N_A_41_384#_c_162_n PM_SKY130_FD_SC_LS__AND3_2%A_41_384#
x_PM_SKY130_FD_SC_LS__AND3_2%VPWR N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_M1004_s
+ N_VPWR_c_249_n N_VPWR_c_250_n N_VPWR_c_251_n N_VPWR_c_252_n N_VPWR_c_253_n
+ N_VPWR_c_254_n VPWR N_VPWR_c_255_n N_VPWR_c_256_n N_VPWR_c_248_n
+ PM_SKY130_FD_SC_LS__AND3_2%VPWR
x_PM_SKY130_FD_SC_LS__AND3_2%X N_X_M1007_s N_X_M1001_d N_X_c_291_n N_X_c_294_n
+ N_X_c_295_n N_X_c_292_n X PM_SKY130_FD_SC_LS__AND3_2%X
x_PM_SKY130_FD_SC_LS__AND3_2%VGND N_VGND_M1003_d N_VGND_M1009_d N_VGND_c_331_n
+ N_VGND_c_332_n N_VGND_c_333_n VGND N_VGND_c_334_n N_VGND_c_335_n
+ N_VGND_c_336_n N_VGND_c_337_n PM_SKY130_FD_SC_LS__AND3_2%VGND
cc_1 VNB N_A_c_56_n 0.00691849f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.485
cc_2 VNB N_A_c_57_n 0.0113576f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.755
cc_3 VNB N_A_c_58_n 0.0324727f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.57
cc_4 VNB N_A_M1006_g 0.0117117f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1
cc_5 VNB A 0.045212f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.47
cc_6 VNB N_A_c_61_n 0.0476697f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.405
cc_7 VNB N_B_c_92_n 0.019964f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.485
cc_8 VNB N_B_c_93_n 0.0152038f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.34
cc_9 VNB B 0.0034927f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.395
cc_10 VNB N_C_c_125_n 0.0185142f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.485
cc_11 VNB N_C_c_126_n 0.0217857f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.34
cc_12 VNB C 0.00354858f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.395
cc_13 VNB N_A_41_384#_M1007_g 0.0222518f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_14 VNB N_A_41_384#_M1009_g 0.0231292f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.405
cc_15 VNB N_A_41_384#_c_159_n 0.0137129f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.462
cc_16 VNB N_A_41_384#_c_160_n 0.0199411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_41_384#_c_161_n 0.00344604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_41_384#_c_162_n 0.0586758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_248_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_X_c_291_n 0.00296545f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1
cc_21 VNB N_X_c_292_n 0.00598001f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.405
cc_22 VNB X 0.00379924f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.405
cc_23 VNB N_VGND_c_331_n 0.0199076f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1
cc_24 VNB N_VGND_c_332_n 0.0451591f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_25 VNB N_VGND_c_333_n 0.0275707f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.47
cc_26 VNB N_VGND_c_334_n 0.0441425f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.405
cc_27 VNB N_VGND_c_335_n 0.0188369f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.405
cc_28 VNB N_VGND_c_336_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.462
cc_29 VNB N_VGND_c_337_n 0.214004f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.462
cc_30 VPB N_A_c_57_n 0.00613573f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.755
cc_31 VPB N_A_c_63_n 0.0274896f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.845
cc_32 VPB N_B_c_92_n 0.0328618f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.485
cc_33 VPB B 0.00303485f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.395
cc_34 VPB N_C_c_126_n 0.0355367f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.34
cc_35 VPB C 0.00165155f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.395
cc_36 VPB N_A_41_384#_c_163_n 0.0167036f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_A_41_384#_c_164_n 0.0174223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_A_41_384#_c_159_n 0.0119354f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.462
cc_39 VPB N_A_41_384#_c_166_n 0.0027152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_41_384#_c_167_n 0.0358627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_41_384#_c_168_n 0.00353992f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_41_384#_c_162_n 0.0297967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_249_n 0.0268291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_250_n 0.0173596f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.405
cc_45 VPB N_VPWR_c_251_n 0.0128289f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.405
cc_46 VPB N_VPWR_c_252_n 0.0632115f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=0.405
cc_47 VPB N_VPWR_c_253_n 0.025575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_254_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.462
cc_49 VPB N_VPWR_c_255_n 0.019175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_256_n 0.0285346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_248_n 0.080923f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_X_c_294_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=0.47
cc_53 VPB N_X_c_295_n 9.66679e-19 $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.405
cc_54 VPB N_X_c_292_n 0.00129283f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.405
cc_55 N_A_c_56_n N_B_c_92_n 0.0168476f $X=0.575 $Y=1.485 $X2=-0.19 $Y2=-0.245
cc_56 N_A_c_63_n N_B_c_92_n 0.025891f $X=0.575 $Y=1.845 $X2=-0.19 $Y2=-0.245
cc_57 N_A_c_58_n N_B_c_93_n 8.67721e-19 $X=0.59 $Y=0.57 $X2=0 $Y2=0
cc_58 N_A_M1006_g N_B_c_93_n 0.0245557f $X=0.59 $Y=1 $X2=0 $Y2=0
cc_59 A N_B_c_93_n 0.0109386f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_60 N_A_c_56_n B 0.00119213f $X=0.575 $Y=1.485 $X2=0 $Y2=0
cc_61 N_A_M1006_g B 0.00223423f $X=0.59 $Y=1 $X2=0 $Y2=0
cc_62 A B 0.01291f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_63 A N_C_c_125_n 0.00108821f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_64 N_A_c_56_n N_A_41_384#_c_159_n 0.00393408f $X=0.575 $Y=1.485 $X2=0 $Y2=0
cc_65 N_A_c_57_n N_A_41_384#_c_159_n 0.00966862f $X=0.575 $Y=1.755 $X2=0 $Y2=0
cc_66 N_A_c_63_n N_A_41_384#_c_159_n 0.00746901f $X=0.575 $Y=1.845 $X2=0 $Y2=0
cc_67 N_A_M1006_g N_A_41_384#_c_159_n 0.0015053f $X=0.59 $Y=1 $X2=0 $Y2=0
cc_68 N_A_c_63_n N_A_41_384#_c_174_n 0.0162305f $X=0.575 $Y=1.845 $X2=0 $Y2=0
cc_69 N_A_M1006_g N_A_41_384#_c_160_n 0.012609f $X=0.59 $Y=1 $X2=0 $Y2=0
cc_70 A N_A_41_384#_c_160_n 0.0277772f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_71 N_A_c_61_n N_A_41_384#_c_160_n 0.00188139f $X=0.515 $Y=0.405 $X2=0 $Y2=0
cc_72 N_A_c_63_n N_A_41_384#_c_167_n 0.0121204f $X=0.575 $Y=1.845 $X2=0 $Y2=0
cc_73 N_A_c_63_n N_A_41_384#_c_168_n 8.6665e-19 $X=0.575 $Y=1.845 $X2=0 $Y2=0
cc_74 N_A_c_63_n N_VPWR_c_249_n 0.00635764f $X=0.575 $Y=1.845 $X2=0 $Y2=0
cc_75 N_A_c_63_n N_VPWR_c_256_n 0.00435405f $X=0.575 $Y=1.845 $X2=0 $Y2=0
cc_76 N_A_c_63_n N_VPWR_c_248_n 0.00484898f $X=0.575 $Y=1.845 $X2=0 $Y2=0
cc_77 A N_VGND_c_331_n 0.0214717f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_78 A N_VGND_c_334_n 0.0794507f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_79 N_A_c_61_n N_VGND_c_334_n 0.0116176f $X=0.515 $Y=0.405 $X2=0 $Y2=0
cc_80 N_A_c_58_n N_VGND_c_337_n 0.00642106f $X=0.59 $Y=0.57 $X2=0 $Y2=0
cc_81 A N_VGND_c_337_n 0.0425626f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_82 N_A_c_61_n N_VGND_c_337_n 0.00862283f $X=0.515 $Y=0.405 $X2=0 $Y2=0
cc_83 N_B_c_93_n N_C_c_125_n 0.0316904f $X=1.16 $Y=1.43 $X2=-0.19 $Y2=-0.245
cc_84 B N_C_c_125_n 0.00818659f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_85 N_B_c_92_n N_C_c_126_n 0.0494194f $X=1.145 $Y=1.845 $X2=0 $Y2=0
cc_86 N_B_c_92_n C 4.10391e-19 $X=1.145 $Y=1.845 $X2=0 $Y2=0
cc_87 B C 0.0282664f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_88 N_B_c_92_n N_A_41_384#_c_159_n 0.00174365f $X=1.145 $Y=1.845 $X2=0 $Y2=0
cc_89 B N_A_41_384#_c_159_n 0.0178438f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_90 N_B_c_92_n N_A_41_384#_c_174_n 0.0134337f $X=1.145 $Y=1.845 $X2=0 $Y2=0
cc_91 B N_A_41_384#_c_174_n 0.0214868f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_92 N_B_c_93_n N_A_41_384#_c_160_n 0.0016883f $X=1.16 $Y=1.43 $X2=0 $Y2=0
cc_93 B N_A_41_384#_c_160_n 0.00709791f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_94 N_B_c_92_n N_A_41_384#_c_167_n 8.56176e-19 $X=1.145 $Y=1.845 $X2=0 $Y2=0
cc_95 N_B_c_92_n N_A_41_384#_c_168_n 0.0105063f $X=1.145 $Y=1.845 $X2=0 $Y2=0
cc_96 B N_A_41_384#_c_168_n 0.00713841f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_97 N_B_c_92_n N_VPWR_c_249_n 0.00615821f $X=1.145 $Y=1.845 $X2=0 $Y2=0
cc_98 N_B_c_92_n N_VPWR_c_253_n 0.00435405f $X=1.145 $Y=1.845 $X2=0 $Y2=0
cc_99 N_B_c_92_n N_VPWR_c_248_n 0.00484898f $X=1.145 $Y=1.845 $X2=0 $Y2=0
cc_100 B A_133_136# 0.00402475f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_101 B A_247_136# 0.00221309f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_102 N_B_c_93_n N_VGND_c_334_n 4.78105e-19 $X=1.16 $Y=1.43 $X2=0 $Y2=0
cc_103 N_C_c_125_n N_A_41_384#_M1007_g 0.0193095f $X=1.55 $Y=1.43 $X2=0 $Y2=0
cc_104 N_C_c_126_n N_A_41_384#_c_163_n 0.0163252f $X=1.595 $Y=1.845 $X2=0 $Y2=0
cc_105 N_C_c_126_n N_A_41_384#_c_191_n 0.0137058f $X=1.595 $Y=1.845 $X2=0 $Y2=0
cc_106 C N_A_41_384#_c_191_n 0.0188937f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_107 N_C_c_126_n N_A_41_384#_c_166_n 0.00388306f $X=1.595 $Y=1.845 $X2=0 $Y2=0
cc_108 C N_A_41_384#_c_166_n 0.00689943f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_109 N_C_c_126_n N_A_41_384#_c_168_n 0.0164545f $X=1.595 $Y=1.845 $X2=0 $Y2=0
cc_110 C N_A_41_384#_c_168_n 0.00254579f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_111 N_C_c_125_n N_A_41_384#_c_161_n 0.00169384f $X=1.55 $Y=1.43 $X2=0 $Y2=0
cc_112 N_C_c_126_n N_A_41_384#_c_161_n 0.00147149f $X=1.595 $Y=1.845 $X2=0 $Y2=0
cc_113 C N_A_41_384#_c_161_n 0.0157355f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_114 N_C_c_126_n N_A_41_384#_c_162_n 0.0149163f $X=1.595 $Y=1.845 $X2=0 $Y2=0
cc_115 C N_A_41_384#_c_162_n 2.91011e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_116 N_C_c_126_n N_VPWR_c_250_n 0.00775644f $X=1.595 $Y=1.845 $X2=0 $Y2=0
cc_117 N_C_c_126_n N_VPWR_c_253_n 0.00435405f $X=1.595 $Y=1.845 $X2=0 $Y2=0
cc_118 N_C_c_126_n N_VPWR_c_248_n 0.00484898f $X=1.595 $Y=1.845 $X2=0 $Y2=0
cc_119 N_C_c_125_n N_VGND_c_331_n 0.0047463f $X=1.55 $Y=1.43 $X2=0 $Y2=0
cc_120 N_C_c_126_n N_VGND_c_331_n 9.95834e-19 $X=1.595 $Y=1.845 $X2=0 $Y2=0
cc_121 C N_VGND_c_331_n 0.00794902f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_122 N_C_c_125_n N_VGND_c_334_n 0.0038748f $X=1.55 $Y=1.43 $X2=0 $Y2=0
cc_123 N_C_c_125_n N_VGND_c_337_n 0.00454494f $X=1.55 $Y=1.43 $X2=0 $Y2=0
cc_124 N_A_41_384#_c_174_n N_VPWR_M1000_d 0.012296f $X=1.205 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_125 N_A_41_384#_c_191_n N_VPWR_M1002_d 0.0211931f $X=2.035 $Y=2.035 $X2=0
+ $Y2=0
cc_126 N_A_41_384#_c_166_n N_VPWR_M1002_d 0.00229907f $X=2.12 $Y=1.95 $X2=0
+ $Y2=0
cc_127 N_A_41_384#_c_174_n N_VPWR_c_249_n 0.0248957f $X=1.205 $Y=2.035 $X2=0
+ $Y2=0
cc_128 N_A_41_384#_c_167_n N_VPWR_c_249_n 0.0191765f $X=0.35 $Y=2.065 $X2=0
+ $Y2=0
cc_129 N_A_41_384#_c_168_n N_VPWR_c_249_n 0.0175495f $X=1.37 $Y=2.115 $X2=0
+ $Y2=0
cc_130 N_A_41_384#_c_163_n N_VPWR_c_250_n 0.0112588f $X=2.315 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A_41_384#_c_191_n N_VPWR_c_250_n 0.0258048f $X=2.035 $Y=2.035 $X2=0
+ $Y2=0
cc_132 N_A_41_384#_c_168_n N_VPWR_c_250_n 0.0223823f $X=1.37 $Y=2.115 $X2=0
+ $Y2=0
cc_133 N_A_41_384#_c_162_n N_VPWR_c_250_n 4.45696e-19 $X=2.6 $Y=1.552 $X2=0
+ $Y2=0
cc_134 N_A_41_384#_c_164_n N_VPWR_c_252_n 0.0269315f $X=2.765 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A_41_384#_c_168_n N_VPWR_c_253_n 0.00794604f $X=1.37 $Y=2.115 $X2=0
+ $Y2=0
cc_136 N_A_41_384#_c_163_n N_VPWR_c_255_n 0.00445602f $X=2.315 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_A_41_384#_c_164_n N_VPWR_c_255_n 0.00422942f $X=2.765 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A_41_384#_c_167_n N_VPWR_c_256_n 0.00798f $X=0.35 $Y=2.065 $X2=0 $Y2=0
cc_139 N_A_41_384#_c_163_n N_VPWR_c_248_n 0.00861719f $X=2.315 $Y=1.765 $X2=0
+ $Y2=0
cc_140 N_A_41_384#_c_164_n N_VPWR_c_248_n 0.00787748f $X=2.765 $Y=1.765 $X2=0
+ $Y2=0
cc_141 N_A_41_384#_c_167_n N_VPWR_c_248_n 0.0105742f $X=0.35 $Y=2.065 $X2=0
+ $Y2=0
cc_142 N_A_41_384#_c_168_n N_VPWR_c_248_n 0.0105585f $X=1.37 $Y=2.115 $X2=0
+ $Y2=0
cc_143 N_A_41_384#_M1007_g N_X_c_291_n 0.00562723f $X=2.13 $Y=0.78 $X2=0 $Y2=0
cc_144 N_A_41_384#_M1009_g N_X_c_291_n 4.72567e-19 $X=2.6 $Y=0.78 $X2=0 $Y2=0
cc_145 N_A_41_384#_c_163_n N_X_c_294_n 0.0159493f $X=2.315 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A_41_384#_c_164_n N_X_c_294_n 0.0118876f $X=2.765 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A_41_384#_c_163_n N_X_c_295_n 0.00187137f $X=2.315 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A_41_384#_c_164_n N_X_c_295_n 0.00198375f $X=2.765 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_41_384#_c_161_n N_X_c_295_n 7.18422e-19 $X=2.22 $Y=1.505 $X2=0 $Y2=0
cc_150 N_A_41_384#_c_162_n N_X_c_295_n 0.00458278f $X=2.6 $Y=1.552 $X2=0 $Y2=0
cc_151 N_A_41_384#_M1007_g N_X_c_292_n 9.76257e-19 $X=2.13 $Y=0.78 $X2=0 $Y2=0
cc_152 N_A_41_384#_c_163_n N_X_c_292_n 5.75089e-19 $X=2.315 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A_41_384#_M1009_g N_X_c_292_n 0.00712292f $X=2.6 $Y=0.78 $X2=0 $Y2=0
cc_154 N_A_41_384#_c_164_n N_X_c_292_n 0.00298674f $X=2.765 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A_41_384#_c_166_n N_X_c_292_n 0.00769572f $X=2.12 $Y=1.95 $X2=0 $Y2=0
cc_156 N_A_41_384#_c_161_n N_X_c_292_n 0.0236573f $X=2.22 $Y=1.505 $X2=0 $Y2=0
cc_157 N_A_41_384#_c_162_n N_X_c_292_n 0.0319436f $X=2.6 $Y=1.552 $X2=0 $Y2=0
cc_158 N_A_41_384#_M1007_g X 0.00442604f $X=2.13 $Y=0.78 $X2=0 $Y2=0
cc_159 N_A_41_384#_M1009_g X 0.0156684f $X=2.6 $Y=0.78 $X2=0 $Y2=0
cc_160 N_A_41_384#_c_161_n X 0.0162347f $X=2.22 $Y=1.505 $X2=0 $Y2=0
cc_161 N_A_41_384#_c_162_n X 0.00550476f $X=2.6 $Y=1.552 $X2=0 $Y2=0
cc_162 N_A_41_384#_M1007_g N_VGND_c_331_n 0.010364f $X=2.13 $Y=0.78 $X2=0 $Y2=0
cc_163 N_A_41_384#_M1009_g N_VGND_c_332_n 0.00878267f $X=2.6 $Y=0.78 $X2=0 $Y2=0
cc_164 N_A_41_384#_c_162_n N_VGND_c_332_n 0.00281053f $X=2.6 $Y=1.552 $X2=0
+ $Y2=0
cc_165 N_A_41_384#_M1009_g N_VGND_c_333_n 0.00565998f $X=2.6 $Y=0.78 $X2=0 $Y2=0
cc_166 N_A_41_384#_M1007_g N_VGND_c_335_n 0.00523933f $X=2.13 $Y=0.78 $X2=0
+ $Y2=0
cc_167 N_A_41_384#_M1009_g N_VGND_c_335_n 0.00548708f $X=2.6 $Y=0.78 $X2=0 $Y2=0
cc_168 N_A_41_384#_M1007_g N_VGND_c_337_n 0.00533081f $X=2.13 $Y=0.78 $X2=0
+ $Y2=0
cc_169 N_A_41_384#_M1009_g N_VGND_c_337_n 0.00533081f $X=2.6 $Y=0.78 $X2=0 $Y2=0
cc_170 N_VPWR_c_250_n N_X_c_294_n 0.0269152f $X=2.04 $Y=2.455 $X2=0 $Y2=0
cc_171 N_VPWR_c_255_n N_X_c_294_n 0.0153846f $X=2.895 $Y=3.33 $X2=0 $Y2=0
cc_172 N_VPWR_c_248_n N_X_c_294_n 0.0126213f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_173 N_VPWR_c_252_n N_X_c_292_n 0.0453496f $X=3.06 $Y=1.985 $X2=0 $Y2=0
cc_174 N_VPWR_c_252_n N_VGND_c_333_n 0.0108898f $X=3.06 $Y=1.985 $X2=0 $Y2=0
cc_175 X N_VGND_M1009_d 0.00398771f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_176 N_X_c_291_n N_VGND_c_331_n 0.0165499f $X=2.345 $Y=0.555 $X2=0 $Y2=0
cc_177 X N_VGND_c_331_n 0.0154525f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_178 N_X_c_291_n N_VGND_c_332_n 0.0016552f $X=2.345 $Y=0.555 $X2=0 $Y2=0
cc_179 X N_VGND_c_332_n 0.00191947f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_180 X N_VGND_c_333_n 0.0300887f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_181 N_X_c_291_n N_VGND_c_335_n 0.0121172f $X=2.345 $Y=0.555 $X2=0 $Y2=0
cc_182 N_X_c_291_n N_VGND_c_337_n 0.0115967f $X=2.345 $Y=0.555 $X2=0 $Y2=0
cc_183 X N_VGND_c_337_n 0.00618074f $X=2.555 $Y=0.84 $X2=0 $Y2=0
