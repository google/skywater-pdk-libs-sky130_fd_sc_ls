* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__mux2i_1 A0 A1 S VGND VNB VPB VPWR Y
M1000 a_426_74# a_114_74# VGND VNB nshort w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=4.6755e+11p ps=3.99e+06u
M1001 Y A0 a_426_74# VNB nshort w=740000u l=150000u
+  ad=5.217e+11p pd=2.89e+06u as=0p ps=0u
M1002 VPWR S a_223_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=5.754e+11p pd=5.09e+06u as=6.272e+11p ps=5.6e+06u
M1003 a_225_74# A1 Y VNB nshort w=740000u l=150000u
+  ad=4.218e+11p pd=4.1e+06u as=0p ps=0u
M1004 Y A0 a_223_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1005 a_399_368# a_114_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.272e+11p pd=5.6e+06u as=0p ps=0u
M1006 a_114_74# S VPWR VPB phighvt w=840000u l=150000u
+  ad=2.31e+11p pd=2.23e+06u as=0p ps=0u
M1007 a_114_74# S VGND VNB nshort w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1008 a_399_368# A1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND S a_225_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
