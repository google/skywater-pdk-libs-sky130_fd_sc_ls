# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__dfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__dfstp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.00000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475000 0.980000 0.805000 1.990000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685000 1.820000 11.465000 2.150000 ;
        RECT 11.100000 0.350000 11.465000 1.130000 ;
        RECT 11.155000 2.150000 11.465000 2.980000 ;
        RECT 11.295000 1.130000 11.465000 1.820000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.855000 1.920000 6.145000 1.965000 ;
        RECT 5.855000 1.965000 8.545000 2.105000 ;
        RECT 5.855000 2.105000 6.145000 2.150000 ;
        RECT 8.255000 1.920000 8.545000 1.965000 ;
        RECT 8.255000 2.105000 8.545000 2.150000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315000 1.180000 1.775000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.000000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.000000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.000000 0.085000 ;
      RECT  0.000000  3.245000 12.000000 3.415000 ;
      RECT  0.115000  0.395000  0.365000 0.765000 ;
      RECT  0.115000  0.765000  0.285000 2.190000 ;
      RECT  0.115000  2.190000  2.615000 2.230000 ;
      RECT  0.115000  2.230000  1.795000 2.360000 ;
      RECT  0.115000  2.360000  0.365000 2.980000 ;
      RECT  0.545000  0.085000  0.795000 0.765000 ;
      RECT  0.565000  2.530000  0.895000 3.245000 ;
      RECT  0.975000  0.350000  1.435000 1.010000 ;
      RECT  0.975000  1.010000  1.145000 1.720000 ;
      RECT  0.975000  1.720000  2.275000 1.890000 ;
      RECT  0.975000  1.890000  1.455000 2.020000 ;
      RECT  1.575000  2.530000  1.905000 3.245000 ;
      RECT  1.615000  0.085000  1.865000 1.010000 ;
      RECT  1.625000  2.060000  2.615000 2.190000 ;
      RECT  1.945000  1.300000  2.275000 1.720000 ;
      RECT  2.045000  0.255000  3.115000 0.425000 ;
      RECT  2.045000  0.425000  2.215000 1.130000 ;
      RECT  2.105000  2.400000  2.275000 2.890000 ;
      RECT  2.105000  2.890000  3.795000 3.060000 ;
      RECT  2.445000  0.595000  2.775000 0.925000 ;
      RECT  2.445000  0.925000  2.615000 2.060000 ;
      RECT  2.445000  2.230000  2.615000 2.260000 ;
      RECT  2.445000  2.260000  2.945000 2.720000 ;
      RECT  2.785000  1.380000  3.115000 2.050000 ;
      RECT  2.945000  0.425000  3.115000 1.380000 ;
      RECT  3.115000  2.260000  3.455000 2.720000 ;
      RECT  3.285000  0.400000  3.615000 1.040000 ;
      RECT  3.285000  1.040000  4.255000 1.210000 ;
      RECT  3.285000  1.210000  3.455000 2.260000 ;
      RECT  3.625000  1.380000  3.915000 2.240000 ;
      RECT  3.625000  2.240000  4.915000 2.410000 ;
      RECT  3.625000  2.410000  3.795000 2.890000 ;
      RECT  4.070000  2.580000  4.575000 2.910000 ;
      RECT  4.070000  2.910000  4.240000 3.245000 ;
      RECT  4.085000  1.210000  4.255000 1.400000 ;
      RECT  4.085000  1.400000  6.245000 1.570000 ;
      RECT  4.230000  1.740000  5.255000 2.070000 ;
      RECT  4.270000  0.085000  4.600000 0.710000 ;
      RECT  4.425000  0.880000  5.160000 1.050000 ;
      RECT  4.425000  1.050000  4.770000 1.230000 ;
      RECT  4.745000  2.410000  4.915000 2.890000 ;
      RECT  4.745000  2.890000  5.690000 3.060000 ;
      RECT  4.770000  0.570000  5.160000 0.880000 ;
      RECT  4.950000  1.220000  6.245000 1.400000 ;
      RECT  5.085000  2.070000  5.255000 2.320000 ;
      RECT  5.085000  2.320000  5.350000 2.720000 ;
      RECT  5.425000  1.790000  6.115000 2.150000 ;
      RECT  5.520000  2.320000  6.585000 2.490000 ;
      RECT  5.520000  2.490000  5.690000 2.890000 ;
      RECT  5.650000  0.085000  6.245000 1.030000 ;
      RECT  5.860000  2.660000  6.110000 3.245000 ;
      RECT  5.915000  1.215000  6.245000 1.220000 ;
      RECT  6.415000  0.280000  7.660000 0.450000 ;
      RECT  6.415000  0.450000  6.585000 1.120000 ;
      RECT  6.415000  1.120000  6.960000 1.450000 ;
      RECT  6.415000  1.450000  6.585000 2.320000 ;
      RECT  6.820000  1.620000  7.320000 1.790000 ;
      RECT  6.820000  1.790000  7.070000 2.550000 ;
      RECT  6.820000  2.550000  7.930000 2.730000 ;
      RECT  6.820000  2.730000  7.470000 2.980000 ;
      RECT  6.825000  0.620000  7.320000 0.950000 ;
      RECT  7.150000  0.950000  7.320000 1.620000 ;
      RECT  7.290000  1.980000  7.660000 2.150000 ;
      RECT  7.290000  2.150000  7.590000 2.380000 ;
      RECT  7.490000  0.450000  7.660000 1.980000 ;
      RECT  7.760000  2.320000  9.470000 2.490000 ;
      RECT  7.760000  2.490000  8.880000 2.550000 ;
      RECT  7.830000  1.070000  9.890000 1.240000 ;
      RECT  7.830000  1.240000  8.145000 2.130000 ;
      RECT  8.100000  2.720000  8.430000 3.245000 ;
      RECT  8.315000  1.480000  8.730000 2.150000 ;
      RECT  8.525000  0.085000  9.360000 0.900000 ;
      RECT  8.630000  2.550000  8.880000 2.980000 ;
      RECT  9.110000  2.660000  9.440000 3.245000 ;
      RECT  9.140000  1.615000  9.470000 2.320000 ;
      RECT  9.530000  0.635000  9.890000 1.070000 ;
      RECT  9.640000  1.240000  9.890000 2.980000 ;
      RECT 10.090000  0.450000 10.420000 1.300000 ;
      RECT 10.090000  1.300000 11.125000 1.630000 ;
      RECT 10.090000  1.630000 10.450000 2.860000 ;
      RECT 10.600000  0.085000 10.930000 1.130000 ;
      RECT 10.655000  2.320000 10.985000 3.245000 ;
      RECT 11.635000  0.085000 11.885000 1.130000 ;
      RECT 11.635000  1.820000 11.885000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  1.950000  6.085000 2.120000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.950000  8.485000 2.120000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
  END
END sky130_fd_sc_ls__dfstp_2
END LIBRARY
