* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__xor3_1 A B C VGND VNB VPB VPWR X
M1000 a_27_134# a_452_288# a_416_86# VNB nshort w=420000u l=150000u
+  ad=4.987e+11p pd=4.17e+06u as=4.475e+11p ps=4.01e+06u
M1001 a_416_86# C a_1215_396# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=3.392e+11p ps=2.34e+06u
M1002 a_416_86# B a_27_134# VPB phighvt w=640000u l=150000u
+  ad=6.2055e+11p pd=4.89e+06u as=4.998e+11p ps=4.51e+06u
M1003 a_384_392# B a_84_108# VPB phighvt w=840000u l=150000u
+  ad=5.784e+11p pd=4.78e+06u as=8.756e+11p ps=5.66e+06u
M1004 a_1215_396# a_1157_298# a_416_86# VPB phighvt w=840000u l=150000u
+  ad=5.082e+11p pd=2.89e+06u as=0p ps=0u
M1005 VGND B a_452_288# VNB nshort w=740000u l=150000u
+  ad=1.3258e+12p pd=8.35e+06u as=2.035e+11p ps=2.03e+06u
M1006 a_27_134# a_452_288# a_384_392# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B a_452_288# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.3176e+12p pd=9.15e+06u as=3.304e+11p ps=2.83e+06u
M1008 a_84_108# a_452_288# a_416_86# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_384_392# B a_27_134# VNB nshort w=640000u l=150000u
+  ad=5.1415e+11p pd=4.38e+06u as=0p ps=0u
M1010 X a_1215_396# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1011 a_416_86# B a_84_108# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=6.252e+11p ps=4.99e+06u
M1012 VPWR C a_1157_298# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.528e+11p ps=2.07e+06u
M1013 a_1215_396# a_1157_298# a_384_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND C a_1157_298# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1015 X a_1215_396# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1016 VPWR a_84_108# a_27_134# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_84_108# a_27_134# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_84_108# a_452_288# a_384_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_384_392# C a_1215_396# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_84_108# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_84_108# A VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
