* NGSPICE file created from sky130_fd_sc_ls__dlymetal6s4s_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dlymetal6s4s_1 A VGND VNB VPB VPWR X
M1000 VGND X a_604_138# VNB nshort w=420000u l=150000u
+  ad=6.828e+11p pd=6.48e+06u as=1.113e+11p ps=1.37e+06u
M1001 a_209_74# a_28_138# VGND VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1002 a_785_74# a_604_138# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=1.043e+12p ps=8.92e+06u
M1003 a_785_74# a_604_138# VGND VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1004 VGND A a_28_138# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 X a_316_138# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1006 VGND a_209_74# a_316_138# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 VPWR a_209_74# a_316_138# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1008 VPWR X a_604_138# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1009 a_209_74# a_28_138# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1010 X a_316_138# VGND VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1011 VPWR A a_28_138# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
.ends

