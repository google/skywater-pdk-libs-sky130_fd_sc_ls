* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__or4b_4 A B C D_N VGND VNB VPB VPWR X
X0 a_496_392# C a_27_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_496_392# a_563_48# a_27_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_27_74# C VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 VGND a_563_48# a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 VPWR A a_116_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_563_48# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 a_27_74# a_563_48# a_496_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_27_392# B a_116_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_116_392# B a_27_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 a_563_48# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_27_392# C a_496_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X20 a_116_392# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
.ends
