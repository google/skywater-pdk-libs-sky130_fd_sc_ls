* File: sky130_fd_sc_ls__einvn_4.spice
* Created: Wed Sep  2 11:06:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__einvn_4.pex.spice"
.subckt sky130_fd_sc_ls__einvn_4  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1013 N_A_114_74#_M1013_d N_TE_B_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_281_74#_M1002_d N_A_114_74#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_281_74#_M1003_d N_A_114_74#_M1003_g N_VGND_M1002_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002.8 A=0.111 P=1.78 MULT=1
MM1009 N_A_281_74#_M1003_d N_A_114_74#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1016 N_A_281_74#_M1016_d N_A_114_74#_M1016_g N_VGND_M1009_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1000 N_A_281_74#_M1016_d N_A_M1000_g N_Z_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1004 N_A_281_74#_M1004_d N_A_M1004_g N_Z_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1073 AS=0.1036 PD=1.03 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1008 N_A_281_74#_M1004_d N_A_M1008_g N_Z_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1073 AS=0.1036 PD=1.03 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1015 N_A_281_74#_M1015_d N_A_M1015_g N_Z_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_114_74#_M1006_d N_TE_B_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1007 N_A_241_368#_M1007_d N_TE_B_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1011 N_A_241_368#_M1011_d N_TE_B_M1011_g N_VPWR_M1007_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75003 A=0.168 P=2.54 MULT=1
MM1012 N_A_241_368#_M1011_d N_TE_B_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1017 N_A_241_368#_M1017_d N_TE_B_M1017_g N_VPWR_M1012_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.6 SB=75002 A=0.168 P=2.54 MULT=1
MM1001 N_Z_M1001_d N_A_M1001_g N_A_241_368#_M1017_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1005 N_Z_M1001_d N_A_M1005_g N_A_241_368#_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1010 N_Z_M1010_d N_A_M1010_g N_A_241_368#_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75003
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1014 N_Z_M1010_d N_A_M1014_g N_A_241_368#_M1014_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.4 SB=75000.2 A=0.168 P=2.54 MULT=1
DX18_noxref VNB VPB NWDIODE A=10.5276 P=15.04
c_60 VNB 0 6.80581e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__einvn_4.pxi.spice"
*
.ends
*
*
