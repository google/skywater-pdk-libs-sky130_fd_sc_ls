* NGSPICE file created from sky130_fd_sc_ls__xnor2_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__xnor2_4 A B VGND VNB VPB VPWR Y
M1000 VPWR A a_950_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=2.77233e+12p pd=1.9e+07u as=1.6688e+12p ps=1.418e+07u
M1001 Y B a_950_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.008e+12p pd=8.52e+06u as=0p ps=0u
M1002 a_511_74# A VGND VNB nshort w=740000u l=150000u
+  ad=1.6317e+12p pd=1.477e+07u as=1.7674e+12p ps=1.293e+07u
M1003 VPWR B a_116_368# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=5.04e+11p ps=4.56e+06u
M1004 VPWR A a_950_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_511_74# a_116_368# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.662e+11p ps=4.22e+06u
M1006 VGND A a_511_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_950_368# B Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_511_74# a_116_368# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_511_74# B VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B a_511_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y a_116_368# a_511_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_74# A VGND VNB nshort w=640000u l=150000u
+  ad=5.44e+11p pd=5.54e+06u as=0p ps=0u
M1013 Y B a_950_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_116_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_116_368# A VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A a_116_368# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A a_511_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_74# B a_116_368# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.24e+11p ps=1.98e+06u
M1019 a_511_74# A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_511_74# B VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_950_368# B Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_116_368# B a_27_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_950_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_116_368# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_950_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_116_368# B VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A a_27_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y a_116_368# a_511_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND B a_511_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

