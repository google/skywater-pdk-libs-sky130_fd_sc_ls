* File: sky130_fd_sc_ls__clkdlyinv5sd2_1.pxi.spice
* Created: Fri Aug 28 13:10:11 2020
* 
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A N_A_M1007_g N_A_c_78_n N_A_c_82_n
+ N_A_M1008_g A A N_A_c_80_n PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A_28_74# N_A_28_74#_M1007_s
+ N_A_28_74#_M1008_s N_A_28_74#_M1009_g N_A_28_74#_M1006_g N_A_28_74#_c_117_n
+ N_A_28_74#_c_123_n N_A_28_74#_c_124_n N_A_28_74#_c_134_n N_A_28_74#_c_118_n
+ N_A_28_74#_c_119_n N_A_28_74#_c_120_n N_A_28_74#_c_121_n
+ PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A_28_74#
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A_288_74# N_A_288_74#_M1006_d
+ N_A_288_74#_M1009_d N_A_288_74#_M1001_g N_A_288_74#_M1000_g
+ N_A_288_74#_c_179_n N_A_288_74#_c_180_n N_A_288_74#_c_181_n
+ N_A_288_74#_c_186_n N_A_288_74#_c_182_n N_A_288_74#_c_183_n
+ PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A_288_74#
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A_549_74# N_A_549_74#_M1000_d
+ N_A_549_74#_M1001_d N_A_549_74#_M1004_g N_A_549_74#_M1003_g
+ N_A_549_74#_c_222_n N_A_549_74#_c_223_n N_A_549_74#_c_224_n
+ N_A_549_74#_c_225_n N_A_549_74#_c_226_n
+ PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A_549_74#
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A_682_74# N_A_682_74#_M1003_s
+ N_A_682_74#_M1004_s N_A_682_74#_M1005_g N_A_682_74#_c_269_n
+ N_A_682_74#_M1002_g N_A_682_74#_c_270_n N_A_682_74#_c_277_n
+ N_A_682_74#_c_271_n N_A_682_74#_c_272_n N_A_682_74#_c_273_n
+ N_A_682_74#_c_274_n N_A_682_74#_c_275_n
+ PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%A_682_74#
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%VPWR N_VPWR_M1008_d N_VPWR_M1001_s
+ N_VPWR_M1004_d N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_327_n VPWR
+ N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_331_n N_VPWR_c_324_n
+ N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n VPWR
+ PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%VPWR
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%Y N_Y_M1005_d N_Y_M1002_d Y Y Y Y Y Y Y Y
+ PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%Y
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%VGND N_VGND_M1007_d N_VGND_M1000_s
+ N_VGND_M1003_d N_VGND_c_391_n N_VGND_c_392_n N_VGND_c_393_n VGND
+ N_VGND_c_394_n N_VGND_c_395_n N_VGND_c_396_n N_VGND_c_397_n N_VGND_c_398_n
+ N_VGND_c_399_n N_VGND_c_400_n N_VGND_c_401_n VGND
+ PM_SKY130_FD_SC_LS__CLKDLYINV5SD2_1%VGND
cc_1 VNB N_A_M1007_g 0.0470899f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.58
cc_2 VNB N_A_c_78_n 0.00974989f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.675
cc_3 VNB A 0.026734f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A_c_80_n 0.0363883f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_5 VNB N_A_28_74#_M1009_g 0.0139918f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_6 VNB N_A_28_74#_M1006_g 0.0379459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_28_74#_c_117_n 0.0226356f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.19
cc_8 VNB N_A_28_74#_c_118_n 0.0206633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_28_74#_c_119_n 0.0121635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_28_74#_c_120_n 0.00294396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_28_74#_c_121_n 0.0477075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_288_74#_M1001_g 0.0186271f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_13 VNB N_A_288_74#_M1000_g 0.049015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_288_74#_c_179_n 0.0268697f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.19
cc_15 VNB N_A_288_74#_c_180_n 0.00978917f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.355
cc_16 VNB N_A_288_74#_c_181_n 0.0255344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_288_74#_c_182_n 0.00614775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_288_74#_c_183_n 0.0633733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_549_74#_M1004_g 0.0158734f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_20 VNB N_A_549_74#_M1003_g 0.0437533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_549_74#_c_222_n 0.0155677f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.19
cc_22 VNB N_A_549_74#_c_223_n 0.0111173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_549_74#_c_224_n 0.0372738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_549_74#_c_225_n 0.00227058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_549_74#_c_226_n 0.0525203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_682_74#_M1005_g 0.0444659f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_27 VNB N_A_682_74#_c_269_n 0.0391593f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_28 VNB N_A_682_74#_c_270_n 0.00814692f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_29 VNB N_A_682_74#_c_271_n 0.00612199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_682_74#_c_272_n 0.00422437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_682_74#_c_273_n 0.0258925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_682_74#_c_274_n 0.0067964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_682_74#_c_275_n 0.00272046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_324_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB Y 0.0204118f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_36 VNB Y 0.0466962f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_37 VNB N_VGND_c_391_n 0.00987431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_392_n 0.0149241f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_39 VNB N_VGND_c_393_n 0.00662038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_394_n 0.0180717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_395_n 0.0296852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_396_n 0.0621707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_397_n 0.0189455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_398_n 0.344385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_399_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_400_n 0.00673217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_401_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VPB N_A_c_78_n 9.82004e-19 $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.675
cc_49 VPB N_A_c_82_n 0.0289243f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_50 VPB A 0.0107514f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_51 VPB N_A_28_74#_M1009_g 0.0409302f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_52 VPB N_A_28_74#_c_123_n 0.0079884f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.295
cc_53 VPB N_A_28_74#_c_124_n 0.0205617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_28_74#_c_120_n 0.00325766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_288_74#_M1001_g 0.0500614f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_56 VPB N_A_288_74#_c_180_n 0.02236f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.355
cc_57 VPB N_A_288_74#_c_186_n 0.00306613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_549_74#_M1004_g 0.0440843f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_59 VPB N_A_549_74#_c_223_n 0.0106835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_682_74#_c_269_n 0.0254953f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_61 VPB N_A_682_74#_c_277_n 0.00967761f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_682_74#_c_271_n 0.0175672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_682_74#_c_272_n 0.00141791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_325_n 0.0101831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_326_n 0.0260677f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.355
cc_66 VPB N_VPWR_c_327_n 0.00777218f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.355
cc_67 VPB N_VPWR_c_328_n 0.018958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_329_n 0.0298867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_330_n 0.0624644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_331_n 0.0184442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_324_n 0.12435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_333_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_334_n 0.00670627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_335_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB Y 0.0121098f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_76 VPB Y 0.0526708f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_77 A N_A_28_74#_M1008_s 0.00256075f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_78 N_A_c_78_n N_A_28_74#_M1009_g 0.00320655f $X=0.495 $Y=1.675 $X2=0 $Y2=0
cc_79 N_A_c_82_n N_A_28_74#_M1009_g 0.0135624f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_80 A N_A_28_74#_M1009_g 0.0011323f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A_c_80_n N_A_28_74#_M1009_g 0.00126282f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_82 N_A_M1007_g N_A_28_74#_M1006_g 0.00808739f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_83 N_A_M1007_g N_A_28_74#_c_117_n 0.0127782f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_84 A N_A_28_74#_c_123_n 0.0237727f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A_c_82_n N_A_28_74#_c_134_n 0.0144812f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_86 A N_A_28_74#_c_134_n 0.0197054f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_87 N_A_c_80_n N_A_28_74#_c_134_n 6.00585e-19 $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_88 N_A_M1007_g N_A_28_74#_c_118_n 0.0120856f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_89 A N_A_28_74#_c_118_n 0.0251751f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_90 N_A_c_80_n N_A_28_74#_c_118_n 0.00146806f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_91 N_A_M1007_g N_A_28_74#_c_119_n 0.00415005f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_92 A N_A_28_74#_c_119_n 0.0289843f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_93 N_A_M1007_g N_A_28_74#_c_120_n 0.0025292f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_94 N_A_c_78_n N_A_28_74#_c_120_n 8.04262e-19 $X=0.495 $Y=1.675 $X2=0 $Y2=0
cc_95 N_A_c_82_n N_A_28_74#_c_120_n 0.00370461f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_96 A N_A_28_74#_c_120_n 0.0427383f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A_c_80_n N_A_28_74#_c_120_n 0.00141272f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_98 N_A_M1007_g N_A_28_74#_c_121_n 0.0021171f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_99 A N_A_28_74#_c_121_n 0.00102763f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_100 N_A_c_80_n N_A_28_74#_c_121_n 0.0170907f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_101 A N_VPWR_M1008_d 0.00135779f $X=0.155 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_102 N_A_c_82_n N_VPWR_c_325_n 0.00426168f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A_c_82_n N_VPWR_c_328_n 0.00461464f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_104 N_A_c_82_n N_VPWR_c_324_n 0.00913361f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A_M1007_g N_VGND_c_391_n 0.00293875f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_106 N_A_M1007_g N_VGND_c_394_n 0.00456766f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_107 N_A_M1007_g N_VGND_c_398_n 0.00456437f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_108 N_A_28_74#_M1006_g N_A_288_74#_c_179_n 0.0110261f $X=1.35 $Y=0.58 $X2=0
+ $Y2=0
cc_109 N_A_28_74#_c_118_n N_A_288_74#_c_179_n 0.0164122f $X=0.975 $Y=0.92 $X2=0
+ $Y2=0
cc_110 N_A_28_74#_c_120_n N_A_288_74#_c_179_n 0.00916028f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_111 N_A_28_74#_c_121_n N_A_288_74#_c_179_n 2.87835e-19 $X=1.35 $Y=1.295 $X2=0
+ $Y2=0
cc_112 N_A_28_74#_M1009_g N_A_288_74#_c_180_n 0.0124318f $X=1.32 $Y=2.46 $X2=0
+ $Y2=0
cc_113 N_A_28_74#_c_120_n N_A_288_74#_c_180_n 0.0406706f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_114 N_A_28_74#_M1009_g N_A_288_74#_c_186_n 0.00707225f $X=1.32 $Y=2.46 $X2=0
+ $Y2=0
cc_115 N_A_28_74#_c_120_n N_A_288_74#_c_182_n 0.0277877f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_116 N_A_28_74#_c_121_n N_A_288_74#_c_182_n 0.00984463f $X=1.35 $Y=1.295 $X2=0
+ $Y2=0
cc_117 N_A_28_74#_c_134_n N_VPWR_M1008_d 0.0250817f $X=0.975 $Y=2.117 $X2=-0.19
+ $Y2=-0.245
cc_118 N_A_28_74#_c_120_n N_VPWR_M1008_d 0.0012063f $X=1.14 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_119 N_A_28_74#_M1009_g N_VPWR_c_325_n 0.0104916f $X=1.32 $Y=2.46 $X2=0 $Y2=0
cc_120 N_A_28_74#_c_134_n N_VPWR_c_325_n 0.0220956f $X=0.975 $Y=2.117 $X2=0
+ $Y2=0
cc_121 N_A_28_74#_M1009_g N_VPWR_c_326_n 0.00458004f $X=1.32 $Y=2.46 $X2=0 $Y2=0
cc_122 N_A_28_74#_c_124_n N_VPWR_c_328_n 0.00593336f $X=0.265 $Y=2.56 $X2=0
+ $Y2=0
cc_123 N_A_28_74#_M1009_g N_VPWR_c_329_n 0.00738282f $X=1.32 $Y=2.46 $X2=0 $Y2=0
cc_124 N_A_28_74#_M1009_g N_VPWR_c_324_n 0.014148f $X=1.32 $Y=2.46 $X2=0 $Y2=0
cc_125 N_A_28_74#_c_124_n N_VPWR_c_324_n 0.00940928f $X=0.265 $Y=2.56 $X2=0
+ $Y2=0
cc_126 N_A_28_74#_M1006_g N_VGND_c_391_n 0.00513169f $X=1.35 $Y=0.58 $X2=0 $Y2=0
cc_127 N_A_28_74#_c_117_n N_VGND_c_391_n 0.0151665f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_128 N_A_28_74#_c_118_n N_VGND_c_391_n 0.0255952f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_129 N_A_28_74#_M1006_g N_VGND_c_392_n 0.0024778f $X=1.35 $Y=0.58 $X2=0 $Y2=0
cc_130 N_A_28_74#_c_117_n N_VGND_c_394_n 0.0170785f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_131 N_A_28_74#_M1006_g N_VGND_c_395_n 0.00553757f $X=1.35 $Y=0.58 $X2=0 $Y2=0
cc_132 N_A_28_74#_M1006_g N_VGND_c_398_n 0.00962875f $X=1.35 $Y=0.58 $X2=0 $Y2=0
cc_133 N_A_28_74#_c_117_n N_VGND_c_398_n 0.0118627f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_134 N_A_28_74#_c_118_n N_VGND_c_398_n 0.0213669f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_135 N_A_288_74#_M1000_g N_A_549_74#_c_222_n 0.0165136f $X=2.655 $Y=0.58 $X2=0
+ $Y2=0
cc_136 N_A_288_74#_c_181_n N_A_549_74#_c_222_n 0.00419423f $X=2.425 $Y=1.305
+ $X2=0 $Y2=0
cc_137 N_A_288_74#_c_181_n N_A_549_74#_c_223_n 0.00419423f $X=2.425 $Y=1.305
+ $X2=0 $Y2=0
cc_138 N_A_288_74#_c_183_n N_A_549_74#_c_223_n 0.0228612f $X=2.655 $Y=1.305
+ $X2=0 $Y2=0
cc_139 N_A_288_74#_c_181_n N_A_549_74#_c_225_n 0.0101411f $X=2.425 $Y=1.305
+ $X2=0 $Y2=0
cc_140 N_A_288_74#_c_183_n N_A_549_74#_c_225_n 0.00534783f $X=2.655 $Y=1.305
+ $X2=0 $Y2=0
cc_141 N_A_288_74#_c_186_n N_VPWR_c_325_n 0.00825858f $X=1.58 $Y=2.815 $X2=0
+ $Y2=0
cc_142 N_A_288_74#_M1001_g N_VPWR_c_326_n 0.0290944f $X=2.62 $Y=2.46 $X2=0 $Y2=0
cc_143 N_A_288_74#_c_180_n N_VPWR_c_326_n 0.0793707f $X=1.58 $Y=2.105 $X2=0
+ $Y2=0
cc_144 N_A_288_74#_c_181_n N_VPWR_c_326_n 0.0151215f $X=2.425 $Y=1.305 $X2=0
+ $Y2=0
cc_145 N_A_288_74#_c_183_n N_VPWR_c_326_n 3.64176e-19 $X=2.655 $Y=1.305 $X2=0
+ $Y2=0
cc_146 N_A_288_74#_c_186_n N_VPWR_c_329_n 0.00976575f $X=1.58 $Y=2.815 $X2=0
+ $Y2=0
cc_147 N_A_288_74#_M1001_g N_VPWR_c_330_n 0.00769107f $X=2.62 $Y=2.46 $X2=0
+ $Y2=0
cc_148 N_A_288_74#_M1001_g N_VPWR_c_324_n 0.0152163f $X=2.62 $Y=2.46 $X2=0 $Y2=0
cc_149 N_A_288_74#_c_186_n N_VPWR_c_324_n 0.0112865f $X=1.58 $Y=2.815 $X2=0
+ $Y2=0
cc_150 N_A_288_74#_c_179_n N_VGND_c_391_n 0.00689121f $X=1.58 $Y=0.58 $X2=0
+ $Y2=0
cc_151 N_A_288_74#_M1000_g N_VGND_c_392_n 0.012646f $X=2.655 $Y=0.58 $X2=0 $Y2=0
cc_152 N_A_288_74#_c_179_n N_VGND_c_392_n 0.0326862f $X=1.58 $Y=0.58 $X2=0 $Y2=0
cc_153 N_A_288_74#_c_181_n N_VGND_c_392_n 0.0165176f $X=2.425 $Y=1.305 $X2=0
+ $Y2=0
cc_154 N_A_288_74#_c_183_n N_VGND_c_392_n 3.84795e-19 $X=2.655 $Y=1.305 $X2=0
+ $Y2=0
cc_155 N_A_288_74#_c_179_n N_VGND_c_395_n 0.0132196f $X=1.58 $Y=0.58 $X2=0 $Y2=0
cc_156 N_A_288_74#_M1000_g N_VGND_c_396_n 0.00553757f $X=2.655 $Y=0.58 $X2=0
+ $Y2=0
cc_157 N_A_288_74#_M1000_g N_VGND_c_398_n 0.0110002f $X=2.655 $Y=0.58 $X2=0
+ $Y2=0
cc_158 N_A_288_74#_c_179_n N_VGND_c_398_n 0.00920999f $X=1.58 $Y=0.58 $X2=0
+ $Y2=0
cc_159 N_A_549_74#_M1003_g N_A_682_74#_M1005_g 0.0193595f $X=4.085 $Y=0.58 $X2=0
+ $Y2=0
cc_160 N_A_549_74#_M1004_g N_A_682_74#_c_269_n 0.0192848f $X=4.045 $Y=2.46 $X2=0
+ $Y2=0
cc_161 N_A_549_74#_c_224_n N_A_682_74#_c_269_n 2.99954e-19 $X=3.84 $Y=1.305
+ $X2=0 $Y2=0
cc_162 N_A_549_74#_c_226_n N_A_682_74#_c_269_n 0.0130085f $X=4.045 $Y=1.305
+ $X2=0 $Y2=0
cc_163 N_A_549_74#_M1003_g N_A_682_74#_c_270_n 0.0127986f $X=4.085 $Y=0.58 $X2=0
+ $Y2=0
cc_164 N_A_549_74#_c_222_n N_A_682_74#_c_270_n 0.0198272f $X=2.885 $Y=0.58 $X2=0
+ $Y2=0
cc_165 N_A_549_74#_M1004_g N_A_682_74#_c_277_n 0.0313626f $X=4.045 $Y=2.46 $X2=0
+ $Y2=0
cc_166 N_A_549_74#_c_223_n N_A_682_74#_c_277_n 0.046582f $X=2.885 $Y=2.105 $X2=0
+ $Y2=0
cc_167 N_A_549_74#_M1004_g N_A_682_74#_c_271_n 0.0265909f $X=4.045 $Y=2.46 $X2=0
+ $Y2=0
cc_168 N_A_549_74#_c_224_n N_A_682_74#_c_271_n 0.0247324f $X=3.84 $Y=1.305 $X2=0
+ $Y2=0
cc_169 N_A_549_74#_c_226_n N_A_682_74#_c_271_n 0.00629507f $X=4.045 $Y=1.305
+ $X2=0 $Y2=0
cc_170 N_A_549_74#_c_223_n N_A_682_74#_c_272_n 0.0073655f $X=2.885 $Y=2.105
+ $X2=0 $Y2=0
cc_171 N_A_549_74#_c_224_n N_A_682_74#_c_272_n 0.0202705f $X=3.84 $Y=1.305 $X2=0
+ $Y2=0
cc_172 N_A_549_74#_M1003_g N_A_682_74#_c_273_n 0.021524f $X=4.085 $Y=0.58 $X2=0
+ $Y2=0
cc_173 N_A_549_74#_c_224_n N_A_682_74#_c_273_n 0.0217376f $X=3.84 $Y=1.305 $X2=0
+ $Y2=0
cc_174 N_A_549_74#_c_226_n N_A_682_74#_c_273_n 0.0075907f $X=4.045 $Y=1.305
+ $X2=0 $Y2=0
cc_175 N_A_549_74#_c_222_n N_A_682_74#_c_274_n 0.0079307f $X=2.885 $Y=0.58 $X2=0
+ $Y2=0
cc_176 N_A_549_74#_c_224_n N_A_682_74#_c_274_n 0.0276549f $X=3.84 $Y=1.305 $X2=0
+ $Y2=0
cc_177 N_A_549_74#_c_226_n N_A_682_74#_c_274_n 7.67879e-19 $X=4.045 $Y=1.305
+ $X2=0 $Y2=0
cc_178 N_A_549_74#_M1003_g N_A_682_74#_c_275_n 0.00400412f $X=4.085 $Y=0.58
+ $X2=0 $Y2=0
cc_179 N_A_549_74#_c_224_n N_A_682_74#_c_275_n 0.00545692f $X=3.84 $Y=1.305
+ $X2=0 $Y2=0
cc_180 N_A_549_74#_c_226_n N_A_682_74#_c_275_n 0.00150236f $X=4.045 $Y=1.305
+ $X2=0 $Y2=0
cc_181 N_A_549_74#_c_223_n N_VPWR_c_326_n 0.0186028f $X=2.885 $Y=2.105 $X2=0
+ $Y2=0
cc_182 N_A_549_74#_M1004_g N_VPWR_c_327_n 0.0185609f $X=4.045 $Y=2.46 $X2=0
+ $Y2=0
cc_183 N_A_549_74#_M1004_g N_VPWR_c_330_n 0.00769107f $X=4.045 $Y=2.46 $X2=0
+ $Y2=0
cc_184 N_A_549_74#_c_223_n N_VPWR_c_330_n 0.00749631f $X=2.885 $Y=2.105 $X2=0
+ $Y2=0
cc_185 N_A_549_74#_M1004_g N_VPWR_c_324_n 0.015182f $X=4.045 $Y=2.46 $X2=0 $Y2=0
cc_186 N_A_549_74#_c_223_n N_VPWR_c_324_n 0.0062048f $X=2.885 $Y=2.105 $X2=0
+ $Y2=0
cc_187 N_A_549_74#_M1003_g N_VGND_c_393_n 0.00781382f $X=4.085 $Y=0.58 $X2=0
+ $Y2=0
cc_188 N_A_549_74#_M1003_g N_VGND_c_396_n 0.00553757f $X=4.085 $Y=0.58 $X2=0
+ $Y2=0
cc_189 N_A_549_74#_c_222_n N_VGND_c_396_n 0.00573605f $X=2.885 $Y=0.58 $X2=0
+ $Y2=0
cc_190 N_A_549_74#_M1003_g N_VGND_c_398_n 0.0109653f $X=4.085 $Y=0.58 $X2=0
+ $Y2=0
cc_191 N_A_549_74#_c_222_n N_VGND_c_398_n 0.00594877f $X=2.885 $Y=0.58 $X2=0
+ $Y2=0
cc_192 N_A_682_74#_c_269_n N_VPWR_c_327_n 0.0163879f $X=4.72 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_A_682_74#_c_277_n N_VPWR_c_327_n 0.0299317f $X=3.535 $Y=2.105 $X2=0
+ $Y2=0
cc_194 N_A_682_74#_c_271_n N_VPWR_c_327_n 0.0255637f $X=4.53 $Y=1.645 $X2=0
+ $Y2=0
cc_195 N_A_682_74#_c_277_n N_VPWR_c_330_n 0.0106198f $X=3.535 $Y=2.105 $X2=0
+ $Y2=0
cc_196 N_A_682_74#_c_269_n N_VPWR_c_331_n 0.00413917f $X=4.72 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_A_682_74#_c_269_n N_VPWR_c_324_n 0.00821389f $X=4.72 $Y=1.765 $X2=0
+ $Y2=0
cc_198 N_A_682_74#_c_277_n N_VPWR_c_324_n 0.00879013f $X=3.535 $Y=2.105 $X2=0
+ $Y2=0
cc_199 N_A_682_74#_M1005_g Y 8.21909e-19 $X=4.71 $Y=0.58 $X2=0 $Y2=0
cc_200 N_A_682_74#_M1005_g Y 0.0124475f $X=4.71 $Y=0.58 $X2=0 $Y2=0
cc_201 N_A_682_74#_c_269_n Y 0.0163621f $X=4.72 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A_682_74#_c_271_n Y 0.0140324f $X=4.53 $Y=1.645 $X2=0 $Y2=0
cc_203 N_A_682_74#_c_273_n Y 0.0133247f $X=4.53 $Y=0.965 $X2=0 $Y2=0
cc_204 N_A_682_74#_c_275_n Y 0.0384675f $X=4.67 $Y=1.46 $X2=0 $Y2=0
cc_205 N_A_682_74#_c_269_n Y 0.00229934f $X=4.72 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A_682_74#_M1005_g N_VGND_c_393_n 0.0112059f $X=4.71 $Y=0.58 $X2=0 $Y2=0
cc_207 N_A_682_74#_c_269_n N_VGND_c_393_n 3.24916e-19 $X=4.72 $Y=1.765 $X2=0
+ $Y2=0
cc_208 N_A_682_74#_c_270_n N_VGND_c_393_n 0.00806009f $X=3.535 $Y=0.565 $X2=0
+ $Y2=0
cc_209 N_A_682_74#_c_273_n N_VGND_c_393_n 0.0218411f $X=4.53 $Y=0.965 $X2=0
+ $Y2=0
cc_210 N_A_682_74#_c_270_n N_VGND_c_396_n 0.0118185f $X=3.535 $Y=0.565 $X2=0
+ $Y2=0
cc_211 N_A_682_74#_M1005_g N_VGND_c_397_n 0.00383152f $X=4.71 $Y=0.58 $X2=0
+ $Y2=0
cc_212 N_A_682_74#_M1005_g N_VGND_c_398_n 0.00761428f $X=4.71 $Y=0.58 $X2=0
+ $Y2=0
cc_213 N_A_682_74#_c_270_n N_VGND_c_398_n 0.0117223f $X=3.535 $Y=0.565 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_327_n Y 0.0476994f $X=4.495 $Y=1.985 $X2=0 $Y2=0
cc_215 N_VPWR_c_331_n Y 0.0234396f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_216 N_VPWR_c_324_n Y 0.0138183f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_217 Y N_VGND_c_393_n 0.0124097f $X=4.95 $Y=0.47 $X2=0 $Y2=0
cc_218 Y N_VGND_c_397_n 0.0155069f $X=4.95 $Y=0.47 $X2=0 $Y2=0
cc_219 Y N_VGND_c_398_n 0.013122f $X=4.95 $Y=0.47 $X2=0 $Y2=0
