* File: sky130_fd_sc_ls__decaphe_2.pxi.spice
* Created: Wed Sep  2 10:59:40 2020
* 
x_PM_SKY130_FD_SC_LS__DECAPHE_2%VGND N_VGND_M1000_g N_VGND_c_14_n N_VGND_c_15_n
+ VGND N_VGND_c_16_n N_VGND_c_17_n N_VGND_c_18_n
+ PM_SKY130_FD_SC_LS__DECAPHE_2%VGND
x_PM_SKY130_FD_SC_LS__DECAPHE_2%VPWR N_VPWR_M1000_s N_VPWR_c_25_n VPWR
+ N_VPWR_c_27_n VPWR PM_SKY130_FD_SC_LS__DECAPHE_2%VPWR
cc_1 VNB N_VGND_M1000_g 0.0027366f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.467
cc_2 VNB N_VGND_c_14_n 0.0123177f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=0.085
cc_3 VNB N_VGND_c_15_n 0.112553f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_VGND_c_16_n 0.0669607f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.465
cc_5 VNB N_VGND_c_17_n 0.0177361f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0
cc_6 VNB N_VGND_c_18_n 0.103415f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0
cc_7 VNB VPWR 0.0442671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VPB N_VGND_M1000_g 0.0346968f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=2.467
cc_9 VPB N_VGND_c_15_n 0.0034656f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_10 VPB N_VPWR_c_25_n 0.113436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_11 VPB VPWR 0.0423048f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_12 VPB N_VPWR_c_27_n 0.021794f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0
cc_13 N_VGND_M1000_g N_VPWR_c_25_n 0.0434328f $X=0.48 $Y=2.467 $X2=0 $Y2=0
cc_14 N_VGND_c_15_n N_VPWR_c_25_n 0.0321444f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_15 N_VGND_c_16_n N_VPWR_c_25_n 0.00187508f $X=0.48 $Y=1.465 $X2=0 $Y2=0
