* File: sky130_fd_sc_ls__maj3_4.pxi.spice
* Created: Wed Sep  2 11:10:03 2020
* 
x_PM_SKY130_FD_SC_LS__MAJ3_4%B N_B_c_152_n N_B_M1011_g N_B_c_144_n N_B_M1016_g
+ N_B_c_153_n N_B_M1022_g N_B_c_145_n N_B_M1023_g N_B_c_154_n N_B_M1001_g
+ N_B_c_146_n N_B_M1024_g N_B_c_147_n N_B_M1030_g N_B_c_155_n N_B_M1005_g
+ N_B_c_156_n N_B_c_198_p B B N_B_c_149_n N_B_c_150_n N_B_c_151_n
+ PM_SKY130_FD_SC_LS__MAJ3_4%B
x_PM_SKY130_FD_SC_LS__MAJ3_4%A N_A_M1013_g N_A_c_259_n N_A_c_275_n N_A_M1014_g
+ N_A_c_260_n N_A_c_261_n N_A_c_262_n N_A_M1029_g N_A_M1019_g N_A_c_264_n
+ N_A_M1006_g N_A_M1004_g N_A_c_266_n N_A_c_267_n N_A_c_268_n N_A_c_279_n
+ N_A_M1028_g N_A_M1009_g N_A_c_270_n N_A_c_271_n N_A_c_280_n N_A_c_272_n A
+ PM_SKY130_FD_SC_LS__MAJ3_4%A
x_PM_SKY130_FD_SC_LS__MAJ3_4%C N_C_c_417_n N_C_c_418_n N_C_c_432_n N_C_M1012_g
+ N_C_M1007_g N_C_c_420_n N_C_c_421_n N_C_c_422_n N_C_M1027_g N_C_M1017_g
+ N_C_c_434_n N_C_M1015_g N_C_M1002_g N_C_c_435_n N_C_M1018_g N_C_M1008_g
+ N_C_c_426_n N_C_c_427_n N_C_c_428_n C N_C_c_429_n N_C_c_430_n
+ PM_SKY130_FD_SC_LS__MAJ3_4%C
x_PM_SKY130_FD_SC_LS__MAJ3_4%A_219_392# N_A_219_392#_M1016_s
+ N_A_219_392#_M1024_s N_A_219_392#_M1002_d N_A_219_392#_M1011_d
+ N_A_219_392#_M1001_d N_A_219_392#_M1015_d N_A_219_392#_c_567_n
+ N_A_219_392#_M1000_g N_A_219_392#_c_556_n N_A_219_392#_M1020_g
+ N_A_219_392#_c_568_n N_A_219_392#_M1003_g N_A_219_392#_c_557_n
+ N_A_219_392#_M1021_g N_A_219_392#_c_569_n N_A_219_392#_M1010_g
+ N_A_219_392#_c_558_n N_A_219_392#_M1025_g N_A_219_392#_c_570_n
+ N_A_219_392#_M1026_g N_A_219_392#_c_559_n N_A_219_392#_M1031_g
+ N_A_219_392#_c_560_n N_A_219_392#_c_561_n N_A_219_392#_c_572_n
+ N_A_219_392#_c_590_n N_A_219_392#_c_687_p N_A_219_392#_c_591_n
+ N_A_219_392#_c_594_n N_A_219_392#_c_595_n N_A_219_392#_c_596_n
+ N_A_219_392#_c_562_n N_A_219_392#_c_573_n N_A_219_392#_c_563_n
+ N_A_219_392#_c_597_n N_A_219_392#_c_598_n N_A_219_392#_c_564_n
+ N_A_219_392#_c_627_n N_A_219_392#_c_565_n N_A_219_392#_c_566_n
+ PM_SKY130_FD_SC_LS__MAJ3_4%A_219_392#
x_PM_SKY130_FD_SC_LS__MAJ3_4%VPWR N_VPWR_M1014_s N_VPWR_M1029_s N_VPWR_M1027_d
+ N_VPWR_M1028_s N_VPWR_M1003_d N_VPWR_M1026_d N_VPWR_c_777_n N_VPWR_c_778_n
+ N_VPWR_c_779_n N_VPWR_c_780_n N_VPWR_c_781_n N_VPWR_c_782_n N_VPWR_c_783_n
+ N_VPWR_c_784_n N_VPWR_c_785_n VPWR N_VPWR_c_786_n N_VPWR_c_787_n
+ N_VPWR_c_788_n N_VPWR_c_789_n N_VPWR_c_790_n N_VPWR_c_791_n N_VPWR_c_792_n
+ N_VPWR_c_793_n N_VPWR_c_776_n PM_SKY130_FD_SC_LS__MAJ3_4%VPWR
x_PM_SKY130_FD_SC_LS__MAJ3_4%A_119_392# N_A_119_392#_M1014_d
+ N_A_119_392#_M1022_s N_A_119_392#_c_894_n N_A_119_392#_c_888_n
+ N_A_119_392#_c_889_n N_A_119_392#_c_892_n
+ PM_SKY130_FD_SC_LS__MAJ3_4%A_119_392#
x_PM_SKY130_FD_SC_LS__MAJ3_4%A_501_392# N_A_501_392#_M1012_s
+ N_A_501_392#_M1005_s N_A_501_392#_c_916_n N_A_501_392#_c_914_n
+ N_A_501_392#_c_915_n N_A_501_392#_c_926_n
+ PM_SKY130_FD_SC_LS__MAJ3_4%A_501_392#
x_PM_SKY130_FD_SC_LS__MAJ3_4%A_905_392# N_A_905_392#_M1006_d
+ N_A_905_392#_M1018_s N_A_905_392#_c_945_n N_A_905_392#_c_941_n
+ N_A_905_392#_c_942_n PM_SKY130_FD_SC_LS__MAJ3_4%A_905_392#
x_PM_SKY130_FD_SC_LS__MAJ3_4%X N_X_M1020_s N_X_M1025_s N_X_M1000_s N_X_M1010_s
+ N_X_c_973_n N_X_c_970_n N_X_c_966_n N_X_c_967_n N_X_c_986_n N_X_c_988_n
+ N_X_c_971_n N_X_c_972_n N_X_c_968_n N_X_c_999_n N_X_c_1015_n X
+ PM_SKY130_FD_SC_LS__MAJ3_4%X
x_PM_SKY130_FD_SC_LS__MAJ3_4%VGND N_VGND_M1013_d N_VGND_M1019_d N_VGND_M1017_d
+ N_VGND_M1009_s N_VGND_M1021_d N_VGND_M1031_d N_VGND_c_1025_n N_VGND_c_1026_n
+ N_VGND_c_1027_n N_VGND_c_1028_n N_VGND_c_1029_n N_VGND_c_1030_n
+ N_VGND_c_1031_n N_VGND_c_1032_n VGND N_VGND_c_1033_n N_VGND_c_1034_n
+ N_VGND_c_1035_n N_VGND_c_1036_n N_VGND_c_1037_n N_VGND_c_1038_n
+ N_VGND_c_1039_n N_VGND_c_1040_n N_VGND_c_1041_n N_VGND_c_1042_n
+ PM_SKY130_FD_SC_LS__MAJ3_4%VGND
x_PM_SKY130_FD_SC_LS__MAJ3_4%A_114_125# N_A_114_125#_M1013_s
+ N_A_114_125#_M1023_d N_A_114_125#_c_1119_n N_A_114_125#_c_1120_n
+ N_A_114_125#_c_1121_n PM_SKY130_FD_SC_LS__MAJ3_4%A_114_125#
x_PM_SKY130_FD_SC_LS__MAJ3_4%A_504_125# N_A_504_125#_M1007_s
+ N_A_504_125#_M1030_d N_A_504_125#_c_1145_n N_A_504_125#_c_1146_n
+ N_A_504_125#_c_1147_n N_A_504_125#_c_1148_n
+ PM_SKY130_FD_SC_LS__MAJ3_4%A_504_125#
x_PM_SKY130_FD_SC_LS__MAJ3_4%A_906_78# N_A_906_78#_M1004_d N_A_906_78#_M1008_s
+ N_A_906_78#_c_1179_n N_A_906_78#_c_1180_n N_A_906_78#_c_1181_n
+ PM_SKY130_FD_SC_LS__MAJ3_4%A_906_78#
cc_1 VNB N_B_c_144_n 0.0157719f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.375
cc_2 VNB N_B_c_145_n 0.0149548f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.375
cc_3 VNB N_B_c_146_n 0.0137321f $X=-0.19 $Y=-0.245 $X2=2.935 $Y2=1.375
cc_4 VNB N_B_c_147_n 0.0160268f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=1.375
cc_5 VNB B 0.00439542f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=1.21
cc_6 VNB N_B_c_149_n 0.0332199f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.63
cc_7 VNB N_B_c_150_n 0.0346107f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=1.63
cc_8 VNB N_B_c_151_n 0.0109019f $X=-0.19 $Y=-0.245 $X2=2.525 $Y2=1.417
cc_9 VNB N_A_M1013_g 0.0308567f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.375
cc_10 VNB N_A_c_259_n 0.0149597f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.945
cc_11 VNB N_A_c_260_n 0.101661f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.375
cc_12 VNB N_A_c_261_n 0.011606f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.945
cc_13 VNB N_A_c_262_n 0.0156618f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.945
cc_14 VNB N_A_M1019_g 0.0327977f $X=-0.19 $Y=-0.245 $X2=2.935 $Y2=0.945
cc_15 VNB N_A_c_264_n 0.0182643f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=1.375
cc_16 VNB N_A_M1004_g 0.0329262f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=1.3
cc_17 VNB N_A_c_266_n 0.0964178f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=1.54
cc_18 VNB N_A_c_267_n 0.0100101f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=1.54
cc_19 VNB N_A_c_268_n 0.00855675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_M1009_g 0.0245517f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.63
cc_21 VNB N_A_c_270_n 0.0162773f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=1.63
cc_22 VNB N_A_c_271_n 0.00852526f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.63
cc_23 VNB N_A_c_272_n 0.00166672f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.54
cc_24 VNB A 0.00579074f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=1.417
cc_25 VNB N_C_c_417_n 0.00583798f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.885
cc_26 VNB N_C_c_418_n 0.0124141f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=2.46
cc_27 VNB N_C_M1007_g 0.0255161f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.46
cc_28 VNB N_C_c_420_n 0.101029f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.375
cc_29 VNB N_C_c_421_n 0.00961946f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.945
cc_30 VNB N_C_c_422_n 0.0246882f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.945
cc_31 VNB N_C_M1017_g 0.0226241f $X=-0.19 $Y=-0.245 $X2=2.935 $Y2=0.945
cc_32 VNB N_C_M1002_g 0.0212185f $X=-0.19 $Y=-0.245 $X2=3.38 $Y2=2.46
cc_33 VNB N_C_M1008_g 0.0187456f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=1.215
cc_34 VNB N_C_c_426_n 0.0149127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_C_c_427_n 0.00184387f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.63
cc_36 VNB N_C_c_428_n 0.00134539f $X=-0.19 $Y=-0.245 $X2=2.88 $Y2=1.63
cc_37 VNB N_C_c_429_n 0.0231761f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.417
cc_38 VNB N_C_c_430_n 0.00463151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_219_392#_c_556_n 0.0177707f $X=-0.19 $Y=-0.245 $X2=3.38 $Y2=1.885
cc_40 VNB N_A_219_392#_c_557_n 0.0161712f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=1.54
cc_41 VNB N_A_219_392#_c_558_n 0.0157856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_219_392#_c_559_n 0.0181907f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.63
cc_43 VNB N_A_219_392#_c_560_n 0.00165849f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.63
cc_44 VNB N_A_219_392#_c_561_n 0.00444125f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.54
cc_45 VNB N_A_219_392#_c_562_n 0.00389952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_219_392#_c_563_n 0.00572055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_219_392#_c_564_n 0.00147192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_219_392#_c_565_n 9.85159e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_219_392#_c_566_n 0.0789898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VPWR_c_776_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_X_c_966_n 0.00302927f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=1.375
cc_52 VNB N_X_c_967_n 0.00762797f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.945
cc_53 VNB N_X_c_968_n 0.0109113f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=1.21
cc_54 VNB X 0.0142018f $X=-0.19 $Y=-0.245 $X2=2.88 $Y2=1.63
cc_55 VNB N_VGND_c_1025_n 0.0110036f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=1.375
cc_56 VNB N_VGND_c_1026_n 0.0505933f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.945
cc_57 VNB N_VGND_c_1027_n 0.0120081f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=1.3
cc_58 VNB N_VGND_c_1028_n 0.00447121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1029_n 0.0122631f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=1.21
cc_60 VNB N_VGND_c_1030_n 0.00730842f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.63
cc_61 VNB N_VGND_c_1031_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.63
cc_62 VNB N_VGND_c_1032_n 0.0305743f $X=-0.19 $Y=-0.245 $X2=2.88 $Y2=1.63
cc_63 VNB N_VGND_c_1033_n 0.0406425f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=1.54
cc_64 VNB N_VGND_c_1034_n 0.0404117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1035_n 0.0393298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1036_n 0.0191053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1037_n 0.016802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1038_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1039_n 0.00510664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1040_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1041_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1042_n 0.423803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_114_125#_c_1119_n 0.0169875f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.885
cc_74 VNB N_A_114_125#_c_1120_n 0.0041948f $X=-0.19 $Y=-0.245 $X2=1.515
+ $Y2=0.945
cc_75 VNB N_A_114_125#_c_1121_n 0.0103612f $X=-0.19 $Y=-0.245 $X2=2.88 $Y2=1.885
cc_76 VNB N_A_504_125#_c_1145_n 8.44865e-19 $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.46
cc_77 VNB N_A_504_125#_c_1146_n 0.012904f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.945
cc_78 VNB N_A_504_125#_c_1147_n 0.00227888f $X=-0.19 $Y=-0.245 $X2=1.515
+ $Y2=0.945
cc_79 VNB N_A_504_125#_c_1148_n 0.00659005f $X=-0.19 $Y=-0.245 $X2=2.88
+ $Y2=1.885
cc_80 VNB N_A_906_78#_c_1179_n 0.0131581f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.885
cc_81 VNB N_A_906_78#_c_1180_n 5.5847e-19 $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.945
cc_82 VNB N_A_906_78#_c_1181_n 0.00287386f $X=-0.19 $Y=-0.245 $X2=2.88 $Y2=1.885
cc_83 VPB N_B_c_152_n 0.0145087f $X=-0.19 $Y=1.66 $X2=1.02 $Y2=1.885
cc_84 VPB N_B_c_153_n 0.0145865f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=1.885
cc_85 VPB N_B_c_154_n 0.0145103f $X=-0.19 $Y=1.66 $X2=2.88 $Y2=1.885
cc_86 VPB N_B_c_155_n 0.0148849f $X=-0.19 $Y=1.66 $X2=3.38 $Y2=1.885
cc_87 VPB N_B_c_156_n 0.00228472f $X=-0.19 $Y=1.66 $X2=1.3 $Y2=1.54
cc_88 VPB B 0.00289288f $X=-0.19 $Y=1.66 $X2=3.035 $Y2=1.21
cc_89 VPB N_B_c_149_n 0.0345401f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=1.63
cc_90 VPB N_B_c_150_n 0.0351375f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=1.63
cc_91 VPB N_A_c_259_n 0.011772f $X=-0.19 $Y=1.66 $X2=1.085 $Y2=0.945
cc_92 VPB N_A_c_275_n 0.0269648f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=1.885
cc_93 VPB N_A_c_262_n 0.0340824f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=0.945
cc_94 VPB N_A_c_264_n 0.0353331f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=1.375
cc_95 VPB N_A_c_268_n 0.0076343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_c_279_n 0.0231953f $X=-0.19 $Y=1.66 $X2=2.525 $Y2=1.215
cc_97 VPB N_A_c_280_n 0.0133023f $X=-0.19 $Y=1.66 $X2=2.88 $Y2=1.63
cc_98 VPB N_A_c_272_n 0.00164609f $X=-0.19 $Y=1.66 $X2=2.955 $Y2=1.54
cc_99 VPB A 0.006713f $X=-0.19 $Y=1.66 $X2=2.64 $Y2=1.417
cc_100 VPB N_C_c_418_n 0.00725229f $X=-0.19 $Y=1.66 $X2=1.02 $Y2=2.46
cc_101 VPB N_C_c_432_n 0.0212057f $X=-0.19 $Y=1.66 $X2=1.02 $Y2=2.46
cc_102 VPB N_C_c_422_n 0.0352552f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=0.945
cc_103 VPB N_C_c_434_n 0.0159383f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=1.375
cc_104 VPB N_C_c_435_n 0.0155164f $X=-0.19 $Y=1.66 $X2=1.3 $Y2=1.54
cc_105 VPB N_C_c_428_n 0.00161416f $X=-0.19 $Y=1.66 $X2=2.88 $Y2=1.63
cc_106 VPB N_C_c_429_n 0.0300497f $X=-0.19 $Y=1.66 $X2=3.12 $Y2=1.417
cc_107 VPB N_C_c_430_n 0.00352284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_219_392#_c_567_n 0.0162875f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=1.375
cc_109 VPB N_A_219_392#_c_568_n 0.0156175f $X=-0.19 $Y=1.66 $X2=1.3 $Y2=1.3
cc_110 VPB N_A_219_392#_c_569_n 0.015079f $X=-0.19 $Y=1.66 $X2=1.465 $Y2=1.215
cc_111 VPB N_A_219_392#_c_570_n 0.0186861f $X=-0.19 $Y=1.66 $X2=1.085 $Y2=1.63
cc_112 VPB N_A_219_392#_c_561_n 0.00246775f $X=-0.19 $Y=1.66 $X2=2.955 $Y2=1.54
cc_113 VPB N_A_219_392#_c_572_n 0.00299985f $X=-0.19 $Y=1.66 $X2=2.955 $Y2=1.54
cc_114 VPB N_A_219_392#_c_573_n 0.00266479f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_219_392#_c_563_n 0.00963371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_219_392#_c_566_n 0.054805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_777_n 0.0111306f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=1.375
cc_118 VPB N_VPWR_c_778_n 0.054022f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=0.945
cc_119 VPB N_VPWR_c_779_n 0.00825864f $X=-0.19 $Y=1.66 $X2=1.3 $Y2=1.54
cc_120 VPB N_VPWR_c_780_n 0.00934999f $X=-0.19 $Y=1.66 $X2=1.465 $Y2=1.215
cc_121 VPB N_VPWR_c_781_n 0.00933855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_782_n 0.0198086f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=1.63
cc_123 VPB N_VPWR_c_783_n 0.00504372f $X=-0.19 $Y=1.66 $X2=2.955 $Y2=1.63
cc_124 VPB N_VPWR_c_784_n 0.0120106f $X=-0.19 $Y=1.66 $X2=2.955 $Y2=1.54
cc_125 VPB N_VPWR_c_785_n 0.0559634f $X=-0.19 $Y=1.66 $X2=3.38 $Y2=1.63
cc_126 VPB N_VPWR_c_786_n 0.0408388f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_787_n 0.0400334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_788_n 0.0436498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_789_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_790_n 0.00497144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_791_n 0.00631788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_792_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_793_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_776_n 0.093429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_119_392#_c_888_n 0.00455202f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=0.945
cc_136 VPB N_A_119_392#_c_889_n 0.0022931f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=0.945
cc_137 VPB N_A_501_392#_c_914_n 0.00498811f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=0.945
cc_138 VPB N_A_501_392#_c_915_n 0.00217391f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=0.945
cc_139 VPB N_A_905_392#_c_941_n 0.00255137f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.46
cc_140 VPB N_A_905_392#_c_942_n 0.00255137f $X=-0.19 $Y=1.66 $X2=2.88 $Y2=2.46
cc_141 VPB N_X_c_970_n 0.00257348f $X=-0.19 $Y=1.66 $X2=2.88 $Y2=2.46
cc_142 VPB N_X_c_971_n 0.00293853f $X=-0.19 $Y=1.66 $X2=1.3 $Y2=1.54
cc_143 VPB N_X_c_972_n 0.00180921f $X=-0.19 $Y=1.66 $X2=1.465 $Y2=1.215
cc_144 N_B_c_144_n N_A_M1013_g 0.0168277f $X=1.085 $Y=1.375 $X2=0 $Y2=0
cc_145 N_B_c_149_n N_A_c_259_n 0.00619213f $X=1.47 $Y=1.63 $X2=0 $Y2=0
cc_146 N_B_c_152_n N_A_c_275_n 0.024506f $X=1.02 $Y=1.885 $X2=0 $Y2=0
cc_147 N_B_c_144_n N_A_c_260_n 0.00737233f $X=1.085 $Y=1.375 $X2=0 $Y2=0
cc_148 N_B_c_145_n N_A_c_260_n 0.00737233f $X=1.515 $Y=1.375 $X2=0 $Y2=0
cc_149 N_B_c_153_n N_A_c_262_n 0.0337462f $X=1.47 $Y=1.885 $X2=0 $Y2=0
cc_150 N_B_c_156_n N_A_c_262_n 2.4772e-19 $X=1.3 $Y=1.54 $X2=0 $Y2=0
cc_151 N_B_c_149_n N_A_c_262_n 0.024583f $X=1.47 $Y=1.63 $X2=0 $Y2=0
cc_152 N_B_c_151_n N_A_c_262_n 0.00125954f $X=2.525 $Y=1.417 $X2=0 $Y2=0
cc_153 N_B_c_145_n N_A_M1019_g 0.0270984f $X=1.515 $Y=1.375 $X2=0 $Y2=0
cc_154 N_B_c_156_n N_A_M1019_g 7.96256e-19 $X=1.3 $Y=1.54 $X2=0 $Y2=0
cc_155 N_B_c_151_n N_A_M1019_g 0.0146196f $X=2.525 $Y=1.417 $X2=0 $Y2=0
cc_156 N_B_c_144_n N_A_c_270_n 7.38627e-19 $X=1.085 $Y=1.375 $X2=0 $Y2=0
cc_157 N_B_c_149_n N_A_c_270_n 0.0100847f $X=1.47 $Y=1.63 $X2=0 $Y2=0
cc_158 N_B_c_154_n N_A_c_280_n 0.00849388f $X=2.88 $Y=1.885 $X2=0 $Y2=0
cc_159 N_B_c_155_n N_A_c_280_n 0.00874123f $X=3.38 $Y=1.885 $X2=0 $Y2=0
cc_160 B N_A_c_280_n 0.0562262f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_161 N_B_c_150_n N_A_c_280_n 0.0210062f $X=3.365 $Y=1.63 $X2=0 $Y2=0
cc_162 N_B_c_151_n N_A_c_280_n 0.00680468f $X=2.525 $Y=1.417 $X2=0 $Y2=0
cc_163 N_B_c_156_n A 0.0105625f $X=1.3 $Y=1.54 $X2=0 $Y2=0
cc_164 B A 0.0162995f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_165 N_B_c_149_n A 0.00162582f $X=1.47 $Y=1.63 $X2=0 $Y2=0
cc_166 N_B_c_151_n A 0.0365244f $X=2.525 $Y=1.417 $X2=0 $Y2=0
cc_167 N_B_c_150_n N_C_c_417_n 0.0230256f $X=3.365 $Y=1.63 $X2=-0.19 $Y2=-0.245
cc_168 N_B_c_151_n N_C_c_417_n 0.0010529f $X=2.525 $Y=1.417 $X2=-0.19 $Y2=-0.245
cc_169 N_B_c_154_n N_C_c_432_n 0.0349777f $X=2.88 $Y=1.885 $X2=0 $Y2=0
cc_170 N_B_c_146_n N_C_M1007_g 0.0197883f $X=2.935 $Y=1.375 $X2=0 $Y2=0
cc_171 B N_C_M1007_g 0.00829523f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_172 N_B_c_151_n N_C_M1007_g 0.0165505f $X=2.525 $Y=1.417 $X2=0 $Y2=0
cc_173 N_B_c_146_n N_C_c_420_n 0.00738071f $X=2.935 $Y=1.375 $X2=0 $Y2=0
cc_174 N_B_c_147_n N_C_c_420_n 0.00737233f $X=3.365 $Y=1.375 $X2=0 $Y2=0
cc_175 N_B_c_155_n N_C_c_422_n 0.0343197f $X=3.38 $Y=1.885 $X2=0 $Y2=0
cc_176 B N_C_c_422_n 2.24587e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_177 N_B_c_150_n N_C_c_422_n 0.0281482f $X=3.365 $Y=1.63 $X2=0 $Y2=0
cc_178 N_B_c_147_n N_C_M1017_g 0.020099f $X=3.365 $Y=1.375 $X2=0 $Y2=0
cc_179 N_B_c_147_n N_C_c_430_n 0.00483014f $X=3.365 $Y=1.375 $X2=0 $Y2=0
cc_180 B N_C_c_430_n 0.029095f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_181 N_B_c_150_n N_C_c_430_n 0.0019154f $X=3.365 $Y=1.63 $X2=0 $Y2=0
cc_182 N_B_c_198_p N_A_219_392#_M1016_s 0.00182762f $X=1.465 $Y=1.215 $X2=-0.19
+ $Y2=-0.245
cc_183 B N_A_219_392#_M1024_s 0.00196283f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_184 N_B_c_144_n N_A_219_392#_c_560_n 0.0163458f $X=1.085 $Y=1.375 $X2=0 $Y2=0
cc_185 N_B_c_145_n N_A_219_392#_c_560_n 0.00434482f $X=1.515 $Y=1.375 $X2=0
+ $Y2=0
cc_186 N_B_c_198_p N_A_219_392#_c_560_n 0.0180006f $X=1.465 $Y=1.215 $X2=0 $Y2=0
cc_187 N_B_c_149_n N_A_219_392#_c_560_n 4.29435e-19 $X=1.47 $Y=1.63 $X2=0 $Y2=0
cc_188 N_B_c_144_n N_A_219_392#_c_561_n 0.00290479f $X=1.085 $Y=1.375 $X2=0
+ $Y2=0
cc_189 N_B_c_156_n N_A_219_392#_c_561_n 0.029127f $X=1.3 $Y=1.54 $X2=0 $Y2=0
cc_190 N_B_c_198_p N_A_219_392#_c_561_n 0.00844566f $X=1.465 $Y=1.215 $X2=0
+ $Y2=0
cc_191 N_B_c_149_n N_A_219_392#_c_561_n 0.0138261f $X=1.47 $Y=1.63 $X2=0 $Y2=0
cc_192 N_B_c_152_n N_A_219_392#_c_572_n 0.0112277f $X=1.02 $Y=1.885 $X2=0 $Y2=0
cc_193 N_B_c_153_n N_A_219_392#_c_572_n 0.00405016f $X=1.47 $Y=1.885 $X2=0 $Y2=0
cc_194 N_B_c_156_n N_A_219_392#_c_572_n 0.0214939f $X=1.3 $Y=1.54 $X2=0 $Y2=0
cc_195 N_B_c_149_n N_A_219_392#_c_572_n 0.0110212f $X=1.47 $Y=1.63 $X2=0 $Y2=0
cc_196 N_B_c_153_n N_A_219_392#_c_590_n 0.00303687f $X=1.47 $Y=1.885 $X2=0 $Y2=0
cc_197 N_B_c_153_n N_A_219_392#_c_591_n 0.0123045f $X=1.47 $Y=1.885 $X2=0 $Y2=0
cc_198 N_B_c_154_n N_A_219_392#_c_591_n 0.0125075f $X=2.88 $Y=1.885 $X2=0 $Y2=0
cc_199 N_B_c_156_n N_A_219_392#_c_591_n 0.00163528f $X=1.3 $Y=1.54 $X2=0 $Y2=0
cc_200 N_B_c_155_n N_A_219_392#_c_594_n 0.00503628f $X=3.38 $Y=1.885 $X2=0 $Y2=0
cc_201 N_B_c_147_n N_A_219_392#_c_595_n 0.0127517f $X=3.365 $Y=1.375 $X2=0 $Y2=0
cc_202 N_B_c_155_n N_A_219_392#_c_596_n 0.00968286f $X=3.38 $Y=1.885 $X2=0 $Y2=0
cc_203 N_B_c_153_n N_A_219_392#_c_597_n 8.12288e-19 $X=1.47 $Y=1.885 $X2=0 $Y2=0
cc_204 N_B_c_155_n N_A_219_392#_c_598_n 4.10389e-19 $X=3.38 $Y=1.885 $X2=0 $Y2=0
cc_205 N_B_c_147_n N_A_219_392#_c_564_n 0.00593229f $X=3.365 $Y=1.375 $X2=0
+ $Y2=0
cc_206 B N_A_219_392#_c_564_n 0.0140293f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_207 N_B_c_150_n N_A_219_392#_c_564_n 4.3034e-19 $X=3.365 $Y=1.63 $X2=0 $Y2=0
cc_208 N_B_c_152_n N_VPWR_c_786_n 0.00278271f $X=1.02 $Y=1.885 $X2=0 $Y2=0
cc_209 N_B_c_153_n N_VPWR_c_786_n 0.00278257f $X=1.47 $Y=1.885 $X2=0 $Y2=0
cc_210 N_B_c_154_n N_VPWR_c_787_n 0.00278257f $X=2.88 $Y=1.885 $X2=0 $Y2=0
cc_211 N_B_c_155_n N_VPWR_c_787_n 0.00278271f $X=3.38 $Y=1.885 $X2=0 $Y2=0
cc_212 N_B_c_152_n N_VPWR_c_776_n 0.00354337f $X=1.02 $Y=1.885 $X2=0 $Y2=0
cc_213 N_B_c_153_n N_VPWR_c_776_n 0.00353905f $X=1.47 $Y=1.885 $X2=0 $Y2=0
cc_214 N_B_c_154_n N_VPWR_c_776_n 0.00354366f $X=2.88 $Y=1.885 $X2=0 $Y2=0
cc_215 N_B_c_155_n N_VPWR_c_776_n 0.00354798f $X=3.38 $Y=1.885 $X2=0 $Y2=0
cc_216 N_B_c_152_n N_A_119_392#_c_888_n 0.0142212f $X=1.02 $Y=1.885 $X2=0 $Y2=0
cc_217 N_B_c_153_n N_A_119_392#_c_888_n 0.0100163f $X=1.47 $Y=1.885 $X2=0 $Y2=0
cc_218 N_B_c_152_n N_A_119_392#_c_892_n 4.94775e-19 $X=1.02 $Y=1.885 $X2=0 $Y2=0
cc_219 N_B_c_153_n N_A_119_392#_c_892_n 0.00522005f $X=1.47 $Y=1.885 $X2=0 $Y2=0
cc_220 N_B_c_154_n N_A_501_392#_c_916_n 0.00516295f $X=2.88 $Y=1.885 $X2=0 $Y2=0
cc_221 N_B_c_155_n N_A_501_392#_c_916_n 2.69714e-19 $X=3.38 $Y=1.885 $X2=0 $Y2=0
cc_222 N_B_c_154_n N_A_501_392#_c_914_n 0.00857759f $X=2.88 $Y=1.885 $X2=0 $Y2=0
cc_223 N_B_c_155_n N_A_501_392#_c_914_n 0.011466f $X=3.38 $Y=1.885 $X2=0 $Y2=0
cc_224 N_B_c_154_n N_A_501_392#_c_915_n 0.00228491f $X=2.88 $Y=1.885 $X2=0 $Y2=0
cc_225 N_B_c_151_n N_VGND_M1019_d 0.00176461f $X=2.525 $Y=1.417 $X2=0 $Y2=0
cc_226 N_B_c_144_n N_VGND_c_1026_n 9.33445e-19 $X=1.085 $Y=1.375 $X2=0 $Y2=0
cc_227 N_B_c_151_n N_VGND_c_1027_n 0.0135055f $X=2.525 $Y=1.417 $X2=0 $Y2=0
cc_228 N_B_c_151_n N_A_114_125#_M1023_d 0.00250873f $X=2.525 $Y=1.417 $X2=0
+ $Y2=0
cc_229 N_B_c_144_n N_A_114_125#_c_1119_n 0.00150539f $X=1.085 $Y=1.375 $X2=0
+ $Y2=0
cc_230 N_B_c_145_n N_A_114_125#_c_1119_n 0.00329102f $X=1.515 $Y=1.375 $X2=0
+ $Y2=0
cc_231 N_B_c_145_n N_A_114_125#_c_1120_n 0.00503319f $X=1.515 $Y=1.375 $X2=0
+ $Y2=0
cc_232 N_B_c_151_n N_A_114_125#_c_1120_n 0.0210243f $X=2.525 $Y=1.417 $X2=0
+ $Y2=0
cc_233 N_B_c_144_n N_A_114_125#_c_1121_n 0.00334268f $X=1.085 $Y=1.375 $X2=0
+ $Y2=0
cc_234 B N_A_504_125#_M1007_s 0.0026453f $X=3.035 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_235 N_B_c_146_n N_A_504_125#_c_1145_n 0.00779152f $X=2.935 $Y=1.375 $X2=0
+ $Y2=0
cc_236 N_B_c_147_n N_A_504_125#_c_1145_n 4.41164e-19 $X=3.365 $Y=1.375 $X2=0
+ $Y2=0
cc_237 N_B_c_150_n N_A_504_125#_c_1145_n 2.01734e-19 $X=3.365 $Y=1.63 $X2=0
+ $Y2=0
cc_238 N_B_c_151_n N_A_504_125#_c_1145_n 0.0214083f $X=2.525 $Y=1.417 $X2=0
+ $Y2=0
cc_239 N_B_c_146_n N_A_504_125#_c_1146_n 0.00307326f $X=2.935 $Y=1.375 $X2=0
+ $Y2=0
cc_240 N_B_c_147_n N_A_504_125#_c_1146_n 0.00152378f $X=3.365 $Y=1.375 $X2=0
+ $Y2=0
cc_241 N_B_c_147_n N_A_504_125#_c_1148_n 0.00187846f $X=3.365 $Y=1.375 $X2=0
+ $Y2=0
cc_242 N_A_M1019_g N_C_c_417_n 0.00678625f $X=2.015 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_243 N_A_c_262_n N_C_c_418_n 0.0195097f $X=1.92 $Y=1.885 $X2=0 $Y2=0
cc_244 A N_C_c_418_n 0.0064364f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_245 N_A_c_262_n N_C_c_432_n 0.0342399f $X=1.92 $Y=1.885 $X2=0 $Y2=0
cc_246 N_A_c_280_n N_C_c_432_n 0.0136312f $X=4.24 $Y=1.96 $X2=0 $Y2=0
cc_247 N_A_M1019_g N_C_M1007_g 0.0190413f $X=2.015 $Y=0.945 $X2=0 $Y2=0
cc_248 N_A_c_267_n N_C_c_420_n 0.021187f $X=4.53 $Y=0.18 $X2=0 $Y2=0
cc_249 N_A_c_260_n N_C_c_421_n 0.0190413f $X=1.94 $Y=0.18 $X2=0 $Y2=0
cc_250 N_A_c_264_n N_C_c_422_n 0.0521082f $X=4.45 $Y=1.885 $X2=0 $Y2=0
cc_251 N_A_c_280_n N_C_c_422_n 0.0140686f $X=4.24 $Y=1.96 $X2=0 $Y2=0
cc_252 N_A_c_272_n N_C_c_422_n 0.00308354f $X=4.405 $Y=1.635 $X2=0 $Y2=0
cc_253 N_A_M1004_g N_C_M1017_g 0.021187f $X=4.455 $Y=0.71 $X2=0 $Y2=0
cc_254 N_A_c_264_n N_C_c_434_n 0.0343789f $X=4.45 $Y=1.885 $X2=0 $Y2=0
cc_255 N_A_c_280_n N_C_c_434_n 0.00211521f $X=4.24 $Y=1.96 $X2=0 $Y2=0
cc_256 N_A_M1004_g N_C_M1002_g 0.0282378f $X=4.455 $Y=0.71 $X2=0 $Y2=0
cc_257 N_A_c_266_n N_C_M1002_g 0.00882199f $X=5.75 $Y=0.18 $X2=0 $Y2=0
cc_258 N_A_c_279_n N_C_c_435_n 0.032254f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_259 N_A_c_266_n N_C_M1008_g 0.00897756f $X=5.75 $Y=0.18 $X2=0 $Y2=0
cc_260 N_A_M1009_g N_C_M1008_g 0.0192578f $X=5.825 $Y=0.915 $X2=0 $Y2=0
cc_261 N_A_c_271_n N_C_M1008_g 0.0083954f $X=5.805 $Y=1.46 $X2=0 $Y2=0
cc_262 N_A_c_264_n N_C_c_426_n 0.00125364f $X=4.45 $Y=1.885 $X2=0 $Y2=0
cc_263 N_A_M1004_g N_C_c_426_n 0.0112003f $X=4.455 $Y=0.71 $X2=0 $Y2=0
cc_264 N_A_c_280_n N_C_c_426_n 0.007338f $X=4.24 $Y=1.96 $X2=0 $Y2=0
cc_265 N_A_c_272_n N_C_c_426_n 0.0253031f $X=4.405 $Y=1.635 $X2=0 $Y2=0
cc_266 N_A_M1004_g N_C_c_427_n 0.00339628f $X=4.455 $Y=0.71 $X2=0 $Y2=0
cc_267 N_A_c_264_n N_C_c_428_n 0.00205988f $X=4.45 $Y=1.885 $X2=0 $Y2=0
cc_268 N_A_c_272_n N_C_c_428_n 0.0251563f $X=4.405 $Y=1.635 $X2=0 $Y2=0
cc_269 N_A_c_264_n N_C_c_429_n 0.0212475f $X=4.45 $Y=1.885 $X2=0 $Y2=0
cc_270 N_A_c_268_n N_C_c_429_n 0.0200681f $X=5.8 $Y=1.795 $X2=0 $Y2=0
cc_271 N_A_c_280_n N_C_c_429_n 2.53908e-19 $X=4.24 $Y=1.96 $X2=0 $Y2=0
cc_272 N_A_c_272_n N_C_c_429_n 0.0019786f $X=4.405 $Y=1.635 $X2=0 $Y2=0
cc_273 N_A_c_264_n N_C_c_430_n 7.92676e-19 $X=4.45 $Y=1.885 $X2=0 $Y2=0
cc_274 N_A_M1004_g N_C_c_430_n 0.00107017f $X=4.455 $Y=0.71 $X2=0 $Y2=0
cc_275 N_A_c_280_n N_C_c_430_n 0.0414297f $X=4.24 $Y=1.96 $X2=0 $Y2=0
cc_276 N_A_c_272_n N_C_c_430_n 0.01436f $X=4.405 $Y=1.635 $X2=0 $Y2=0
cc_277 N_A_c_280_n N_A_219_392#_M1001_d 0.00250873f $X=4.24 $Y=1.96 $X2=0 $Y2=0
cc_278 N_A_c_268_n N_A_219_392#_c_567_n 0.00449613f $X=5.8 $Y=1.795 $X2=0 $Y2=0
cc_279 N_A_c_279_n N_A_219_392#_c_567_n 0.0178001f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_280 N_A_M1009_g N_A_219_392#_c_556_n 0.0170887f $X=5.825 $Y=0.915 $X2=0 $Y2=0
cc_281 N_A_M1013_g N_A_219_392#_c_560_n 0.00241064f $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_282 N_A_c_260_n N_A_219_392#_c_560_n 2.56684e-19 $X=1.94 $Y=0.18 $X2=0 $Y2=0
cc_283 N_A_M1013_g N_A_219_392#_c_561_n 0.00381203f $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_284 N_A_c_270_n N_A_219_392#_c_561_n 0.0112956f $X=0.515 $Y=1.49 $X2=0 $Y2=0
cc_285 N_A_c_275_n N_A_219_392#_c_572_n 0.00273184f $X=0.52 $Y=1.885 $X2=0 $Y2=0
cc_286 N_A_c_262_n N_A_219_392#_c_572_n 7.87646e-19 $X=1.92 $Y=1.885 $X2=0 $Y2=0
cc_287 N_A_c_262_n N_A_219_392#_c_590_n 8.04986e-19 $X=1.92 $Y=1.885 $X2=0 $Y2=0
cc_288 N_A_c_262_n N_A_219_392#_c_591_n 0.0169039f $X=1.92 $Y=1.885 $X2=0 $Y2=0
cc_289 N_A_c_280_n N_A_219_392#_c_591_n 0.0354782f $X=4.24 $Y=1.96 $X2=0 $Y2=0
cc_290 A N_A_219_392#_c_591_n 0.0227073f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_291 N_A_M1004_g N_A_219_392#_c_595_n 0.0123829f $X=4.455 $Y=0.71 $X2=0 $Y2=0
cc_292 N_A_c_266_n N_A_219_392#_c_595_n 7.06373e-19 $X=5.75 $Y=0.18 $X2=0 $Y2=0
cc_293 N_A_c_264_n N_A_219_392#_c_596_n 0.0157796f $X=4.45 $Y=1.885 $X2=0 $Y2=0
cc_294 N_A_c_280_n N_A_219_392#_c_596_n 0.0704772f $X=4.24 $Y=1.96 $X2=0 $Y2=0
cc_295 N_A_M1009_g N_A_219_392#_c_562_n 0.0036791f $X=5.825 $Y=0.915 $X2=0 $Y2=0
cc_296 N_A_c_271_n N_A_219_392#_c_562_n 7.34435e-19 $X=5.805 $Y=1.46 $X2=0 $Y2=0
cc_297 N_A_c_268_n N_A_219_392#_c_573_n 0.00443587f $X=5.8 $Y=1.795 $X2=0 $Y2=0
cc_298 N_A_c_279_n N_A_219_392#_c_573_n 0.00139183f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_299 N_A_c_268_n N_A_219_392#_c_563_n 0.0165223f $X=5.8 $Y=1.795 $X2=0 $Y2=0
cc_300 N_A_c_271_n N_A_219_392#_c_563_n 0.0115597f $X=5.805 $Y=1.46 $X2=0 $Y2=0
cc_301 N_A_c_280_n N_A_219_392#_c_598_n 0.0198661f $X=4.24 $Y=1.96 $X2=0 $Y2=0
cc_302 N_A_c_264_n N_A_219_392#_c_627_n 8.79478e-19 $X=4.45 $Y=1.885 $X2=0 $Y2=0
cc_303 N_A_c_279_n N_A_219_392#_c_627_n 0.00238646f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_304 N_A_c_268_n N_A_219_392#_c_566_n 0.0150136f $X=5.8 $Y=1.795 $X2=0 $Y2=0
cc_305 N_A_c_271_n N_A_219_392#_c_566_n 0.00634523f $X=5.805 $Y=1.46 $X2=0 $Y2=0
cc_306 N_A_c_280_n N_VPWR_M1029_s 2.34434e-19 $X=4.24 $Y=1.96 $X2=0 $Y2=0
cc_307 A N_VPWR_M1029_s 0.00317248f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_308 N_A_c_280_n N_VPWR_M1027_d 0.00337505f $X=4.24 $Y=1.96 $X2=0 $Y2=0
cc_309 N_A_c_275_n N_VPWR_c_778_n 0.0103974f $X=0.52 $Y=1.885 $X2=0 $Y2=0
cc_310 N_A_c_262_n N_VPWR_c_779_n 0.00300056f $X=1.92 $Y=1.885 $X2=0 $Y2=0
cc_311 N_A_c_264_n N_VPWR_c_780_n 0.00574337f $X=4.45 $Y=1.885 $X2=0 $Y2=0
cc_312 N_A_c_279_n N_VPWR_c_781_n 0.0116208f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_313 N_A_c_275_n N_VPWR_c_786_n 0.0044313f $X=0.52 $Y=1.885 $X2=0 $Y2=0
cc_314 N_A_c_262_n N_VPWR_c_786_n 0.0044313f $X=1.92 $Y=1.885 $X2=0 $Y2=0
cc_315 N_A_c_264_n N_VPWR_c_788_n 0.00445602f $X=4.45 $Y=1.885 $X2=0 $Y2=0
cc_316 N_A_c_279_n N_VPWR_c_788_n 0.00445602f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_317 N_A_c_275_n N_VPWR_c_776_n 0.00857418f $X=0.52 $Y=1.885 $X2=0 $Y2=0
cc_318 N_A_c_262_n N_VPWR_c_776_n 0.0085404f $X=1.92 $Y=1.885 $X2=0 $Y2=0
cc_319 N_A_c_264_n N_VPWR_c_776_n 0.00858504f $X=4.45 $Y=1.885 $X2=0 $Y2=0
cc_320 N_A_c_279_n N_VPWR_c_776_n 0.00858228f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_321 N_A_c_275_n N_A_119_392#_c_894_n 0.00862798f $X=0.52 $Y=1.885 $X2=0 $Y2=0
cc_322 N_A_c_262_n N_A_119_392#_c_888_n 0.00323938f $X=1.92 $Y=1.885 $X2=0 $Y2=0
cc_323 N_A_c_275_n N_A_119_392#_c_889_n 0.00350568f $X=0.52 $Y=1.885 $X2=0 $Y2=0
cc_324 N_A_c_262_n N_A_119_392#_c_892_n 0.00396652f $X=1.92 $Y=1.885 $X2=0 $Y2=0
cc_325 N_A_c_280_n N_A_501_392#_M1012_s 0.00198204f $X=4.24 $Y=1.96 $X2=-0.19
+ $Y2=-0.245
cc_326 N_A_c_280_n N_A_501_392#_M1005_s 0.00251484f $X=4.24 $Y=1.96 $X2=0 $Y2=0
cc_327 N_A_c_264_n N_A_905_392#_c_941_n 0.00542733f $X=4.45 $Y=1.885 $X2=0 $Y2=0
cc_328 N_A_c_279_n N_A_905_392#_c_942_n 0.00594165f $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_329 N_A_c_279_n N_X_c_973_n 4.56552e-19 $X=5.8 $Y=1.885 $X2=0 $Y2=0
cc_330 N_A_M1013_g N_VGND_c_1026_n 0.0239301f $X=0.495 $Y=0.945 $X2=0 $Y2=0
cc_331 N_A_c_261_n N_VGND_c_1026_n 0.00763335f $X=0.57 $Y=0.18 $X2=0 $Y2=0
cc_332 N_A_c_260_n N_VGND_c_1027_n 0.00600873f $X=1.94 $Y=0.18 $X2=0 $Y2=0
cc_333 N_A_c_267_n N_VGND_c_1028_n 0.00599801f $X=4.53 $Y=0.18 $X2=0 $Y2=0
cc_334 N_A_c_266_n N_VGND_c_1029_n 0.0131476f $X=5.75 $Y=0.18 $X2=0 $Y2=0
cc_335 N_A_c_261_n N_VGND_c_1033_n 0.0395853f $X=0.57 $Y=0.18 $X2=0 $Y2=0
cc_336 N_A_c_267_n N_VGND_c_1035_n 0.0361594f $X=4.53 $Y=0.18 $X2=0 $Y2=0
cc_337 N_A_c_260_n N_VGND_c_1042_n 0.0432928f $X=1.94 $Y=0.18 $X2=0 $Y2=0
cc_338 N_A_c_261_n N_VGND_c_1042_n 0.00749832f $X=0.57 $Y=0.18 $X2=0 $Y2=0
cc_339 N_A_c_266_n N_VGND_c_1042_n 0.0391765f $X=5.75 $Y=0.18 $X2=0 $Y2=0
cc_340 N_A_c_267_n N_VGND_c_1042_n 0.00546436f $X=4.53 $Y=0.18 $X2=0 $Y2=0
cc_341 N_A_c_260_n N_A_114_125#_c_1119_n 0.0163379f $X=1.94 $Y=0.18 $X2=0 $Y2=0
cc_342 N_A_M1019_g N_A_114_125#_c_1119_n 0.00609242f $X=2.015 $Y=0.945 $X2=0
+ $Y2=0
cc_343 N_A_M1019_g N_A_114_125#_c_1120_n 0.00850643f $X=2.015 $Y=0.945 $X2=0
+ $Y2=0
cc_344 N_A_M1013_g N_A_114_125#_c_1121_n 0.0063893f $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_345 N_A_c_260_n N_A_114_125#_c_1121_n 0.007046f $X=1.94 $Y=0.18 $X2=0 $Y2=0
cc_346 N_A_M1004_g N_A_906_78#_c_1179_n 4.61883e-19 $X=4.455 $Y=0.71 $X2=0 $Y2=0
cc_347 N_A_c_266_n N_A_906_78#_c_1179_n 0.01728f $X=5.75 $Y=0.18 $X2=0 $Y2=0
cc_348 N_A_M1009_g N_A_906_78#_c_1179_n 0.00591191f $X=5.825 $Y=0.915 $X2=0
+ $Y2=0
cc_349 N_A_M1009_g N_A_906_78#_c_1180_n 0.00848181f $X=5.825 $Y=0.915 $X2=0
+ $Y2=0
cc_350 N_A_M1004_g N_A_906_78#_c_1181_n 0.00674166f $X=4.455 $Y=0.71 $X2=0 $Y2=0
cc_351 N_A_c_266_n N_A_906_78#_c_1181_n 0.00710114f $X=5.75 $Y=0.18 $X2=0 $Y2=0
cc_352 N_A_c_267_n N_A_906_78#_c_1181_n 2.05582e-19 $X=4.53 $Y=0.18 $X2=0 $Y2=0
cc_353 N_C_c_432_n N_A_219_392#_c_591_n 0.0150958f $X=2.43 $Y=1.885 $X2=0 $Y2=0
cc_354 N_C_c_422_n N_A_219_392#_c_594_n 7.18055e-19 $X=3.88 $Y=1.885 $X2=0 $Y2=0
cc_355 N_C_c_420_n N_A_219_392#_c_595_n 3.38974e-19 $X=3.88 $Y=0.18 $X2=0 $Y2=0
cc_356 N_C_c_422_n N_A_219_392#_c_595_n 7.25114e-19 $X=3.88 $Y=1.885 $X2=0 $Y2=0
cc_357 N_C_M1017_g N_A_219_392#_c_595_n 0.0126701f $X=3.955 $Y=0.71 $X2=0 $Y2=0
cc_358 N_C_M1002_g N_A_219_392#_c_595_n 0.0104894f $X=4.965 $Y=0.915 $X2=0 $Y2=0
cc_359 N_C_c_426_n N_A_219_392#_c_595_n 0.056185f $X=4.755 $Y=1.215 $X2=0 $Y2=0
cc_360 N_C_c_428_n N_A_219_392#_c_595_n 0.00421159f $X=5.055 $Y=1.635 $X2=0
+ $Y2=0
cc_361 N_C_c_429_n N_A_219_392#_c_595_n 2.02977e-19 $X=5.35 $Y=1.677 $X2=0 $Y2=0
cc_362 N_C_c_430_n N_A_219_392#_c_595_n 0.0386737f $X=3.747 $Y=1.215 $X2=0 $Y2=0
cc_363 N_C_c_422_n N_A_219_392#_c_596_n 0.0156265f $X=3.88 $Y=1.885 $X2=0 $Y2=0
cc_364 N_C_c_434_n N_A_219_392#_c_596_n 0.00900921f $X=4.9 $Y=1.885 $X2=0 $Y2=0
cc_365 N_C_c_428_n N_A_219_392#_c_596_n 0.00642995f $X=5.055 $Y=1.635 $X2=0
+ $Y2=0
cc_366 N_C_M1002_g N_A_219_392#_c_562_n 0.00103641f $X=4.965 $Y=0.915 $X2=0
+ $Y2=0
cc_367 N_C_M1008_g N_A_219_392#_c_562_n 0.016944f $X=5.395 $Y=0.915 $X2=0 $Y2=0
cc_368 N_C_c_426_n N_A_219_392#_c_562_n 0.0100252f $X=4.755 $Y=1.215 $X2=0 $Y2=0
cc_369 N_C_c_427_n N_A_219_392#_c_562_n 0.00549671f $X=4.84 $Y=1.47 $X2=0 $Y2=0
cc_370 N_C_c_428_n N_A_219_392#_c_562_n 0.0273574f $X=5.055 $Y=1.635 $X2=0 $Y2=0
cc_371 N_C_c_429_n N_A_219_392#_c_562_n 0.00961323f $X=5.35 $Y=1.677 $X2=0 $Y2=0
cc_372 N_C_c_434_n N_A_219_392#_c_573_n 4.14699e-19 $X=4.9 $Y=1.885 $X2=0 $Y2=0
cc_373 N_C_c_435_n N_A_219_392#_c_573_n 0.00213029f $X=5.35 $Y=1.885 $X2=0 $Y2=0
cc_374 N_C_c_428_n N_A_219_392#_c_573_n 0.00911816f $X=5.055 $Y=1.635 $X2=0
+ $Y2=0
cc_375 N_C_c_429_n N_A_219_392#_c_573_n 0.00595618f $X=5.35 $Y=1.677 $X2=0 $Y2=0
cc_376 N_C_M1017_g N_A_219_392#_c_564_n 8.55015e-19 $X=3.955 $Y=0.71 $X2=0 $Y2=0
cc_377 N_C_c_434_n N_A_219_392#_c_627_n 0.00549003f $X=4.9 $Y=1.885 $X2=0 $Y2=0
cc_378 N_C_c_435_n N_A_219_392#_c_627_n 0.0153752f $X=5.35 $Y=1.885 $X2=0 $Y2=0
cc_379 N_C_c_428_n N_A_219_392#_c_627_n 0.0181464f $X=5.055 $Y=1.635 $X2=0 $Y2=0
cc_380 N_C_c_429_n N_A_219_392#_c_627_n 0.00663744f $X=5.35 $Y=1.677 $X2=0 $Y2=0
cc_381 N_C_c_432_n N_VPWR_c_779_n 0.00358761f $X=2.43 $Y=1.885 $X2=0 $Y2=0
cc_382 N_C_c_422_n N_VPWR_c_780_n 0.00402278f $X=3.88 $Y=1.885 $X2=0 $Y2=0
cc_383 N_C_c_432_n N_VPWR_c_787_n 0.0044313f $X=2.43 $Y=1.885 $X2=0 $Y2=0
cc_384 N_C_c_422_n N_VPWR_c_787_n 0.0044313f $X=3.88 $Y=1.885 $X2=0 $Y2=0
cc_385 N_C_c_434_n N_VPWR_c_788_n 0.00320914f $X=4.9 $Y=1.885 $X2=0 $Y2=0
cc_386 N_C_c_435_n N_VPWR_c_788_n 0.00320914f $X=5.35 $Y=1.885 $X2=0 $Y2=0
cc_387 N_C_c_432_n N_VPWR_c_776_n 0.00853368f $X=2.43 $Y=1.885 $X2=0 $Y2=0
cc_388 N_C_c_422_n N_VPWR_c_776_n 0.00854258f $X=3.88 $Y=1.885 $X2=0 $Y2=0
cc_389 N_C_c_434_n N_VPWR_c_776_n 0.00401319f $X=4.9 $Y=1.885 $X2=0 $Y2=0
cc_390 N_C_c_435_n N_VPWR_c_776_n 0.00401319f $X=5.35 $Y=1.885 $X2=0 $Y2=0
cc_391 N_C_c_432_n N_A_501_392#_c_916_n 0.00351786f $X=2.43 $Y=1.885 $X2=0 $Y2=0
cc_392 N_C_c_422_n N_A_501_392#_c_914_n 0.00395612f $X=3.88 $Y=1.885 $X2=0 $Y2=0
cc_393 N_C_c_432_n N_A_501_392#_c_915_n 0.00369135f $X=2.43 $Y=1.885 $X2=0 $Y2=0
cc_394 N_C_c_422_n N_A_501_392#_c_926_n 0.00354606f $X=3.88 $Y=1.885 $X2=0 $Y2=0
cc_395 N_C_c_434_n N_A_905_392#_c_945_n 0.00937718f $X=4.9 $Y=1.885 $X2=0 $Y2=0
cc_396 N_C_c_435_n N_A_905_392#_c_945_n 0.0103693f $X=5.35 $Y=1.885 $X2=0 $Y2=0
cc_397 N_C_c_434_n N_A_905_392#_c_941_n 0.00633305f $X=4.9 $Y=1.885 $X2=0 $Y2=0
cc_398 N_C_c_435_n N_A_905_392#_c_941_n 8.31475e-19 $X=5.35 $Y=1.885 $X2=0 $Y2=0
cc_399 N_C_c_434_n N_A_905_392#_c_942_n 8.31475e-19 $X=4.9 $Y=1.885 $X2=0 $Y2=0
cc_400 N_C_c_435_n N_A_905_392#_c_942_n 0.00645035f $X=5.35 $Y=1.885 $X2=0 $Y2=0
cc_401 N_C_c_421_n N_VGND_c_1027_n 0.00600873f $X=2.52 $Y=0.18 $X2=0 $Y2=0
cc_402 N_C_c_420_n N_VGND_c_1028_n 0.00640572f $X=3.88 $Y=0.18 $X2=0 $Y2=0
cc_403 N_C_M1017_g N_VGND_c_1028_n 0.00661284f $X=3.955 $Y=0.71 $X2=0 $Y2=0
cc_404 N_C_c_421_n N_VGND_c_1034_n 0.0393818f $X=2.52 $Y=0.18 $X2=0 $Y2=0
cc_405 N_C_c_420_n N_VGND_c_1042_n 0.0359131f $X=3.88 $Y=0.18 $X2=0 $Y2=0
cc_406 N_C_c_421_n N_VGND_c_1042_n 0.00912007f $X=2.52 $Y=0.18 $X2=0 $Y2=0
cc_407 N_C_c_430_n N_A_504_125#_M1030_d 0.00277483f $X=3.747 $Y=1.215 $X2=0
+ $Y2=0
cc_408 N_C_M1007_g N_A_504_125#_c_1145_n 0.00853196f $X=2.445 $Y=0.945 $X2=0
+ $Y2=0
cc_409 N_C_c_420_n N_A_504_125#_c_1146_n 0.009817f $X=3.88 $Y=0.18 $X2=0 $Y2=0
cc_410 N_C_M1007_g N_A_504_125#_c_1147_n 0.00609242f $X=2.445 $Y=0.945 $X2=0
+ $Y2=0
cc_411 N_C_c_420_n N_A_504_125#_c_1147_n 0.00635148f $X=3.88 $Y=0.18 $X2=0 $Y2=0
cc_412 N_C_c_420_n N_A_504_125#_c_1148_n 0.007046f $X=3.88 $Y=0.18 $X2=0 $Y2=0
cc_413 N_C_M1017_g N_A_504_125#_c_1148_n 0.00379633f $X=3.955 $Y=0.71 $X2=0
+ $Y2=0
cc_414 N_C_c_426_n N_A_906_78#_M1004_d 0.00205112f $X=4.755 $Y=1.215 $X2=-0.19
+ $Y2=-0.245
cc_415 N_C_M1002_g N_A_906_78#_c_1179_n 0.00156411f $X=4.965 $Y=0.915 $X2=0
+ $Y2=0
cc_416 N_C_M1008_g N_A_906_78#_c_1179_n 0.00307819f $X=5.395 $Y=0.915 $X2=0
+ $Y2=0
cc_417 N_C_M1002_g N_A_906_78#_c_1180_n 4.53718e-19 $X=4.965 $Y=0.915 $X2=0
+ $Y2=0
cc_418 N_C_M1008_g N_A_906_78#_c_1180_n 0.00833548f $X=5.395 $Y=0.915 $X2=0
+ $Y2=0
cc_419 N_C_M1002_g N_A_906_78#_c_1181_n 0.00204725f $X=4.965 $Y=0.915 $X2=0
+ $Y2=0
cc_420 N_A_219_392#_c_591_n N_VPWR_M1029_s 0.00559435f $X=2.99 $Y=2.3 $X2=0
+ $Y2=0
cc_421 N_A_219_392#_c_596_n N_VPWR_M1027_d 0.00692629f $X=4.96 $Y=2.3 $X2=0
+ $Y2=0
cc_422 N_A_219_392#_c_572_n N_VPWR_c_778_n 0.00451331f $X=1.252 $Y=2.045 $X2=0
+ $Y2=0
cc_423 N_A_219_392#_c_591_n N_VPWR_c_779_n 0.019282f $X=2.99 $Y=2.3 $X2=0 $Y2=0
cc_424 N_A_219_392#_c_596_n N_VPWR_c_780_n 0.0248957f $X=4.96 $Y=2.3 $X2=0 $Y2=0
cc_425 N_A_219_392#_c_567_n N_VPWR_c_781_n 0.00857122f $X=6.305 $Y=1.765 $X2=0
+ $Y2=0
cc_426 N_A_219_392#_c_573_n N_VPWR_c_781_n 0.00127934f $X=5.475 $Y=1.97 $X2=0
+ $Y2=0
cc_427 N_A_219_392#_c_563_n N_VPWR_c_781_n 0.0149363f $X=6.985 $Y=1.51 $X2=0
+ $Y2=0
cc_428 N_A_219_392#_c_627_n N_VPWR_c_781_n 0.0144107f $X=5.125 $Y=2.215 $X2=0
+ $Y2=0
cc_429 N_A_219_392#_c_566_n N_VPWR_c_781_n 0.00102184f $X=7.655 $Y=1.555 $X2=0
+ $Y2=0
cc_430 N_A_219_392#_c_567_n N_VPWR_c_782_n 0.00445602f $X=6.305 $Y=1.765 $X2=0
+ $Y2=0
cc_431 N_A_219_392#_c_568_n N_VPWR_c_782_n 0.00445602f $X=6.755 $Y=1.765 $X2=0
+ $Y2=0
cc_432 N_A_219_392#_c_568_n N_VPWR_c_783_n 0.00595264f $X=6.755 $Y=1.765 $X2=0
+ $Y2=0
cc_433 N_A_219_392#_c_569_n N_VPWR_c_783_n 0.0124472f $X=7.205 $Y=1.765 $X2=0
+ $Y2=0
cc_434 N_A_219_392#_c_570_n N_VPWR_c_783_n 5.69946e-19 $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_435 N_A_219_392#_c_569_n N_VPWR_c_785_n 6.1988e-19 $X=7.205 $Y=1.765 $X2=0
+ $Y2=0
cc_436 N_A_219_392#_c_570_n N_VPWR_c_785_n 0.0181898f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_437 N_A_219_392#_c_566_n N_VPWR_c_785_n 4.41799e-19 $X=7.655 $Y=1.555 $X2=0
+ $Y2=0
cc_438 N_A_219_392#_c_569_n N_VPWR_c_789_n 0.00413917f $X=7.205 $Y=1.765 $X2=0
+ $Y2=0
cc_439 N_A_219_392#_c_570_n N_VPWR_c_789_n 0.00413917f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_440 N_A_219_392#_c_567_n N_VPWR_c_776_n 0.00857585f $X=6.305 $Y=1.765 $X2=0
+ $Y2=0
cc_441 N_A_219_392#_c_568_n N_VPWR_c_776_n 0.00857589f $X=6.755 $Y=1.765 $X2=0
+ $Y2=0
cc_442 N_A_219_392#_c_569_n N_VPWR_c_776_n 0.00817726f $X=7.205 $Y=1.765 $X2=0
+ $Y2=0
cc_443 N_A_219_392#_c_570_n N_VPWR_c_776_n 0.00817726f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_444 N_A_219_392#_c_572_n N_A_119_392#_M1014_d 0.00206372f $X=1.252 $Y=2.045
+ $X2=-0.19 $Y2=-0.245
cc_445 N_A_219_392#_c_591_n N_A_119_392#_M1022_s 0.00907415f $X=2.99 $Y=2.3
+ $X2=0 $Y2=0
cc_446 N_A_219_392#_c_572_n N_A_119_392#_c_894_n 0.00756635f $X=1.252 $Y=2.045
+ $X2=0 $Y2=0
cc_447 N_A_219_392#_M1011_d N_A_119_392#_c_888_n 0.00197722f $X=1.095 $Y=1.96
+ $X2=0 $Y2=0
cc_448 N_A_219_392#_c_687_p N_A_119_392#_c_888_n 0.014173f $X=1.245 $Y=2.57
+ $X2=0 $Y2=0
cc_449 N_A_219_392#_c_591_n N_A_119_392#_c_888_n 0.0032335f $X=2.99 $Y=2.3 $X2=0
+ $Y2=0
cc_450 N_A_219_392#_c_597_n N_A_119_392#_c_888_n 4.1793e-19 $X=1.252 $Y=2.3
+ $X2=0 $Y2=0
cc_451 N_A_219_392#_c_591_n N_A_119_392#_c_892_n 0.0168928f $X=2.99 $Y=2.3 $X2=0
+ $Y2=0
cc_452 N_A_219_392#_c_591_n N_A_501_392#_M1012_s 0.00395925f $X=2.99 $Y=2.3
+ $X2=-0.19 $Y2=-0.245
cc_453 N_A_219_392#_c_596_n N_A_501_392#_M1005_s 0.00494496f $X=4.96 $Y=2.3
+ $X2=0 $Y2=0
cc_454 N_A_219_392#_c_591_n N_A_501_392#_c_916_n 0.0168119f $X=2.99 $Y=2.3 $X2=0
+ $Y2=0
cc_455 N_A_219_392#_M1001_d N_A_501_392#_c_914_n 0.00250873f $X=2.955 $Y=1.96
+ $X2=0 $Y2=0
cc_456 N_A_219_392#_c_591_n N_A_501_392#_c_914_n 0.00365467f $X=2.99 $Y=2.3
+ $X2=0 $Y2=0
cc_457 N_A_219_392#_c_594_n N_A_501_392#_c_914_n 0.0185388f $X=3.155 $Y=2.65
+ $X2=0 $Y2=0
cc_458 N_A_219_392#_c_596_n N_A_501_392#_c_914_n 0.00365467f $X=4.96 $Y=2.3
+ $X2=0 $Y2=0
cc_459 N_A_219_392#_c_596_n N_A_501_392#_c_926_n 0.0197899f $X=4.96 $Y=2.3 $X2=0
+ $Y2=0
cc_460 N_A_219_392#_c_596_n N_A_905_392#_M1006_d 0.00879078f $X=4.96 $Y=2.3
+ $X2=-0.19 $Y2=-0.245
cc_461 N_A_219_392#_c_627_n N_A_905_392#_M1018_s 0.00337882f $X=5.125 $Y=2.215
+ $X2=0 $Y2=0
cc_462 N_A_219_392#_M1015_d N_A_905_392#_c_945_n 0.00510213f $X=4.975 $Y=1.96
+ $X2=0 $Y2=0
cc_463 N_A_219_392#_c_596_n N_A_905_392#_c_945_n 0.00809975f $X=4.96 $Y=2.3
+ $X2=0 $Y2=0
cc_464 N_A_219_392#_c_627_n N_A_905_392#_c_945_n 0.0206694f $X=5.125 $Y=2.215
+ $X2=0 $Y2=0
cc_465 N_A_219_392#_c_596_n N_A_905_392#_c_941_n 0.0165436f $X=4.96 $Y=2.3 $X2=0
+ $Y2=0
cc_466 N_A_219_392#_c_627_n N_A_905_392#_c_942_n 0.0040151f $X=5.125 $Y=2.215
+ $X2=0 $Y2=0
cc_467 N_A_219_392#_c_567_n N_X_c_973_n 0.00284497f $X=6.305 $Y=1.765 $X2=0
+ $Y2=0
cc_468 N_A_219_392#_c_568_n N_X_c_973_n 4.27055e-19 $X=6.755 $Y=1.765 $X2=0
+ $Y2=0
cc_469 N_A_219_392#_c_563_n N_X_c_973_n 0.0219683f $X=6.985 $Y=1.51 $X2=0 $Y2=0
cc_470 N_A_219_392#_c_566_n N_X_c_973_n 0.00654661f $X=7.655 $Y=1.555 $X2=0
+ $Y2=0
cc_471 N_A_219_392#_c_567_n N_X_c_970_n 0.010008f $X=6.305 $Y=1.765 $X2=0 $Y2=0
cc_472 N_A_219_392#_c_568_n N_X_c_970_n 0.0119295f $X=6.755 $Y=1.765 $X2=0 $Y2=0
cc_473 N_A_219_392#_c_569_n N_X_c_970_n 7.34739e-19 $X=7.205 $Y=1.765 $X2=0
+ $Y2=0
cc_474 N_A_219_392#_c_557_n N_X_c_967_n 0.0120699f $X=6.805 $Y=1.345 $X2=0 $Y2=0
cc_475 N_A_219_392#_c_558_n N_X_c_967_n 0.014204f $X=7.235 $Y=1.345 $X2=0 $Y2=0
cc_476 N_A_219_392#_c_559_n N_X_c_967_n 0.0140021f $X=7.665 $Y=1.345 $X2=0 $Y2=0
cc_477 N_A_219_392#_c_563_n N_X_c_967_n 0.0289012f $X=6.985 $Y=1.51 $X2=0 $Y2=0
cc_478 N_A_219_392#_c_566_n N_X_c_967_n 0.0046356f $X=7.655 $Y=1.555 $X2=0 $Y2=0
cc_479 N_A_219_392#_c_563_n N_X_c_986_n 0.0187104f $X=6.985 $Y=1.51 $X2=0 $Y2=0
cc_480 N_A_219_392#_c_566_n N_X_c_986_n 0.00325866f $X=7.655 $Y=1.555 $X2=0
+ $Y2=0
cc_481 N_A_219_392#_c_568_n N_X_c_988_n 0.0119563f $X=6.755 $Y=1.765 $X2=0 $Y2=0
cc_482 N_A_219_392#_c_569_n N_X_c_988_n 0.0145869f $X=7.205 $Y=1.765 $X2=0 $Y2=0
cc_483 N_A_219_392#_c_563_n N_X_c_988_n 0.0290464f $X=6.985 $Y=1.51 $X2=0 $Y2=0
cc_484 N_A_219_392#_c_566_n N_X_c_988_n 0.00779721f $X=7.655 $Y=1.555 $X2=0
+ $Y2=0
cc_485 N_A_219_392#_c_569_n N_X_c_971_n 0.00186003f $X=7.205 $Y=1.765 $X2=0
+ $Y2=0
cc_486 N_A_219_392#_c_570_n N_X_c_971_n 0.00146913f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_487 N_A_219_392#_c_563_n N_X_c_971_n 0.00160647f $X=6.985 $Y=1.51 $X2=0 $Y2=0
cc_488 N_A_219_392#_c_566_n N_X_c_971_n 0.0101615f $X=7.655 $Y=1.555 $X2=0 $Y2=0
cc_489 N_A_219_392#_c_569_n N_X_c_972_n 0.00424451f $X=7.205 $Y=1.765 $X2=0
+ $Y2=0
cc_490 N_A_219_392#_c_570_n N_X_c_972_n 0.00334744f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_491 N_A_219_392#_c_566_n N_X_c_968_n 0.0196476f $X=7.655 $Y=1.555 $X2=0 $Y2=0
cc_492 N_A_219_392#_c_563_n N_X_c_999_n 0.0128914f $X=6.985 $Y=1.51 $X2=0 $Y2=0
cc_493 N_A_219_392#_c_566_n N_X_c_999_n 0.00780004f $X=7.655 $Y=1.555 $X2=0
+ $Y2=0
cc_494 N_A_219_392#_c_559_n X 0.0116155f $X=7.665 $Y=1.345 $X2=0 $Y2=0
cc_495 N_A_219_392#_c_563_n X 0.00383354f $X=6.985 $Y=1.51 $X2=0 $Y2=0
cc_496 N_A_219_392#_c_595_n N_VGND_M1017_d 0.00488427f $X=5.095 $Y=0.875 $X2=0
+ $Y2=0
cc_497 N_A_219_392#_c_560_n N_VGND_c_1026_n 0.00804752f $X=0.88 $Y=0.96 $X2=0
+ $Y2=0
cc_498 N_A_219_392#_c_561_n N_VGND_c_1026_n 0.0137788f $X=0.88 $Y=1.875 $X2=0
+ $Y2=0
cc_499 N_A_219_392#_c_595_n N_VGND_c_1028_n 0.0204925f $X=5.095 $Y=0.875 $X2=0
+ $Y2=0
cc_500 N_A_219_392#_c_556_n N_VGND_c_1029_n 0.00178995f $X=6.335 $Y=1.345 $X2=0
+ $Y2=0
cc_501 N_A_219_392#_c_563_n N_VGND_c_1029_n 0.0211465f $X=6.985 $Y=1.51 $X2=0
+ $Y2=0
cc_502 N_A_219_392#_c_566_n N_VGND_c_1029_n 0.00148787f $X=7.655 $Y=1.555 $X2=0
+ $Y2=0
cc_503 N_A_219_392#_c_556_n N_VGND_c_1030_n 4.3896e-19 $X=6.335 $Y=1.345 $X2=0
+ $Y2=0
cc_504 N_A_219_392#_c_557_n N_VGND_c_1030_n 0.00830759f $X=6.805 $Y=1.345 $X2=0
+ $Y2=0
cc_505 N_A_219_392#_c_558_n N_VGND_c_1030_n 0.0106161f $X=7.235 $Y=1.345 $X2=0
+ $Y2=0
cc_506 N_A_219_392#_c_559_n N_VGND_c_1030_n 0.0013836f $X=7.665 $Y=1.345 $X2=0
+ $Y2=0
cc_507 N_A_219_392#_c_558_n N_VGND_c_1032_n 0.0013836f $X=7.235 $Y=1.345 $X2=0
+ $Y2=0
cc_508 N_A_219_392#_c_559_n N_VGND_c_1032_n 0.0116796f $X=7.665 $Y=1.345 $X2=0
+ $Y2=0
cc_509 N_A_219_392#_c_556_n N_VGND_c_1036_n 0.00490845f $X=6.335 $Y=1.345 $X2=0
+ $Y2=0
cc_510 N_A_219_392#_c_557_n N_VGND_c_1036_n 0.00407914f $X=6.805 $Y=1.345 $X2=0
+ $Y2=0
cc_511 N_A_219_392#_c_558_n N_VGND_c_1037_n 0.00407914f $X=7.235 $Y=1.345 $X2=0
+ $Y2=0
cc_512 N_A_219_392#_c_559_n N_VGND_c_1037_n 0.00407914f $X=7.665 $Y=1.345 $X2=0
+ $Y2=0
cc_513 N_A_219_392#_c_556_n N_VGND_c_1042_n 0.00506877f $X=6.335 $Y=1.345 $X2=0
+ $Y2=0
cc_514 N_A_219_392#_c_557_n N_VGND_c_1042_n 0.00425776f $X=6.805 $Y=1.345 $X2=0
+ $Y2=0
cc_515 N_A_219_392#_c_558_n N_VGND_c_1042_n 0.00425776f $X=7.235 $Y=1.345 $X2=0
+ $Y2=0
cc_516 N_A_219_392#_c_559_n N_VGND_c_1042_n 0.00425776f $X=7.665 $Y=1.345 $X2=0
+ $Y2=0
cc_517 N_A_219_392#_c_560_n N_VGND_c_1042_n 8.2431e-19 $X=0.88 $Y=0.96 $X2=0
+ $Y2=0
cc_518 N_A_219_392#_c_595_n N_VGND_c_1042_n 0.0140608f $X=5.095 $Y=0.875 $X2=0
+ $Y2=0
cc_519 N_A_219_392#_c_560_n N_A_114_125#_M1013_s 0.00391632f $X=0.88 $Y=0.96
+ $X2=-0.19 $Y2=-0.245
cc_520 N_A_219_392#_c_561_n N_A_114_125#_M1013_s 0.00431621f $X=0.88 $Y=1.875
+ $X2=-0.19 $Y2=-0.245
cc_521 N_A_219_392#_c_560_n N_A_114_125#_c_1119_n 0.0304906f $X=0.88 $Y=0.96
+ $X2=0 $Y2=0
cc_522 N_A_219_392#_c_560_n N_A_114_125#_c_1120_n 0.0149198f $X=0.88 $Y=0.96
+ $X2=0 $Y2=0
cc_523 N_A_219_392#_c_560_n N_A_114_125#_c_1121_n 0.0143885f $X=0.88 $Y=0.96
+ $X2=0 $Y2=0
cc_524 N_A_219_392#_c_595_n N_A_504_125#_M1030_d 0.00709487f $X=5.095 $Y=0.875
+ $X2=0 $Y2=0
cc_525 N_A_219_392#_c_564_n N_A_504_125#_c_1145_n 0.0128619f $X=3.15 $Y=0.78
+ $X2=0 $Y2=0
cc_526 N_A_219_392#_c_595_n N_A_504_125#_c_1146_n 0.00580283f $X=5.095 $Y=0.875
+ $X2=0 $Y2=0
cc_527 N_A_219_392#_c_564_n N_A_504_125#_c_1146_n 0.0185913f $X=3.15 $Y=0.78
+ $X2=0 $Y2=0
cc_528 N_A_219_392#_c_595_n N_A_504_125#_c_1148_n 0.0245465f $X=5.095 $Y=0.875
+ $X2=0 $Y2=0
cc_529 N_A_219_392#_c_564_n N_A_504_125#_c_1148_n 0.00111461f $X=3.15 $Y=0.78
+ $X2=0 $Y2=0
cc_530 N_A_219_392#_c_595_n N_A_906_78#_M1004_d 0.00493556f $X=5.095 $Y=0.875
+ $X2=-0.19 $Y2=-0.245
cc_531 N_A_219_392#_c_562_n N_A_906_78#_M1008_s 0.00171779f $X=5.475 $Y=1.675
+ $X2=0 $Y2=0
cc_532 N_A_219_392#_c_595_n N_A_906_78#_c_1179_n 0.00775961f $X=5.095 $Y=0.875
+ $X2=0 $Y2=0
cc_533 N_A_219_392#_c_565_n N_A_906_78#_c_1179_n 0.0129666f $X=5.18 $Y=0.76
+ $X2=0 $Y2=0
cc_534 N_A_219_392#_c_562_n N_A_906_78#_c_1180_n 0.00497798f $X=5.475 $Y=1.675
+ $X2=0 $Y2=0
cc_535 N_A_219_392#_c_563_n N_A_906_78#_c_1180_n 0.00856441f $X=6.985 $Y=1.51
+ $X2=0 $Y2=0
cc_536 N_A_219_392#_c_595_n N_A_906_78#_c_1181_n 0.0201615f $X=5.095 $Y=0.875
+ $X2=0 $Y2=0
cc_537 N_VPWR_c_778_n N_A_119_392#_c_894_n 0.0462323f $X=0.295 $Y=2.105 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_779_n N_A_119_392#_c_888_n 0.0123076f $X=2.15 $Y=2.72 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_786_n N_A_119_392#_c_888_n 0.0621395f $X=2.06 $Y=3.33 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_776_n N_A_119_392#_c_888_n 0.0346106f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_778_n N_A_119_392#_c_889_n 0.012272f $X=0.295 $Y=2.105 $X2=0
+ $Y2=0
cc_542 N_VPWR_c_786_n N_A_119_392#_c_889_n 0.0236039f $X=2.06 $Y=3.33 $X2=0
+ $Y2=0
cc_543 N_VPWR_c_776_n N_A_119_392#_c_889_n 0.012761f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_544 N_VPWR_c_779_n N_A_119_392#_c_892_n 0.0235051f $X=2.15 $Y=2.72 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_780_n N_A_501_392#_c_914_n 0.0119239f $X=4.155 $Y=2.72 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_787_n N_A_501_392#_c_914_n 0.0654114f $X=3.99 $Y=3.33 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_776_n N_A_501_392#_c_914_n 0.0365591f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_779_n N_A_501_392#_c_915_n 0.0117551f $X=2.15 $Y=2.72 $X2=0
+ $Y2=0
cc_549 N_VPWR_c_787_n N_A_501_392#_c_915_n 0.0230852f $X=3.99 $Y=3.33 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_776_n N_A_501_392#_c_915_n 0.0126044f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_788_n N_A_905_392#_c_945_n 0.00940922f $X=5.94 $Y=3.33 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_776_n N_A_905_392#_c_945_n 0.0153148f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_553 N_VPWR_c_780_n N_A_905_392#_c_941_n 0.0153184f $X=4.155 $Y=2.72 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_788_n N_A_905_392#_c_941_n 0.0140716f $X=5.94 $Y=3.33 $X2=0
+ $Y2=0
cc_555 N_VPWR_c_776_n N_A_905_392#_c_941_n 0.0117933f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_781_n N_A_905_392#_c_942_n 0.0285262f $X=6.025 $Y=2.105 $X2=0
+ $Y2=0
cc_557 N_VPWR_c_788_n N_A_905_392#_c_942_n 0.0140716f $X=5.94 $Y=3.33 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_776_n N_A_905_392#_c_942_n 0.0117933f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_781_n N_X_c_970_n 0.0360825f $X=6.025 $Y=2.105 $X2=0 $Y2=0
cc_560 N_VPWR_c_782_n N_X_c_970_n 0.014552f $X=6.895 $Y=3.33 $X2=0 $Y2=0
cc_561 N_VPWR_c_783_n N_X_c_970_n 0.0533352f $X=6.98 $Y=2.35 $X2=0 $Y2=0
cc_562 N_VPWR_c_776_n N_X_c_970_n 0.0119791f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_563 N_VPWR_M1003_d N_X_c_988_n 0.0037816f $X=6.83 $Y=1.84 $X2=0 $Y2=0
cc_564 N_VPWR_c_783_n N_X_c_988_n 0.0154248f $X=6.98 $Y=2.35 $X2=0 $Y2=0
cc_565 N_VPWR_c_785_n N_X_c_971_n 0.00162356f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_566 N_VPWR_c_783_n N_X_c_972_n 0.0507202f $X=6.98 $Y=2.35 $X2=0 $Y2=0
cc_567 N_VPWR_c_785_n N_X_c_972_n 0.0628522f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_568 N_VPWR_c_789_n N_X_c_972_n 0.00749631f $X=7.715 $Y=3.33 $X2=0 $Y2=0
cc_569 N_VPWR_c_776_n N_X_c_972_n 0.0062048f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_570 N_VPWR_c_785_n N_X_c_968_n 0.0287715f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_571 N_VPWR_c_785_n N_X_c_1015_n 0.0123817f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_572 N_VPWR_c_778_n N_VGND_c_1026_n 0.00901122f $X=0.295 $Y=2.105 $X2=0 $Y2=0
cc_573 N_X_c_967_n N_VGND_M1021_d 0.00330483f $X=7.805 $Y=1.09 $X2=0 $Y2=0
cc_574 N_X_c_967_n N_VGND_M1031_d 0.00286145f $X=7.805 $Y=1.09 $X2=0 $Y2=0
cc_575 X N_VGND_M1031_d 9.02712e-19 $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_576 N_X_c_966_n N_VGND_c_1029_n 0.00126499f $X=6.59 $Y=0.64 $X2=0 $Y2=0
cc_577 N_X_c_966_n N_VGND_c_1030_n 0.0136308f $X=6.59 $Y=0.64 $X2=0 $Y2=0
cc_578 N_X_c_967_n N_VGND_c_1030_n 0.0170777f $X=7.805 $Y=1.09 $X2=0 $Y2=0
cc_579 N_X_c_967_n N_VGND_c_1032_n 0.023215f $X=7.805 $Y=1.09 $X2=0 $Y2=0
cc_580 N_X_c_966_n N_VGND_c_1036_n 0.00734888f $X=6.59 $Y=0.64 $X2=0 $Y2=0
cc_581 N_X_c_966_n N_VGND_c_1042_n 0.00845298f $X=6.59 $Y=0.64 $X2=0 $Y2=0
cc_582 N_VGND_c_1027_n N_A_114_125#_c_1119_n 0.0130055f $X=2.23 $Y=0.78 $X2=0
+ $Y2=0
cc_583 N_VGND_c_1033_n N_A_114_125#_c_1119_n 0.0633823f $X=2.145 $Y=0 $X2=0
+ $Y2=0
cc_584 N_VGND_c_1042_n N_A_114_125#_c_1119_n 0.0341125f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_585 N_VGND_c_1027_n N_A_114_125#_c_1120_n 0.0256104f $X=2.23 $Y=0.78 $X2=0
+ $Y2=0
cc_586 N_VGND_c_1026_n N_A_114_125#_c_1121_n 0.0269092f $X=0.28 $Y=0.77 $X2=0
+ $Y2=0
cc_587 N_VGND_c_1033_n N_A_114_125#_c_1121_n 0.0210718f $X=2.145 $Y=0 $X2=0
+ $Y2=0
cc_588 N_VGND_c_1042_n N_A_114_125#_c_1121_n 0.0111709f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_589 N_VGND_c_1027_n N_A_504_125#_c_1145_n 0.0251774f $X=2.23 $Y=0.78 $X2=0
+ $Y2=0
cc_590 N_VGND_c_1034_n N_A_504_125#_c_1146_n 0.0369458f $X=4.005 $Y=0 $X2=0
+ $Y2=0
cc_591 N_VGND_c_1042_n N_A_504_125#_c_1146_n 0.0203602f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_592 N_VGND_c_1027_n N_A_504_125#_c_1147_n 0.0130055f $X=2.23 $Y=0.78 $X2=0
+ $Y2=0
cc_593 N_VGND_c_1034_n N_A_504_125#_c_1147_n 0.0261721f $X=4.005 $Y=0 $X2=0
+ $Y2=0
cc_594 N_VGND_c_1042_n N_A_504_125#_c_1147_n 0.013484f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_595 N_VGND_c_1028_n N_A_504_125#_c_1148_n 0.0176811f $X=4.17 $Y=0.535 $X2=0
+ $Y2=0
cc_596 N_VGND_c_1034_n N_A_504_125#_c_1148_n 0.0210718f $X=4.005 $Y=0 $X2=0
+ $Y2=0
cc_597 N_VGND_c_1042_n N_A_504_125#_c_1148_n 0.0111709f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_598 N_VGND_c_1029_n N_A_906_78#_c_1179_n 0.0133372f $X=6.12 $Y=0.64 $X2=0
+ $Y2=0
cc_599 N_VGND_c_1035_n N_A_906_78#_c_1179_n 0.0617759f $X=5.955 $Y=0 $X2=0 $Y2=0
cc_600 N_VGND_c_1042_n N_A_906_78#_c_1179_n 0.0317974f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_601 N_VGND_c_1029_n N_A_906_78#_c_1180_n 0.0256144f $X=6.12 $Y=0.64 $X2=0
+ $Y2=0
cc_602 N_VGND_c_1028_n N_A_906_78#_c_1181_n 0.0192332f $X=4.17 $Y=0.535 $X2=0
+ $Y2=0
cc_603 N_VGND_c_1035_n N_A_906_78#_c_1181_n 0.0213621f $X=5.955 $Y=0 $X2=0 $Y2=0
cc_604 N_VGND_c_1042_n N_A_906_78#_c_1181_n 0.0110227f $X=7.92 $Y=0 $X2=0 $Y2=0
