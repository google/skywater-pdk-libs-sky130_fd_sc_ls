* File: sky130_fd_sc_ls__dlrtn_1.spice
* Created: Wed Sep  2 11:03:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dlrtn_1.pex.spice"
.subckt sky130_fd_sc_ls__dlrtn_1  VNB VPB D GATE_N RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_D_M1012_g N_A_27_136#_M1012_s VNB NSHORT L=0.15 W=0.55
+ AD=0.171076 AS=0.15675 PD=1.27054 PS=1.67 NRD=55.86 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1001 N_A_232_98#_M1001_d N_GATE_N_M1001_g N_VGND_M1012_d VNB NSHORT L=0.15
+ W=0.74 AD=0.1961 AS=0.230174 PD=2.01 PS=1.70946 NRD=0 NRS=41.52 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_232_98#_M1015_g N_A_357_392#_M1015_s VNB NSHORT L=0.15
+ W=0.74 AD=0.426921 AS=0.2109 PD=2.06449 PS=2.05 NRD=84.624 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1011 A_681_74# N_A_27_136#_M1011_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.369229 PD=0.88 PS=1.78551 NRD=12.18 NRS=15.936 M=1 R=4.26667
+ SA=75001.3 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1017 N_A_654_392#_M1017_d N_A_232_98#_M1017_g A_681_74# VNB NSHORT L=0.15
+ W=0.64 AD=0.115623 AS=0.0768 PD=1.16528 PS=0.88 NRD=8.436 NRS=12.18 M=1
+ R=4.26667 SA=75001.7 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1007 A_854_74# N_A_357_392#_M1007_g N_A_654_392#_M1017_d VNB NSHORT L=0.15
+ W=0.42 AD=0.05775 AS=0.0758774 PD=0.695 PS=0.764717 NRD=23.568 NRS=0 M=1 R=2.8
+ SA=75002.1 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_897_406#_M1004_g A_854_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.1239 AS=0.05775 PD=1.43 PS=0.695 NRD=1.428 NRS=23.568 M=1 R=2.8
+ SA=75002.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 A_1139_74# N_A_654_392#_M1013_g N_A_897_406#_M1013_s VNB NSHORT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_RESET_B_M1008_g A_1139_74# VNB NSHORT L=0.15 W=0.74
+ AD=0.163525 AS=0.0888 PD=1.185 PS=0.98 NRD=12.972 NRS=10.536 M=1 R=4.93333
+ SA=75000.6 SB=75000.9 A=0.111 P=1.78 MULT=1
MM1014 N_Q_M1014_d N_A_897_406#_M1014_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2701 AS=0.163525 PD=2.21 PS=1.185 NRD=12.972 NRS=12.972 M=1 R=4.93333
+ SA=75001.2 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_D_M1000_g N_A_27_136#_M1000_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.198125 AS=0.2478 PD=1.315 PS=2.27 NRD=22.261 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1019 N_A_232_98#_M1019_d N_GATE_N_M1019_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.198125 PD=2.27 PS=1.315 NRD=2.3443 NRS=22.261 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_A_232_98#_M1009_g N_A_357_392#_M1009_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.225202 AS=0.2478 PD=1.46087 PS=2.27 NRD=49.9592 NRS=2.3443
+ M=1 R=5.6 SA=75000.2 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1005 A_570_392# N_A_27_136#_M1005_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.268098 PD=1.27 PS=1.73913 NRD=15.7403 NRS=19.6803 M=1 R=6.66667
+ SA=75000.8 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1002 N_A_654_392#_M1002_d N_A_357_392#_M1002_g A_570_392# VPB PHIGHVT L=0.15
+ W=1 AD=0.283732 AS=0.135 PD=2.17606 PS=1.27 NRD=2.9353 NRS=15.7403 M=1
+ R=6.66667 SA=75001.2 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1003 A_793_508# N_A_232_98#_M1003_g N_A_654_392#_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.11235 AS=0.119168 PD=0.955 PS=0.913944 NRD=99.6623 NRS=107.286 M=1
+ R=2.8 SA=75001.8 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1018 N_VPWR_M1018_d N_A_897_406#_M1018_g A_793_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.132152 AS=0.11235 PD=1.11507 PS=0.955 NRD=4.6886 NRS=99.6623 M=1 R=2.8
+ SA=75002.4 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1010 N_A_897_406#_M1010_d N_A_654_392#_M1010_g N_VPWR_M1018_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.235 AS=0.314648 PD=1.47 PS=2.65493 NRD=18.715 NRS=1.9503 M=1
+ R=6.66667 SA=75001.2 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1016 N_VPWR_M1016_d N_RESET_B_M1016_g N_A_897_406#_M1010_d VPB PHIGHVT L=0.15
+ W=1 AD=0.224717 AS=0.235 PD=1.46698 PS=1.47 NRD=19.0302 NRS=18.715 M=1
+ R=6.66667 SA=75001.8 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1006 N_Q_M1006_d N_A_897_406#_M1006_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.251683 PD=2.83 PS=1.64302 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=14.0988 P=18.88
*
.include "sky130_fd_sc_ls__dlrtn_1.pxi.spice"
*
.ends
*
*
