# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__maj3_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__maj3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.180000 1.795000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.305000 1.245000 2.975000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.215000 1.245000 3.715000 1.300000 ;
        RECT 3.215000 1.300000 4.535000 1.630000 ;
        RECT 3.215000 1.630000 3.715000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 0.350000 0.895000 1.130000 ;
        RECT 0.555000 1.130000 0.725000 1.820000 ;
        RECT 0.555000 1.820000 0.915000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.135000  0.085000 0.385000 1.130000 ;
      RECT 0.135000  1.820000 0.385000 3.245000 ;
      RECT 0.895000  1.320000 1.255000 1.650000 ;
      RECT 1.075000  0.085000 1.795000 1.010000 ;
      RECT 1.085000  1.650000 1.255000 1.780000 ;
      RECT 1.085000  1.780000 2.135000 1.950000 ;
      RECT 1.085000  2.120000 1.780000 3.245000 ;
      RECT 1.965000  0.350000 2.760000 0.905000 ;
      RECT 1.965000  0.905000 4.660000 1.075000 ;
      RECT 1.965000  1.075000 2.135000 1.780000 ;
      RECT 1.965000  1.950000 4.685000 2.120000 ;
      RECT 1.965000  2.120000 2.785000 2.755000 ;
      RECT 3.340000  0.085000 3.840000 0.680000 ;
      RECT 3.485000  2.290000 3.815000 3.245000 ;
      RECT 4.330000  0.350000 4.660000 0.905000 ;
      RECT 4.330000  1.075000 4.660000 1.130000 ;
      RECT 4.355000  1.820000 4.685000 1.950000 ;
      RECT 4.355000  2.120000 4.685000 2.860000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_ls__maj3_2
