* NGSPICE file created from sky130_fd_sc_ls__dfrtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
M1000 VGND a_2010_409# Q VNB nshort w=740000u l=150000u
+  ad=2.10185e+12p pd=1.715e+07u as=4.847e+11p ps=4.27e+06u
M1001 a_1350_392# a_494_392# a_834_355# VNB nshort w=740000u l=150000u
+  ad=4.58e+11p pd=3.28e+06u as=9.435e+11p ps=4.03e+06u
M1002 VGND RESET_B a_124_78# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1003 a_2010_409# a_1350_392# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=3.136e+12p ps=2.402e+07u
M1004 a_494_392# a_299_392# VGND VNB nshort w=740000u l=150000u
+  ad=2.0255e+11p pd=2.07e+06u as=0p ps=0u
M1005 VPWR a_2010_409# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=7.224e+11p ps=5.77e+06u
M1006 a_699_463# a_494_392# a_37_78# VPB phighvt w=420000u l=150000u
+  ad=2.478e+11p pd=2.86e+06u as=2.478e+11p ps=2.86e+06u
M1007 a_1627_493# a_494_392# a_1350_392# VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=6.724e+11p ps=4.47e+06u
M1008 VGND CLK a_299_392# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.4175e+11p ps=2.14e+06u
M1009 a_834_355# a_699_463# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR CLK a_299_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=3.223e+11p ps=2.75e+06u
M1011 a_789_463# a_299_392# a_699_463# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1012 a_124_78# D a_37_78# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1013 a_2010_409# a_1350_392# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1014 a_1678_395# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1015 a_834_355# a_699_463# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1016 VGND a_2010_409# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_494_392# a_299_392# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1018 a_890_138# a_834_355# a_812_138# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.008e+11p ps=1.32e+06u
M1019 Q a_2010_409# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_1678_395# a_1647_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1021 a_37_78# D VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR RESET_B a_37_78# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_1350_392# a_1678_395# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1350_392# a_299_392# a_834_355# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_699_463# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_834_355# a_789_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1678_395# a_1350_392# a_1827_81# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1028 Q a_2010_409# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND RESET_B a_890_138# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_1350_392# a_2010_409# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_2010_409# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Q a_2010_409# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1827_81# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_812_138# a_494_392# a_699_463# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1035 a_1647_81# a_299_392# a_1350_392# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Q a_2010_409# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_699_463# a_299_392# a_37_78# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR a_1678_395# a_1627_493# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

