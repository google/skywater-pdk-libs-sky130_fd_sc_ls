* File: sky130_fd_sc_ls__sedfxtp_2.pex.spice
* Created: Wed Sep  2 11:29:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%D 2 3 5 8 12 13 18 19 21 23
c42 23 0 2.2081e-19 $X=0.525 $Y=1.99
c43 18 0 1.59585e-19 $X=0.525 $Y=1.145
r44 21 23 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.825
+ $X2=0.525 $Y2=1.99
r45 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.825 $X2=0.525 $Y2=1.825
r46 18 21 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=0.525 $Y=1.145
+ $X2=0.525 $Y2=1.825
r47 18 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.145 $X2=0.525 $Y2=1.145
r48 13 22 4.85239 $w=3.78e-07 $l=1.6e-07 $layer=LI1_cond $X=0.615 $Y=1.665
+ $X2=0.615 $Y2=1.825
r49 12 13 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.615 $Y=1.295
+ $X2=0.615 $Y2=1.665
r50 12 19 4.54912 $w=3.78e-07 $l=1.5e-07 $layer=LI1_cond $X=0.615 $Y=1.295
+ $X2=0.615 $Y2=1.145
r51 11 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=0.98
+ $X2=0.525 $Y2=1.145
r52 8 11 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.615 $Y=0.58 $X2=0.615
+ $Y2=0.98
r53 3 5 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.57 $Y=2.245
+ $X2=0.57 $Y2=2.64
r54 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.57 $Y=2.155 $X2=0.57
+ $Y2=2.245
r55 2 23 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.57 $Y=2.155
+ $X2=0.57 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%A_180_290# 1 2 7 9 12 14 18 19 20 21 22 23
+ 26 30 32 34 44
c107 44 0 1.26127e-19 $X=2.425 $Y=1.685
c108 34 0 7.02076e-20 $X=2.22 $Y=1.685
c109 32 0 7.48038e-20 $X=2.22 $Y=1.95
c110 23 0 3.52195e-20 $X=1.305 $Y=2.035
c111 21 0 1.59585e-19 $X=1.305 $Y=1.065
c112 19 0 1.74672e-19 $X=1.14 $Y=1.615
r113 35 44 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=2.22 $Y=1.685
+ $X2=2.425 $Y2=1.685
r114 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.22
+ $Y=1.685 $X2=2.22 $Y2=1.685
r115 32 37 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.22 $Y=2.035
+ $X2=1.895 $Y2=2.035
r116 32 34 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.22 $Y=1.95
+ $X2=2.22 $Y2=1.685
r117 28 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=2.12
+ $X2=1.895 $Y2=2.035
r118 28 30 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.895 $Y=2.12
+ $X2=1.895 $Y2=2.515
r119 24 26 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=1.74 $Y=0.98
+ $X2=1.74 $Y2=0.775
r120 22 37 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=2.035
+ $X2=1.895 $Y2=2.035
r121 22 23 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.81 $Y=2.035
+ $X2=1.305 $Y2=2.035
r122 20 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.615 $Y=1.065
+ $X2=1.74 $Y2=0.98
r123 20 21 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.615 $Y=1.065
+ $X2=1.305 $Y2=1.065
r124 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.14
+ $Y=1.615 $X2=1.14 $Y2=1.615
r125 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.14 $Y=1.95
+ $X2=1.305 $Y2=2.035
r126 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.14 $Y=1.95
+ $X2=1.14 $Y2=1.615
r127 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.14 $Y=1.15
+ $X2=1.305 $Y2=1.065
r128 15 18 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.14 $Y=1.15
+ $X2=1.14 $Y2=1.615
r129 14 19 41.6085 $w=4.05e-07 $l=3.03e-07 $layer=POLY_cond $X=1.102 $Y=1.918
+ $X2=1.102 $Y2=1.615
r130 10 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.425 $Y=1.52
+ $X2=2.425 $Y2=1.685
r131 10 12 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=2.425 $Y=1.52
+ $X2=2.425 $Y2=0.775
r132 7 14 49.5642 $w=3.18e-07 $l=3.78884e-07 $layer=POLY_cond $X=0.99 $Y=2.245
+ $X2=1.102 $Y2=1.918
r133 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.99 $Y=2.245
+ $X2=0.99 $Y2=2.64
r134 2 30 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=2.315 $X2=1.895 $Y2=2.515
r135 1 26 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.635
+ $Y=0.565 $X2=1.78 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%DE 3 5 6 10 11 12 13 15 16 18 19 21 23 25
+ 27 28 31 32 33
c93 33 0 7.48038e-20 $X=1.68 $Y=1.65
c94 32 0 1.3237e-19 $X=1.68 $Y=1.485
c95 25 0 7.02076e-20 $X=1.995 $Y=1.135
r96 31 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.485
+ $X2=1.68 $Y2=1.65
r97 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.485 $X2=1.68 $Y2=1.485
r98 28 32 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=1.485
r99 21 23 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.8 $Y=2.24 $X2=2.8
+ $Y2=2.635
r100 20 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=2.165
+ $X2=2.12 $Y2=2.165
r101 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.725 $Y=2.165
+ $X2=2.8 $Y2=2.24
r102 19 20 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.725 $Y=2.165
+ $X2=2.195 $Y2=2.165
r103 16 27 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.24
+ $X2=2.12 $Y2=2.165
r104 16 18 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.12 $Y=2.24
+ $X2=2.12 $Y2=2.635
r105 13 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.995 $Y=1.06
+ $X2=1.995 $Y2=1.135
r106 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.995 $Y=1.06
+ $X2=1.995 $Y2=0.775
r107 11 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.045 $Y=2.165
+ $X2=2.12 $Y2=2.165
r108 11 12 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.045 $Y=2.165
+ $X2=1.815 $Y2=2.165
r109 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.74 $Y=2.09
+ $X2=1.815 $Y2=2.165
r110 10 33 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.74 $Y=2.09
+ $X2=1.74 $Y2=1.65
r111 7 25 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=1.68 $Y=1.135
+ $X2=1.995 $Y2=1.135
r112 7 31 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=1.68 $Y=1.21
+ $X2=1.68 $Y2=1.485
r113 5 7 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.135
+ $X2=1.68 $Y2=1.135
r114 5 6 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.515 $Y=1.135
+ $X2=1.08 $Y2=1.135
r115 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.005 $Y=1.06
+ $X2=1.08 $Y2=1.135
r116 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.005 $Y=1.06
+ $X2=1.005 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%A_548_87# 1 2 9 12 13 15 16 18 19 20 21 23
+ 25 26 30 35 37 39 45 47 49 50 51 57 58 64 65
c252 50 0 1.30591e-19 $X=14.975 $Y=1.665
c253 49 0 1.70806e-19 $X=14.665 $Y=1.665
c254 25 0 3.76658e-20 $X=13.765 $Y=2.05
c255 13 0 1.85697e-19 $X=3.19 $Y=2.24
c256 12 0 1.26127e-19 $X=3.19 $Y=2.15
r257 63 65 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=2.905 $Y=1.68
+ $X2=3.19 $Y2=1.68
r258 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.905
+ $Y=1.68 $X2=2.905 $Y2=1.68
r259 60 63 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.815 $Y=1.68
+ $X2=2.905 $Y2=1.68
r260 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=1.665
+ $X2=15.12 $Y2=1.665
r261 54 64 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.64 $Y=1.68
+ $X2=2.905 $Y2=1.68
r262 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=1.665
r263 51 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.665
+ $X2=2.64 $Y2=1.665
r264 50 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.975 $Y=1.665
+ $X2=15.12 $Y2=1.665
r265 50 51 15.0866 $w=1.4e-07 $l=1.219e-05 $layer=MET1_cond $X=14.975 $Y=1.665
+ $X2=2.785 $Y2=1.665
r266 48 58 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=14.75 $Y=1.665
+ $X2=15.12 $Y2=1.665
r267 48 49 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.75 $Y=1.665
+ $X2=14.665 $Y2=1.665
r268 44 45 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=14.532 $Y=1.12
+ $X2=14.532 $Y2=1.29
r269 39 42 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=13.675 $Y=2.215
+ $X2=13.675 $Y2=2.385
r270 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.675
+ $Y=2.215 $X2=13.675 $Y2=2.215
r271 37 47 3.58051 $w=2.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=14.665 $Y=2.3
+ $X2=14.575 $Y2=2.385
r272 36 49 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=14.665 $Y=1.78
+ $X2=14.665 $Y2=1.665
r273 36 37 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=14.665 $Y=1.78
+ $X2=14.665 $Y2=2.3
r274 35 49 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=14.665 $Y=1.55
+ $X2=14.665 $Y2=1.665
r275 35 45 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=14.665 $Y=1.55
+ $X2=14.665 $Y2=1.29
r276 30 44 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=14.48 $Y=0.58
+ $X2=14.48 $Y2=1.12
r277 27 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.84 $Y=2.385
+ $X2=13.675 $Y2=2.385
r278 26 47 2.90867 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=14.4 $Y=2.385
+ $X2=14.575 $Y2=2.385
r279 26 27 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=14.4 $Y=2.385
+ $X2=13.84 $Y2=2.385
r280 25 40 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=13.765 $Y=2.05
+ $X2=13.675 $Y2=2.215
r281 24 25 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=13.765 $Y=1.015
+ $X2=13.765 $Y2=2.05
r282 21 40 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=13.63 $Y=2.465
+ $X2=13.675 $Y2=2.215
r283 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.63 $Y=2.465
+ $X2=13.63 $Y2=2.75
r284 19 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.69 $Y=0.94
+ $X2=13.765 $Y2=1.015
r285 19 20 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=13.69 $Y=0.94
+ $X2=13.235 $Y2=0.94
r286 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.16 $Y=0.865
+ $X2=13.235 $Y2=0.94
r287 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.16 $Y=0.865
+ $X2=13.16 $Y2=0.58
r288 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.19 $Y=2.24
+ $X2=3.19 $Y2=2.635
r289 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.19 $Y=2.15 $X2=3.19
+ $Y2=2.24
r290 11 65 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.845
+ $X2=3.19 $Y2=1.68
r291 11 12 118.556 $w=1.8e-07 $l=3.05e-07 $layer=POLY_cond $X=3.19 $Y=1.845
+ $X2=3.19 $Y2=2.15
r292 7 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=1.515
+ $X2=2.815 $Y2=1.68
r293 7 9 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.815 $Y=1.515
+ $X2=2.815 $Y2=0.775
r294 2 47 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=14.415
+ $Y=2.32 $X2=14.565 $Y2=2.465
r295 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=14.34
+ $Y=0.37 $X2=14.48 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%A_663_87# 1 2 7 9 10 11 12 14 17 18 21 22
+ 27 28 30 31 35 36 41 43 47
c110 41 0 1.05969e-19 $X=4.55 $Y=0.805
c111 12 0 1.43112e-19 $X=5.74 $Y=2.2
r112 44 47 5.10825 $w=4.78e-07 $l=2.05e-07 $layer=LI1_cond $X=4.21 $Y=2.495
+ $X2=4.415 $Y2=2.495
r113 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.785
+ $Y=1.58 $X2=5.785 $Y2=1.58
r114 33 35 14.5686 $w=2.63e-07 $l=3.35e-07 $layer=LI1_cond $X=5.752 $Y=1.915
+ $X2=5.752 $Y2=1.58
r115 32 43 2.40986 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=4.295 $Y=2
+ $X2=4.152 $Y2=2
r116 31 33 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=5.62 $Y=2
+ $X2=5.752 $Y2=1.915
r117 31 32 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=5.62 $Y=2
+ $X2=4.295 $Y2=2
r118 30 44 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=4.21 $Y=2.255
+ $X2=4.21 $Y2=2.495
r119 29 43 4.02809 $w=2.27e-07 $l=1.1025e-07 $layer=LI1_cond $X=4.21 $Y=2.085
+ $X2=4.152 $Y2=2
r120 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.21 $Y=2.085
+ $X2=4.21 $Y2=2.255
r121 27 28 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.13
+ $Y=1.78 $X2=4.13 $Y2=1.78
r122 25 43 4.02809 $w=2.27e-07 $l=8.5e-08 $layer=LI1_cond $X=4.152 $Y=1.915
+ $X2=4.152 $Y2=2
r123 25 27 5.45894 $w=2.83e-07 $l=1.35e-07 $layer=LI1_cond $X=4.152 $Y=1.915
+ $X2=4.152 $Y2=1.78
r124 24 27 31.1362 $w=2.83e-07 $l=7.7e-07 $layer=LI1_cond $X=4.152 $Y=1.01
+ $X2=4.152 $Y2=1.78
r125 21 22 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.13
+ $Y=0.42 $X2=4.13 $Y2=0.42
r126 19 41 11.3252 $w=4.03e-07 $l=3.98e-07 $layer=LI1_cond $X=4.152 $Y=0.807
+ $X2=4.55 $Y2=0.807
r127 19 24 2.81058 $w=2.85e-07 $l=2.03e-07 $layer=LI1_cond $X=4.152 $Y=0.807
+ $X2=4.152 $Y2=1.01
r128 19 21 7.48077 $w=2.83e-07 $l=1.85e-07 $layer=LI1_cond $X=4.152 $Y=0.605
+ $X2=4.152 $Y2=0.42
r129 18 36 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.785 $Y=1.92
+ $X2=5.785 $Y2=1.58
r130 16 28 99.6709 $w=3.3e-07 $l=5.7e-07 $layer=POLY_cond $X=4.13 $Y=1.21
+ $X2=4.13 $Y2=1.78
r131 16 17 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.13 $Y=1.21
+ $X2=4.13 $Y2=1.135
r132 15 22 111.911 $w=3.3e-07 $l=6.4e-07 $layer=POLY_cond $X=4.13 $Y=1.06
+ $X2=4.13 $Y2=0.42
r133 15 17 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.13 $Y=1.06
+ $X2=4.13 $Y2=1.135
r134 12 18 50.3582 $w=2.68e-07 $l=3.01662e-07 $layer=POLY_cond $X=5.74 $Y=2.2
+ $X2=5.785 $Y2=1.92
r135 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.74 $Y=2.2
+ $X2=5.74 $Y2=2.595
r136 10 17 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.965 $Y=1.135
+ $X2=4.13 $Y2=1.135
r137 10 11 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.965 $Y=1.135
+ $X2=3.465 $Y2=1.135
r138 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.39 $Y=1.06
+ $X2=3.465 $Y2=1.135
r139 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.39 $Y=1.06 $X2=3.39
+ $Y2=0.775
r140 2 47 600 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=2.275 $X2=4.415 $Y2=2.495
r141 1 41 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=4.405
+ $Y=0.625 $X2=4.55 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%SCD 3 6 7 9 10 13
c43 13 0 8.67074e-20 $X=5.245 $Y=1.58
c44 3 0 3.01793e-19 $X=5.265 $Y=0.835
r45 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.245 $Y=1.58
+ $X2=5.245 $Y2=1.745
r46 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.245 $Y=1.58
+ $X2=5.245 $Y2=1.415
r47 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.245
+ $Y=1.58 $X2=5.245 $Y2=1.58
r48 10 14 7.49192 $w=4.53e-07 $l=2.85e-07 $layer=LI1_cond $X=5.182 $Y=1.295
+ $X2=5.182 $Y2=1.58
r49 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.32 $Y=2.2 $X2=5.32
+ $Y2=2.595
r50 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.32 $Y=2.11 $X2=5.32
+ $Y2=2.2
r51 6 16 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=5.32 $Y=2.11
+ $X2=5.32 $Y2=1.745
r52 3 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.265 $Y=0.835
+ $X2=5.265 $Y2=1.415
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%SCE 1 3 4 5 7 8 11 15 16 17 20 22 25 26
c85 26 0 2.82531e-19 $X=4.67 $Y=1.345
c86 20 0 1.9935e-19 $X=5.625 $Y=0.835
r87 25 28 40.6969 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.672 $Y=1.345
+ $X2=4.672 $Y2=1.51
r88 25 27 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.672 $Y=1.345
+ $X2=4.672 $Y2=1.18
r89 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.67
+ $Y=1.345 $X2=4.67 $Y2=1.345
r90 22 26 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=4.56 $Y=1.345
+ $X2=4.67 $Y2=1.345
r91 18 20 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.625 $Y=0.255
+ $X2=5.625 $Y2=0.835
r92 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.55 $Y=0.18
+ $X2=5.625 $Y2=0.255
r93 16 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.55 $Y=0.18
+ $X2=4.84 $Y2=0.18
r94 15 27 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=4.765 $Y=0.835
+ $X2=4.765 $Y2=1.18
r95 12 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.765 $Y=0.255
+ $X2=4.84 $Y2=0.18
r96 12 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.765 $Y=0.255
+ $X2=4.765 $Y2=0.835
r97 9 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.64 $Y=2.99
+ $X2=4.64 $Y2=2.595
r98 8 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.64 $Y=2.2 $X2=4.64
+ $Y2=2.595
r99 7 8 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.64 $Y=2.11 $X2=4.64
+ $Y2=2.2
r100 7 28 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=4.64 $Y=2.11 $X2=4.64
+ $Y2=1.51
r101 4 9 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=4.55 $Y=3.105
+ $X2=4.64 $Y2=2.99
r102 4 5 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=4.55 $Y=3.105
+ $X2=3.715 $Y2=3.105
r103 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.64 $Y=3.03
+ $X2=3.715 $Y2=3.105
r104 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.64 $Y=3.03
+ $X2=3.64 $Y2=2.635
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%CLK 1 3 4 6 7
c34 7 0 1.22168e-20 $X=6.48 $Y=1.295
r35 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.56
+ $Y=1.385 $X2=6.56 $Y2=1.385
r36 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.56 $Y=1.295 $X2=6.56
+ $Y2=1.385
r37 4 10 65.7037 $w=3.49e-07 $l=4.22137e-07 $layer=POLY_cond $X=6.755 $Y=1.745
+ $X2=6.62 $Y2=1.385
r38 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.755 $Y=1.745
+ $X2=6.755 $Y2=2.38
r39 1 10 38.7725 $w=3.49e-07 $l=1.67481e-07 $layer=POLY_cond $X=6.625 $Y=1.22
+ $X2=6.62 $Y2=1.385
r40 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.625 $Y=1.22 $X2=6.625
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%A_1538_74# 1 2 7 9 10 12 15 18 19 21 24 26
+ 27 28 33 34 38 41 42 43 45 46 47 49 52 53 55 57 58 61 62 63 66 68 69 73
c237 73 0 2.65373e-20 $X=13.285 $Y=1.42
c238 61 0 1.50148e-19 $X=8.84 $Y=2.185
c239 53 0 1.80054e-19 $X=12.205 $Y=1.635
c240 33 0 1.39112e-19 $X=8.73 $Y=1.82
c241 19 0 1.48476e-19 $X=13.21 $Y=2.465
r242 73 86 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.285 $Y=1.42
+ $X2=13.285 $Y2=1.585
r243 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.285
+ $Y=1.42 $X2=13.285 $Y2=1.42
r244 69 72 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=13.285 $Y=1.275
+ $X2=13.285 $Y2=1.42
r245 66 77 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=9.49 $Y=1.18
+ $X2=9.285 $Y2=1.18
r246 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.49
+ $Y=1.18 $X2=9.49 $Y2=1.18
r247 62 65 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=9.49 $Y=0.935
+ $X2=9.49 $Y2=1.18
r248 62 63 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=9.49 $Y=0.935
+ $X2=9.49 $Y2=0.85
r249 61 76 52.3552 $w=2.9e-07 $l=3.15e-07 $layer=POLY_cond $X=8.84 $Y=2.242
+ $X2=9.155 $Y2=2.242
r250 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.84
+ $Y=2.185 $X2=8.84 $Y2=2.185
r251 58 60 3.16509 $w=4.24e-07 $l=1.1e-07 $layer=LI1_cond $X=8.73 $Y=2.085
+ $X2=8.84 $Y2=2.085
r252 56 68 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.37 $Y=1.275
+ $X2=12.205 $Y2=1.275
r253 55 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.12 $Y=1.275
+ $X2=13.285 $Y2=1.275
r254 55 56 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=13.12 $Y=1.275
+ $X2=12.37 $Y2=1.275
r255 53 82 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.205 $Y=1.635
+ $X2=12.205 $Y2=1.47
r256 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.205
+ $Y=1.635 $X2=12.205 $Y2=1.635
r257 50 68 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.205 $Y=1.36
+ $X2=12.205 $Y2=1.275
r258 50 52 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=12.205 $Y=1.36
+ $X2=12.205 $Y2=1.635
r259 49 68 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=12.125 $Y=1.19
+ $X2=12.205 $Y2=1.275
r260 48 49 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=12.125 $Y=1.02
+ $X2=12.125 $Y2=1.19
r261 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.04 $Y=0.935
+ $X2=12.125 $Y2=1.02
r262 46 47 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=12.04 $Y=0.935
+ $X2=11.465 $Y2=0.935
r263 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.38 $Y=0.85
+ $X2=11.465 $Y2=0.935
r264 44 45 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=11.38 $Y=0.425
+ $X2=11.38 $Y2=0.85
r265 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.295 $Y=0.34
+ $X2=11.38 $Y2=0.425
r266 42 43 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.295 $Y=0.34
+ $X2=10.705 $Y2=0.34
r267 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.62 $Y=0.425
+ $X2=10.705 $Y2=0.34
r268 40 41 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=10.62 $Y=0.425
+ $X2=10.62 $Y2=0.85
r269 39 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.655 $Y=0.935
+ $X2=9.49 $Y2=0.935
r270 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.535 $Y=0.935
+ $X2=10.62 $Y2=0.85
r271 38 39 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=10.535 $Y=0.935
+ $X2=9.655 $Y2=0.935
r272 36 63 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.41 $Y=0.425
+ $X2=9.41 $Y2=0.85
r273 35 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.815 $Y=0.34
+ $X2=8.73 $Y2=0.34
r274 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.325 $Y=0.34
+ $X2=9.41 $Y2=0.425
r275 34 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.325 $Y=0.34
+ $X2=8.815 $Y2=0.34
r276 33 58 6.13403 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=8.73 $Y=1.82
+ $X2=8.73 $Y2=2.085
r277 32 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.73 $Y=0.425
+ $X2=8.73 $Y2=0.34
r278 32 33 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=8.73 $Y=0.425
+ $X2=8.73 $Y2=1.82
r279 28 58 2.60462 $w=4.24e-07 $l=1.16619e-07 $layer=LI1_cond $X=8.645 $Y=2.01
+ $X2=8.73 $Y2=2.085
r280 28 30 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=8.645 $Y=2.01
+ $X2=8.37 $Y2=2.01
r281 26 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.645 $Y=0.34
+ $X2=8.73 $Y2=0.34
r282 26 27 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=8.645 $Y=0.34
+ $X2=7.995 $Y2=0.34
r283 22 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.83 $Y=0.425
+ $X2=7.995 $Y2=0.34
r284 22 24 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.83 $Y=0.425
+ $X2=7.83 $Y2=0.515
r285 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.21 $Y=2.465
+ $X2=13.21 $Y2=2.75
r286 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=13.21 $Y=2.375
+ $X2=13.21 $Y2=2.465
r287 18 86 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=13.21 $Y=2.375
+ $X2=13.21 $Y2=1.585
r288 15 82 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=12.295 $Y=0.69
+ $X2=12.295 $Y2=1.47
r289 10 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.285 $Y=1.015
+ $X2=9.285 $Y2=1.18
r290 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.285 $Y=1.015
+ $X2=9.285 $Y2=0.695
r291 7 76 18.1727 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=9.155 $Y=2.465
+ $X2=9.155 $Y2=2.242
r292 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.155 $Y=2.465
+ $X2=9.155 $Y2=2.75
r293 2 30 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=8.22
+ $Y=1.84 $X2=8.37 $Y2=2.01
r294 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.69
+ $Y=0.37 $X2=7.83 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%A_1340_74# 1 2 11 13 15 17 18 22 24 27 28
+ 30 31 33 36 38 39 42 45 46 49 50 55 56 59 65
c188 59 0 1.50148e-19 $X=9.69 $Y=2.185
c189 56 0 1.22168e-20 $X=7.45 $Y=1.695
c190 46 0 1.48476e-19 $X=12.56 $Y=2.475
c191 27 0 1.39112e-19 $X=9.58 $Y=2.02
r192 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.745
+ $Y=1.635 $X2=12.745 $Y2=1.635
r193 62 65 5.12197 $w=2.23e-07 $l=1e-07 $layer=LI1_cond $X=12.645 $Y=1.642
+ $X2=12.745 $Y2=1.642
r194 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.69
+ $Y=2.185 $X2=9.69 $Y2=2.185
r195 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.45
+ $Y=1.695 $X2=7.45 $Y2=1.695
r196 53 55 8.3904 $w=6.68e-07 $l=4.7e-07 $layer=LI1_cond $X=6.98 $Y=1.865
+ $X2=7.45 $Y2=1.865
r197 48 62 2.38091 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=12.645 $Y=1.755
+ $X2=12.645 $Y2=1.642
r198 48 49 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=12.645 $Y=1.755
+ $X2=12.645 $Y2=2.39
r199 47 59 12.3706 $w=2.86e-07 $l=3.69188e-07 $layer=LI1_cond $X=9.885 $Y=2.475
+ $X2=9.705 $Y2=2.185
r200 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.56 $Y=2.475
+ $X2=12.645 $Y2=2.39
r201 46 47 174.519 $w=1.68e-07 $l=2.675e-06 $layer=LI1_cond $X=12.56 $Y=2.475
+ $X2=9.885 $Y2=2.475
r202 45 53 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=6.98 $Y=1.53
+ $X2=6.98 $Y2=1.865
r203 45 50 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.98 $Y=1.53
+ $X2=6.98 $Y2=1.01
r204 40 50 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=6.87 $Y=0.815
+ $X2=6.87 $Y2=1.01
r205 40 42 8.86495 $w=3.88e-07 $l=3e-07 $layer=LI1_cond $X=6.87 $Y=0.815
+ $X2=6.87 $Y2=0.515
r206 34 66 38.5562 $w=2.99e-07 $l=1.77059e-07 $layer=POLY_cond $X=12.77 $Y=1.47
+ $X2=12.745 $Y2=1.635
r207 34 36 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=12.77 $Y=1.47
+ $X2=12.77 $Y2=0.58
r208 31 66 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=12.67 $Y=1.885
+ $X2=12.745 $Y2=1.635
r209 31 33 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.67 $Y=1.885
+ $X2=12.67 $Y2=2.46
r210 28 60 56.6494 $w=3.06e-07 $l=3.15278e-07 $layer=POLY_cond $X=9.605 $Y=2.465
+ $X2=9.68 $Y2=2.185
r211 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.605 $Y=2.465
+ $X2=9.605 $Y2=2.75
r212 27 60 38.535 $w=3.06e-07 $l=2.09105e-07 $layer=POLY_cond $X=9.58 $Y=2.02
+ $X2=9.68 $Y2=2.185
r213 26 27 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=9.58 $Y=1.765
+ $X2=9.58 $Y2=2.02
r214 25 39 17.0838 $w=1.85e-07 $l=9.08295e-08 $layer=POLY_cond $X=8.68 $Y=1.69
+ $X2=8.605 $Y2=1.655
r215 24 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.505 $Y=1.69
+ $X2=9.58 $Y2=1.765
r216 24 25 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=9.505 $Y=1.69
+ $X2=8.68 $Y2=1.69
r217 20 39 8.32657 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=8.605 $Y=1.545
+ $X2=8.605 $Y2=1.655
r218 20 22 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=8.605 $Y=1.545
+ $X2=8.605 $Y2=0.695
r219 19 38 14.6817 $w=2.2e-07 $l=7.5e-08 $layer=POLY_cond $X=8.22 $Y=1.655
+ $X2=8.145 $Y2=1.655
r220 18 39 17.0838 $w=1.85e-07 $l=7.5e-08 $layer=POLY_cond $X=8.53 $Y=1.655
+ $X2=8.605 $Y2=1.655
r221 18 19 90.4236 $w=2.2e-07 $l=3.1e-07 $layer=POLY_cond $X=8.53 $Y=1.655
+ $X2=8.22 $Y2=1.655
r222 15 38 10.8713 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=8.145 $Y=1.765
+ $X2=8.145 $Y2=1.655
r223 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.145 $Y=1.765
+ $X2=8.145 $Y2=2.4
r224 14 56 8.65449 $w=2.2e-07 $l=2.06961e-07 $layer=POLY_cond $X=7.69 $Y=1.655
+ $X2=7.487 $Y2=1.647
r225 13 38 14.6817 $w=2.2e-07 $l=7.5e-08 $layer=POLY_cond $X=8.07 $Y=1.655
+ $X2=8.145 $Y2=1.655
r226 13 14 110.842 $w=2.2e-07 $l=3.8e-07 $layer=POLY_cond $X=8.07 $Y=1.655
+ $X2=7.69 $Y2=1.655
r227 9 56 16.755 $w=2.77e-07 $l=1.77088e-07 $layer=POLY_cond $X=7.615 $Y=1.53
+ $X2=7.487 $Y2=1.647
r228 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.615 $Y=1.53
+ $X2=7.615 $Y2=0.74
r229 2 53 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=6.83
+ $Y=1.82 $X2=6.98 $Y2=2
r230 1 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.7
+ $Y=0.37 $X2=6.84 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%A_1979_71# 1 2 9 12 13 15 18 19 20 22 23
+ 25 26 30 33 36 37 43 47 49 53
c106 36 0 1.80054e-19 $X=11.635 $Y=1.355
r107 45 47 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=10.915 $Y=2.135
+ $X2=11.04 $Y2=2.135
r108 41 53 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=10.08 $Y=1.34
+ $X2=10.155 $Y2=1.34
r109 41 50 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=10.08 $Y=1.34
+ $X2=9.97 $Y2=1.34
r110 40 43 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=10.08 $Y=1.34
+ $X2=10.245 $Y2=1.34
r111 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.08
+ $Y=1.34 $X2=10.08 $Y2=1.34
r112 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.635
+ $Y=1.355 $X2=11.635 $Y2=1.355
r113 34 49 2.53577 $w=3.3e-07 $l=3.22102e-07 $layer=LI1_cond $X=11.125 $Y=1.355
+ $X2=10.875 $Y2=1.19
r114 34 36 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=11.125 $Y=1.355
+ $X2=11.635 $Y2=1.355
r115 33 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.04 $Y=2.05
+ $X2=11.04 $Y2=2.135
r116 32 49 3.59786 $w=1.7e-07 $l=4.04166e-07 $layer=LI1_cond $X=11.04 $Y=1.52
+ $X2=10.875 $Y2=1.19
r117 32 33 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=11.04 $Y=1.52
+ $X2=11.04 $Y2=2.05
r118 28 49 3.59786 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=11 $Y=1.19
+ $X2=10.875 $Y2=1.19
r119 28 30 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=11 $Y=1.19 $X2=11
+ $Y2=0.81
r120 26 49 2.53577 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.875 $Y=1.275
+ $X2=10.875 $Y2=1.19
r121 26 43 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=10.875 $Y=1.275
+ $X2=10.245 $Y2=1.275
r122 23 25 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=11.935 $Y=1.11
+ $X2=11.935 $Y2=0.69
r123 20 22 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=11.71 $Y=1.885
+ $X2=11.71 $Y2=2.46
r124 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.71 $Y=1.795
+ $X2=11.71 $Y2=1.885
r125 18 23 40.1667 $w=2.7e-07 $l=3.76032e-07 $layer=POLY_cond $X=11.71 $Y=1.39
+ $X2=11.935 $Y2=1.11
r126 18 37 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=11.71 $Y=1.39
+ $X2=11.635 $Y2=1.39
r127 18 19 106.895 $w=1.8e-07 $l=2.75e-07 $layer=POLY_cond $X=11.71 $Y=1.52
+ $X2=11.71 $Y2=1.795
r128 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.155 $Y=2.465
+ $X2=10.155 $Y2=2.75
r129 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.155 $Y=2.375
+ $X2=10.155 $Y2=2.465
r130 11 53 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.155 $Y=1.505
+ $X2=10.155 $Y2=1.34
r131 11 12 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=10.155 $Y=1.505
+ $X2=10.155 $Y2=2.375
r132 7 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.97 $Y=1.175
+ $X2=9.97 $Y2=1.34
r133 7 9 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.97 $Y=1.175
+ $X2=9.97 $Y2=0.695
r134 2 45 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.765
+ $Y=1.99 $X2=10.915 $Y2=2.135
r135 1 30 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=10.82
+ $Y=0.37 $X2=10.96 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%A_1736_97# 1 2 7 9 12 16 20 21 26 27 30
r85 30 33 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=10.62 $Y=1.665
+ $X2=10.62 $Y2=1.745
r86 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.62
+ $Y=1.665 $X2=10.62 $Y2=1.665
r87 26 27 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=9.365 $Y=2.75
+ $X2=9.365 $Y2=2.52
r88 22 24 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=9.07 $Y=1.745 $X2=9.27
+ $Y2=1.745
r89 21 24 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=9.355 $Y=1.745
+ $X2=9.27 $Y2=1.745
r90 20 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.455 $Y=1.745
+ $X2=10.62 $Y2=1.745
r91 20 21 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=10.455 $Y=1.745
+ $X2=9.355 $Y2=1.745
r92 18 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.27 $Y=1.83
+ $X2=9.27 $Y2=1.745
r93 18 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.27 $Y=1.83 $X2=9.27
+ $Y2=2.52
r94 14 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.07 $Y=1.66
+ $X2=9.07 $Y2=1.745
r95 14 16 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=9.07 $Y=1.66 $X2=9.07
+ $Y2=0.76
r96 10 31 38.5818 $w=3.27e-07 $l=2.12238e-07 $layer=POLY_cond $X=10.745 $Y=1.5
+ $X2=10.637 $Y2=1.665
r97 10 12 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=10.745 $Y=1.5
+ $X2=10.745 $Y2=0.69
r98 7 31 51.1109 $w=3.27e-07 $l=2.75227e-07 $layer=POLY_cond $X=10.69 $Y=1.915
+ $X2=10.637 $Y2=1.665
r99 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.69 $Y=1.915
+ $X2=10.69 $Y2=2.41
r100 2 26 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=9.23
+ $Y=2.54 $X2=9.38 $Y2=2.75
r101 1 16 182 $w=1.7e-07 $l=5.09264e-07 $layer=licon1_NDIFF $count=1 $X=8.68
+ $Y=0.485 $X2=9.07 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%A_2474_74# 1 2 9 11 13 14 18 20 22 25 27
+ 29 31 32 35 39 41 42 45 47 48 50 51 54 56 57
c168 41 0 3.76658e-20 $X=13.62 $Y=0.935
r169 56 59 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=14.245 $Y=1.625
+ $X2=14.245 $Y2=1.84
r170 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=14.245
+ $Y=1.625 $X2=14.245 $Y2=1.625
r171 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.79 $Y=1.84
+ $X2=13.705 $Y2=1.84
r172 51 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.08 $Y=1.84
+ $X2=14.245 $Y2=1.84
r173 51 52 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=14.08 $Y=1.84
+ $X2=13.79 $Y2=1.84
r174 50 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.705 $Y=1.755
+ $X2=13.705 $Y2=1.84
r175 49 50 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=13.705 $Y=1.02
+ $X2=13.705 $Y2=1.755
r176 47 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.62 $Y=1.84
+ $X2=13.705 $Y2=1.84
r177 47 48 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.62 $Y=1.84
+ $X2=13.25 $Y2=1.84
r178 43 48 9.70699 $w=2.57e-07 $l=2.14126e-07 $layer=LI1_cond $X=13.075 $Y=1.927
+ $X2=13.25 $Y2=1.84
r179 43 45 21.4025 $w=3.48e-07 $l=6.5e-07 $layer=LI1_cond $X=13.075 $Y=2.1
+ $X2=13.075 $Y2=2.75
r180 41 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.62 $Y=0.935
+ $X2=13.705 $Y2=1.02
r181 41 42 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=13.62 $Y=0.935
+ $X2=12.72 $Y2=0.935
r182 37 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.555 $Y=0.85
+ $X2=12.72 $Y2=0.935
r183 37 39 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=12.555 $Y=0.85
+ $X2=12.555 $Y2=0.58
r184 35 36 8.95356 $w=3.23e-07 $l=6e-08 $layer=POLY_cond $X=15.755 $Y=1.562
+ $X2=15.815 $Y2=1.562
r185 34 35 60.4365 $w=3.23e-07 $l=4.05e-07 $layer=POLY_cond $X=15.35 $Y=1.562
+ $X2=15.755 $Y2=1.562
r186 33 34 3.73065 $w=3.23e-07 $l=2.5e-08 $layer=POLY_cond $X=15.325 $Y=1.562
+ $X2=15.35 $Y2=1.562
r187 32 57 54.4068 $w=3.5e-07 $l=3.3e-07 $layer=POLY_cond $X=14.255 $Y=1.955
+ $X2=14.255 $Y2=1.625
r188 30 57 2.47304 $w=3.5e-07 $l=1.5e-08 $layer=POLY_cond $X=14.255 $Y=1.61
+ $X2=14.255 $Y2=1.625
r189 30 31 20.4101 $w=2.5e-07 $l=2.38485e-07 $layer=POLY_cond $X=14.255 $Y=1.61
+ $X2=14.08 $Y2=1.46
r190 27 36 20.7134 $w=1.5e-07 $l=2.03e-07 $layer=POLY_cond $X=15.815 $Y=1.765
+ $X2=15.815 $Y2=1.562
r191 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=15.815 $Y=1.765
+ $X2=15.815 $Y2=2.4
r192 23 35 20.7134 $w=1.5e-07 $l=2.02e-07 $layer=POLY_cond $X=15.755 $Y=1.36
+ $X2=15.755 $Y2=1.562
r193 23 25 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=15.755 $Y=1.36
+ $X2=15.755 $Y2=0.74
r194 20 34 20.7134 $w=1.5e-07 $l=2.03e-07 $layer=POLY_cond $X=15.35 $Y=1.765
+ $X2=15.35 $Y2=1.562
r195 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=15.35 $Y=1.765
+ $X2=15.35 $Y2=2.4
r196 16 33 20.7134 $w=1.5e-07 $l=2.02e-07 $layer=POLY_cond $X=15.325 $Y=1.36
+ $X2=15.325 $Y2=1.562
r197 16 18 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=15.325 $Y=1.36
+ $X2=15.325 $Y2=0.74
r198 15 31 5.30422 $w=2.5e-07 $l=3.62284e-07 $layer=POLY_cond $X=14.43 $Y=1.485
+ $X2=14.08 $Y2=1.46
r199 14 33 13.7803 $w=3.23e-07 $l=1.08185e-07 $layer=POLY_cond $X=15.25 $Y=1.485
+ $X2=15.325 $Y2=1.562
r200 14 15 203.732 $w=2.5e-07 $l=8.2e-07 $layer=POLY_cond $X=15.25 $Y=1.485
+ $X2=14.43 $Y2=1.485
r201 11 32 49.5674 $w=2.82e-07 $l=3.29773e-07 $layer=POLY_cond $X=14.34 $Y=2.245
+ $X2=14.255 $Y2=1.955
r202 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=14.34 $Y=2.245
+ $X2=14.34 $Y2=2.64
r203 7 31 20.4101 $w=2.5e-07 $l=2.29619e-07 $layer=POLY_cond $X=14.265 $Y=1.36
+ $X2=14.08 $Y2=1.46
r204 7 9 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=14.265 $Y=1.36
+ $X2=14.265 $Y2=0.58
r205 2 45 600 $w=1.7e-07 $l=9.02053e-07 $layer=licon1_PDIFF $count=1 $X=12.745
+ $Y=1.96 $X2=12.985 $Y2=2.75
r206 1 39 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=12.37
+ $Y=0.37 $X2=12.555 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%A_40_464# 1 2 3 4 14 17 19 22 23 24 26 27
+ 28 30 33 36 40 42 46 50 52
c127 19 0 1.8559e-19 $X=1.47 $Y=2.375
r128 48 50 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.255 $Y=1.26
+ $X2=3.415 $Y2=1.26
r129 44 46 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.1 $Y=0.84
+ $X2=3.255 $Y2=0.84
r130 37 40 5.98039 $w=4.58e-07 $l=2.3e-07 $layer=LI1_cond $X=0.17 $Y=0.58
+ $X2=0.4 $Y2=0.58
r131 36 52 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.415 $Y=2.29
+ $X2=3.375 $Y2=2.375
r132 35 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=1.345
+ $X2=3.415 $Y2=1.26
r133 35 36 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=3.415 $Y=1.345
+ $X2=3.415 $Y2=2.29
r134 33 52 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=2.46
+ $X2=3.375 $Y2=2.375
r135 30 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.255 $Y=1.175
+ $X2=3.255 $Y2=1.26
r136 29 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=1.005
+ $X2=3.255 $Y2=0.84
r137 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.255 $Y=1.005
+ $X2=3.255 $Y2=1.175
r138 27 52 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.25 $Y=2.375
+ $X2=3.375 $Y2=2.375
r139 27 28 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.25 $Y=2.375
+ $X2=2.32 $Y2=2.375
r140 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.235 $Y=2.46
+ $X2=2.32 $Y2=2.375
r141 25 26 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.235 $Y=2.46
+ $X2=2.235 $Y2=2.905
r142 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.15 $Y=2.99
+ $X2=2.235 $Y2=2.905
r143 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.15 $Y=2.99
+ $X2=1.64 $Y2=2.99
r144 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.555 $Y=2.905
+ $X2=1.64 $Y2=2.99
r145 21 22 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.555 $Y=2.46
+ $X2=1.555 $Y2=2.905
r146 20 42 3.41642 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.51 $Y=2.375
+ $X2=0.297 $Y2=2.375
r147 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.47 $Y=2.375
+ $X2=1.555 $Y2=2.46
r148 19 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.47 $Y=2.375
+ $X2=0.51 $Y2=2.375
r149 15 42 3.17288 $w=2.97e-07 $l=8.5e-08 $layer=LI1_cond $X=0.297 $Y=2.46
+ $X2=0.297 $Y2=2.375
r150 15 17 0.135582 $w=4.23e-07 $l=5e-09 $layer=LI1_cond $X=0.297 $Y=2.46
+ $X2=0.297 $Y2=2.465
r151 14 42 3.17288 $w=2.97e-07 $l=1.64085e-07 $layer=LI1_cond $X=0.17 $Y=2.29
+ $X2=0.297 $Y2=2.375
r152 13 37 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.17 $Y=0.81 $X2=0.17
+ $Y2=0.58
r153 13 14 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=0.17 $Y=0.81
+ $X2=0.17 $Y2=2.29
r154 4 33 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.265
+ $Y=2.315 $X2=3.415 $Y2=2.46
r155 3 17 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.2
+ $Y=2.32 $X2=0.345 $Y2=2.465
r156 2 44 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=2.89
+ $Y=0.565 $X2=3.1 $Y2=0.84
r157 1 40 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.255
+ $Y=0.37 $X2=0.4 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49
+ 53 57 61 65 69 71 74 75 77 78 79 81 86 91 96 101 106 124 128 134 137 140 143
+ 146 149 152 156
c183 65 0 1.04054e-19 $X=15.125 $Y=2.035
c184 3 0 9.53964e-20 $X=4.715 $Y=2.275
r185 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=3.33
+ $X2=16.08 $Y2=3.33
r186 152 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r187 149 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r188 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r189 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r190 140 141 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r191 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r192 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r193 132 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=16.08 $Y2=3.33
r194 132 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=15.12 $Y2=3.33
r195 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r196 129 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.29 $Y=3.33
+ $X2=15.125 $Y2=3.33
r197 129 131 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=15.29 $Y=3.33
+ $X2=15.6 $Y2=3.33
r198 128 155 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=15.875 $Y=3.33
+ $X2=16.097 $Y2=3.33
r199 128 131 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=15.875 $Y=3.33
+ $X2=15.6 $Y2=3.33
r200 127 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r201 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r202 124 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.96 $Y=3.33
+ $X2=15.125 $Y2=3.33
r203 124 126 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=14.96 $Y=3.33
+ $X2=14.64 $Y2=3.33
r204 123 127 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.64 $Y2=3.33
r205 122 123 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r206 120 123 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=13.68 $Y2=3.33
r207 119 122 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=11.76 $Y=3.33
+ $X2=13.68 $Y2=3.33
r208 119 120 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r209 117 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r210 117 150 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.32 $Y2=3.33
r211 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r212 114 149 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.545 $Y=3.33
+ $X2=10.38 $Y2=3.33
r213 114 116 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=10.545 $Y=3.33
+ $X2=11.28 $Y2=3.33
r214 113 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r215 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r216 110 113 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.84 $Y2=3.33
r217 109 112 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=9.84 $Y2=3.33
r218 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r219 107 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.085 $Y=3.33
+ $X2=7.92 $Y2=3.33
r220 107 109 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.085 $Y=3.33
+ $X2=8.4 $Y2=3.33
r221 106 149 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.215 $Y=3.33
+ $X2=10.38 $Y2=3.33
r222 106 112 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.215 $Y=3.33
+ $X2=9.84 $Y2=3.33
r223 105 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r224 105 144 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r225 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r226 102 143 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=6.527 $Y2=3.33
r227 102 104 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=7.44 $Y2=3.33
r228 101 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=3.33
+ $X2=7.92 $Y2=3.33
r229 101 104 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.755 $Y=3.33
+ $X2=7.44 $Y2=3.33
r230 100 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r231 100 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r232 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r233 97 140 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.26 $Y=3.33
+ $X2=5.135 $Y2=3.33
r234 97 99 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.26 $Y=3.33 $X2=6
+ $Y2=3.33
r235 96 143 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=6.36 $Y=3.33
+ $X2=6.527 $Y2=3.33
r236 96 99 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.36 $Y=3.33 $X2=6
+ $Y2=3.33
r237 95 141 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r238 95 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r239 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r240 92 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=2.615 $Y2=3.33
r241 92 94 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=3.12 $Y2=3.33
r242 91 140 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.01 $Y=3.33
+ $X2=5.135 $Y2=3.33
r243 91 94 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=5.01 $Y=3.33
+ $X2=3.12 $Y2=3.33
r244 90 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r245 90 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r246 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r247 87 134 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.3 $Y=3.33
+ $X2=1.175 $Y2=3.33
r248 87 89 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.3 $Y=3.33 $X2=2.16
+ $Y2=3.33
r249 86 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.49 $Y=3.33
+ $X2=2.615 $Y2=3.33
r250 86 89 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.49 $Y=3.33
+ $X2=2.16 $Y2=3.33
r251 84 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r252 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r253 81 134 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.05 $Y=3.33
+ $X2=1.175 $Y2=3.33
r254 81 83 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.05 $Y=3.33
+ $X2=0.72 $Y2=3.33
r255 79 110 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=8.16 $Y=3.33
+ $X2=8.4 $Y2=3.33
r256 79 147 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=8.16 $Y=3.33
+ $X2=7.92 $Y2=3.33
r257 77 122 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=13.69 $Y=3.33
+ $X2=13.68 $Y2=3.33
r258 77 78 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=13.69 $Y=3.33
+ $X2=13.96 $Y2=3.33
r259 76 126 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=14.23 $Y=3.33
+ $X2=14.64 $Y2=3.33
r260 76 78 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=14.23 $Y=3.33
+ $X2=13.96 $Y2=3.33
r261 74 116 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=11.31 $Y=3.33
+ $X2=11.28 $Y2=3.33
r262 74 75 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=11.31 $Y=3.33
+ $X2=11.48 $Y2=3.33
r263 73 119 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=11.65 $Y=3.33
+ $X2=11.76 $Y2=3.33
r264 73 75 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=11.65 $Y=3.33
+ $X2=11.48 $Y2=3.33
r265 69 155 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=16.04 $Y=3.245
+ $X2=16.097 $Y2=3.33
r266 69 71 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=16.04 $Y=3.245
+ $X2=16.04 $Y2=2.405
r267 65 68 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=15.125 $Y=2.035
+ $X2=15.125 $Y2=2.815
r268 63 152 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.125 $Y=3.245
+ $X2=15.125 $Y2=3.33
r269 63 68 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=15.125 $Y=3.245
+ $X2=15.125 $Y2=2.815
r270 59 78 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=13.96 $Y=3.245
+ $X2=13.96 $Y2=3.33
r271 59 61 9.52433 $w=5.38e-07 $l=4.3e-07 $layer=LI1_cond $X=13.96 $Y=3.245
+ $X2=13.96 $Y2=2.815
r272 55 75 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=11.48 $Y=3.245
+ $X2=11.48 $Y2=3.33
r273 55 57 14.575 $w=3.38e-07 $l=4.3e-07 $layer=LI1_cond $X=11.48 $Y=3.245
+ $X2=11.48 $Y2=2.815
r274 51 149 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.38 $Y=3.245
+ $X2=10.38 $Y2=3.33
r275 51 53 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.38 $Y=3.245
+ $X2=10.38 $Y2=2.815
r276 47 146 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=3.33
r277 47 49 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=2.805
r278 43 143 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=6.527 $Y=3.245
+ $X2=6.527 $Y2=3.33
r279 43 45 15.4806 $w=3.33e-07 $l=4.5e-07 $layer=LI1_cond $X=6.527 $Y=3.245
+ $X2=6.527 $Y2=2.795
r280 39 140 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.135 $Y=3.245
+ $X2=5.135 $Y2=3.33
r281 39 41 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=5.135 $Y=3.245
+ $X2=5.135 $Y2=2.765
r282 35 137 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=3.245
+ $X2=2.615 $Y2=3.33
r283 35 37 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.615 $Y=3.245
+ $X2=2.615 $Y2=2.8
r284 31 134 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=3.245
+ $X2=1.175 $Y2=3.33
r285 31 33 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=1.175 $Y=3.245
+ $X2=1.175 $Y2=2.805
r286 10 71 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=15.89
+ $Y=1.84 $X2=16.04 $Y2=2.405
r287 9 68 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=14.98
+ $Y=1.84 $X2=15.125 $Y2=2.815
r288 9 65 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=14.98
+ $Y=1.84 $X2=15.125 $Y2=2.035
r289 8 61 600 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_PDIFF $count=1 $X=13.705
+ $Y=2.54 $X2=13.96 $Y2=2.815
r290 7 57 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=11.33
+ $Y=1.96 $X2=11.48 $Y2=2.815
r291 6 53 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=10.23
+ $Y=2.54 $X2=10.38 $Y2=2.815
r292 5 49 600 $w=1.7e-07 $l=1.03496e-06 $layer=licon1_PDIFF $count=1 $X=7.775
+ $Y=1.84 $X2=7.92 $Y2=2.805
r293 4 45 600 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=1.82 $X2=6.525 $Y2=2.795
r294 3 41 600 $w=1.7e-07 $l=6.52917e-07 $layer=licon1_PDIFF $count=1 $X=4.715
+ $Y=2.275 $X2=5.095 $Y2=2.765
r295 2 37 600 $w=1.7e-07 $l=6.47708e-07 $layer=licon1_PDIFF $count=1 $X=2.195
+ $Y=2.315 $X2=2.575 $Y2=2.8
r296 1 33 600 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=1 $X=1.065
+ $Y=2.32 $X2=1.215 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%A_693_113# 1 2 3 4 5 6 21 24 25 26 28 29
+ 30 35 38 39 40 41 45 47 51 54 57 59 62 65 67 68
c172 62 0 1.43112e-19 $X=6.012 $Y=2.255
c173 57 0 1.85697e-19 $X=3.81 $Y=2.295
c174 25 0 9.53964e-20 $X=4.67 $Y=2.99
r175 68 70 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=8.34 $Y=2.455
+ $X2=8.34 $Y2=2.605
r176 64 65 0.949071 $w=4.23e-07 $l=3.5e-08 $layer=LI1_cond $X=6.012 $Y=2.42
+ $X2=6.012 $Y2=2.455
r177 56 57 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=3.755 $Y=1.005
+ $X2=3.755 $Y2=2.295
r178 54 56 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.675 $Y=0.775
+ $X2=3.675 $Y2=1.005
r179 49 51 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=8.89 $Y=2.69 $X2=8.89
+ $Y2=2.75
r180 48 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.425 $Y=2.605
+ $X2=8.34 $Y2=2.605
r181 47 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.765 $Y=2.605
+ $X2=8.89 $Y2=2.69
r182 47 48 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=8.765 $Y=2.605
+ $X2=8.425 $Y2=2.605
r183 43 45 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=8.35 $Y=1.48
+ $X2=8.35 $Y2=0.76
r184 42 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.035 $Y=2.455
+ $X2=7.95 $Y2=2.455
r185 41 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.255 $Y=2.455
+ $X2=8.34 $Y2=2.455
r186 41 42 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.255 $Y=2.455
+ $X2=8.035 $Y2=2.455
r187 39 43 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.225 $Y=1.565
+ $X2=8.35 $Y2=1.48
r188 39 40 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=8.225 $Y=1.565
+ $X2=8.035 $Y2=1.565
r189 38 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.95 $Y=2.37
+ $X2=7.95 $Y2=2.455
r190 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.95 $Y=1.65
+ $X2=8.035 $Y2=1.565
r191 37 38 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=7.95 $Y=1.65
+ $X2=7.95 $Y2=2.37
r192 36 65 6.14847 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=6.225 $Y=2.455
+ $X2=6.012 $Y2=2.455
r193 35 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.865 $Y=2.455
+ $X2=7.95 $Y2=2.455
r194 35 36 106.995 $w=1.68e-07 $l=1.64e-06 $layer=LI1_cond $X=7.865 $Y=2.455
+ $X2=6.225 $Y2=2.455
r195 33 59 10.6395 $w=3.44e-07 $l=3.98748e-07 $layer=LI1_cond $X=6.14 $Y=1.065
+ $X2=5.84 $Y2=0.835
r196 33 62 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=6.14 $Y=1.065
+ $X2=6.14 $Y2=2.255
r197 29 64 2.1693 $w=4.23e-07 $l=8e-08 $layer=LI1_cond $X=6.012 $Y=2.34
+ $X2=6.012 $Y2=2.42
r198 29 62 6.59116 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=6.012 $Y=2.34
+ $X2=6.012 $Y2=2.255
r199 29 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.8 $Y=2.34 $X2=4.84
+ $Y2=2.34
r200 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.755 $Y=2.425
+ $X2=4.84 $Y2=2.34
r201 27 28 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.755 $Y=2.425
+ $X2=4.755 $Y2=2.905
r202 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.67 $Y=2.99
+ $X2=4.755 $Y2=2.905
r203 25 26 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.67 $Y=2.99
+ $X2=3.95 $Y2=2.99
r204 22 26 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.81 $Y=2.905
+ $X2=3.95 $Y2=2.99
r205 22 24 18.3156 $w=2.78e-07 $l=4.45e-07 $layer=LI1_cond $X=3.81 $Y=2.905
+ $X2=3.81 $Y2=2.46
r206 21 57 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=3.81 $Y=2.435
+ $X2=3.81 $Y2=2.295
r207 21 24 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.81 $Y=2.435
+ $X2=3.81 $Y2=2.46
r208 6 51 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=8.785
+ $Y=2.54 $X2=8.93 $Y2=2.75
r209 5 64 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=5.815
+ $Y=2.275 $X2=5.965 $Y2=2.42
r210 4 24 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.715
+ $Y=2.315 $X2=3.865 $Y2=2.46
r211 3 45 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=8.245
+ $Y=0.485 $X2=8.39 $Y2=0.76
r212 2 59 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.7
+ $Y=0.625 $X2=5.84 $Y2=0.835
r213 1 54 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=3.465
+ $Y=0.565 $X2=3.675 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%Q 1 2 9 12 15 17 18 19
r33 23 25 0.0398693 $w=5.98e-07 $l=2e-09 $layer=LI1_cond $X=15.58 $Y=1.85
+ $X2=15.582 $Y2=1.85
r34 18 19 9.56863 $w=5.98e-07 $l=4.8e-07 $layer=LI1_cond $X=15.6 $Y=1.85
+ $X2=16.08 $Y2=1.85
r35 18 25 0.358824 $w=5.98e-07 $l=1.8e-08 $layer=LI1_cond $X=15.6 $Y=1.85
+ $X2=15.582 $Y2=1.85
r36 13 25 6.03242 $w=2.45e-07 $l=3e-07 $layer=LI1_cond $X=15.582 $Y=2.15
+ $X2=15.582 $Y2=1.85
r37 13 15 12.23 $w=2.43e-07 $l=2.6e-07 $layer=LI1_cond $X=15.582 $Y=2.15
+ $X2=15.582 $Y2=2.41
r38 12 25 6.03242 $w=2.45e-07 $l=3e-07 $layer=LI1_cond $X=15.582 $Y=1.55
+ $X2=15.582 $Y2=1.85
r39 12 17 19.7562 $w=2.43e-07 $l=4.2e-07 $layer=LI1_cond $X=15.582 $Y=1.55
+ $X2=15.582 $Y2=1.13
r40 7 17 6.55101 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=15.54 $Y=0.965
+ $X2=15.54 $Y2=1.13
r41 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=15.54 $Y=0.965
+ $X2=15.54 $Y2=0.515
r42 2 23 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=15.425
+ $Y=1.84 $X2=15.58 $Y2=1.985
r43 2 15 300 $w=1.7e-07 $l=6.42845e-07 $layer=licon1_PDIFF $count=2 $X=15.425
+ $Y=1.84 $X2=15.58 $Y2=2.41
r44 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.4
+ $Y=0.37 $X2=15.54 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SEDFXTP_2%VGND 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49
+ 53 57 61 63 65 68 69 70 72 77 82 94 98 103 116 121 127 130 133 136 139 142 147
+ 150 152 156
c186 45 0 1.9935e-19 $X=6.405 $Y=0.515
c187 33 0 1.74672e-19 $X=1.22 $Y=0.58
r188 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=0
+ $X2=16.08 $Y2=0
r189 152 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r190 149 150 11.2171 $w=7.63e-07 $l=1.65e-07 $layer=LI1_cond $X=13.98 $Y=0.297
+ $X2=14.145 $Y2=0.297
r191 145 149 4.6905 $w=7.63e-07 $l=3e-07 $layer=LI1_cond $X=13.68 $Y=0.297
+ $X2=13.98 $Y2=0.297
r192 145 147 15.9858 $w=7.63e-07 $l=4.7e-07 $layer=LI1_cond $X=13.68 $Y=0.297
+ $X2=13.21 $Y2=0.297
r193 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r194 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r195 139 140 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r196 136 137 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r197 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r198 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r199 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r200 125 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=16.08 $Y2=0
r201 125 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=15.12 $Y2=0
r202 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r203 122 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.205 $Y=0
+ $X2=15.04 $Y2=0
r204 122 124 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=15.205 $Y=0
+ $X2=15.6 $Y2=0
r205 121 155 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=15.875 $Y=0
+ $X2=16.097 $Y2=0
r206 121 124 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=15.875 $Y=0
+ $X2=15.6 $Y2=0
r207 120 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.12 $Y2=0
r208 120 146 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=13.68 $Y2=0
r209 119 150 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=14.64 $Y=0
+ $X2=14.145 $Y2=0
r210 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r211 116 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.875 $Y=0
+ $X2=15.04 $Y2=0
r212 116 119 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=14.875 $Y=0
+ $X2=14.64 $Y2=0
r213 115 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r214 114 147 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=13.2 $Y=0
+ $X2=13.21 $Y2=0
r215 114 115 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r216 112 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r217 112 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r218 111 114 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r219 111 112 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r220 109 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.885 $Y=0
+ $X2=11.76 $Y2=0
r221 109 111 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=11.885 $Y=0
+ $X2=12.24 $Y2=0
r222 107 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r223 107 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.32 $Y2=0
r224 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r225 104 139 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=10.365 $Y=0
+ $X2=10.232 $Y2=0
r226 104 106 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=10.365 $Y=0
+ $X2=11.28 $Y2=0
r227 103 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.635 $Y=0
+ $X2=11.76 $Y2=0
r228 103 106 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=11.635 $Y=0
+ $X2=11.28 $Y2=0
r229 102 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r230 101 102 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r231 99 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.485 $Y=0
+ $X2=7.36 $Y2=0
r232 99 101 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=7.485 $Y=0
+ $X2=9.84 $Y2=0
r233 98 139 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=10.1 $Y=0
+ $X2=10.232 $Y2=0
r234 98 101 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=10.1 $Y=0 $X2=9.84
+ $Y2=0
r235 97 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r236 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r237 94 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.235 $Y=0
+ $X2=7.36 $Y2=0
r238 94 96 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.235 $Y=0
+ $X2=6.96 $Y2=0
r239 93 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r240 93 134 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r241 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r242 90 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.215 $Y=0
+ $X2=5.05 $Y2=0
r243 90 92 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=5.215 $Y=0 $X2=6
+ $Y2=0
r244 89 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r245 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r246 86 89 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r247 86 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r248 85 88 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r249 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r250 83 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.21 $Y2=0
r251 83 85 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.64 $Y2=0
r252 82 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.885 $Y=0
+ $X2=5.05 $Y2=0
r253 82 88 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.885 $Y=0
+ $X2=4.56 $Y2=0
r254 81 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r255 81 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r256 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r257 78 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0
+ $X2=1.22 $Y2=0
r258 78 80 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r259 77 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=2.21 $Y2=0
r260 77 80 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=1.68 $Y2=0
r261 75 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r262 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r263 72 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=1.22 $Y2=0
r264 72 74 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r265 70 102 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=8.16 $Y=0
+ $X2=9.84 $Y2=0
r266 70 137 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=8.16 $Y=0
+ $X2=7.44 $Y2=0
r267 68 92 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.235 $Y=0 $X2=6
+ $Y2=0
r268 68 69 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.235 $Y=0 $X2=6.365
+ $Y2=0
r269 67 96 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=6.495 $Y=0
+ $X2=6.96 $Y2=0
r270 67 69 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.495 $Y=0 $X2=6.365
+ $Y2=0
r271 63 155 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=16.04 $Y=0.085
+ $X2=16.097 $Y2=0
r272 63 65 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=16.04 $Y=0.085
+ $X2=16.04 $Y2=0.515
r273 59 152 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.04 $Y=0.085
+ $X2=15.04 $Y2=0
r274 59 61 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=15.04 $Y=0.085
+ $X2=15.04 $Y2=0.515
r275 55 142 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.76 $Y=0.085
+ $X2=11.76 $Y2=0
r276 55 57 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.76 $Y=0.085
+ $X2=11.76 $Y2=0.515
r277 51 139 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=10.232 $Y=0.085
+ $X2=10.232 $Y2=0
r278 51 53 18.7 $w=2.63e-07 $l=4.3e-07 $layer=LI1_cond $X=10.232 $Y=0.085
+ $X2=10.232 $Y2=0.515
r279 47 136 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0
r280 47 49 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0.515
r281 43 69 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.365 $Y=0.085
+ $X2=6.365 $Y2=0
r282 43 45 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=6.365 $Y=0.085
+ $X2=6.365 $Y2=0.515
r283 39 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.05 $Y=0.085
+ $X2=5.05 $Y2=0
r284 39 41 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=5.05 $Y=0.085
+ $X2=5.05 $Y2=0.805
r285 35 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0
r286 35 37 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0.775
r287 31 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r288 31 33 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.58
r289 10 65 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=15.83
+ $Y=0.37 $X2=16.04 $Y2=0.515
r290 9 61 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=14.895
+ $Y=0.37 $X2=15.04 $Y2=0.515
r291 8 149 91 $w=1.7e-07 $l=8.14279e-07 $layer=licon1_NDIFF $count=2 $X=13.235
+ $Y=0.37 $X2=13.98 $Y2=0.515
r292 7 57 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=11.575
+ $Y=0.37 $X2=11.72 $Y2=0.515
r293 6 53 182 $w=1.7e-07 $l=2.39531e-07 $layer=licon1_NDIFF $count=1 $X=10.045
+ $Y=0.485 $X2=10.27 $Y2=0.515
r294 5 49 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.255
+ $Y=0.37 $X2=7.4 $Y2=0.515
r295 4 45 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=6.255
+ $Y=0.37 $X2=6.405 $Y2=0.515
r296 3 41 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=4.84
+ $Y=0.625 $X2=5.05 $Y2=0.805
r297 2 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.565 $X2=2.21 $Y2=0.775
r298 1 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.37 $X2=1.22 $Y2=0.58
.ends

