* NGSPICE file created from sky130_fd_sc_ls__xor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__xor2_1 A B VGND VNB VPB VPWR X
M1000 VGND B a_194_125# VNB nshort w=550000u l=150000u
+  ad=8.846e+11p pd=6.8e+06u as=3.5475e+11p ps=2.39e+06u
M1001 a_455_87# A VGND VNB nshort w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1002 X B a_455_87# VNB nshort w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1003 a_194_125# B a_158_392# VPB phighvt w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=2.7e+11p ps=2.54e+06u
M1004 a_355_368# B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=7.672e+11p pd=5.85e+06u as=7.654e+11p ps=5.67e+06u
M1005 a_194_125# A VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_158_392# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_355_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_194_125# a_355_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.864e+11p pd=2.93e+06u as=0p ps=0u
M1009 VGND a_194_125# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

