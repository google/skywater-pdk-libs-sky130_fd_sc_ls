# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__decaphe_18
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__decaphe_18 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.640000 0.085000 ;
        RECT 0.085000  0.085000 8.555000 1.080000 ;
        RECT 0.085000  1.080000 1.155000 1.600000 ;
        RECT 2.205000  1.080000 2.895000 1.600000 ;
        RECT 3.965000  1.080000 4.655000 1.600000 ;
        RECT 5.725000  1.080000 6.415000 1.600000 ;
        RECT 7.485000  1.080000 8.555000 1.600000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.640000 3.415000 ;
        RECT 0.085000 1.770000 8.555000 3.245000 ;
        RECT 1.325000 1.250000 2.015000 1.770000 ;
        RECT 3.085000 1.250000 3.775000 1.770000 ;
        RECT 4.845000 1.250000 5.535000 1.770000 ;
        RECT 6.605000 1.250000 7.295000 1.770000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
END sky130_fd_sc_ls__decaphe_18
