* NGSPICE file created from sky130_fd_sc_ls__ebufn_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__ebufn_4 A TE_B VGND VNB VPB VPWR Z
M1000 a_208_74# TE_B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=1.036e+12p ps=8.57e+06u
M1001 a_348_368# TE_B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=1.6632e+12p pd=1.417e+07u as=0p ps=0u
M1002 Z a_27_368# a_348_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1003 VGND A a_27_368# VNB nshort w=740000u l=150000u
+  ad=6.216e+11p pd=6.12e+06u as=2.109e+11p ps=2.05e+06u
M1004 a_378_74# a_27_368# Z VNB nshort w=740000u l=150000u
+  ad=1.0323e+12p pd=1.019e+07u as=4.292e+11p ps=4.12e+06u
M1005 VGND a_208_74# a_378_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_378_74# a_208_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR TE_B a_348_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_348_368# a_27_368# Z VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR TE_B a_348_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_208_74# a_378_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_208_74# TE_B VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1012 a_348_368# TE_B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_378_74# a_27_368# Z VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Z a_27_368# a_378_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1016 a_378_74# a_208_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Z a_27_368# a_348_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Z a_27_368# a_378_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_348_368# a_27_368# Z VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

