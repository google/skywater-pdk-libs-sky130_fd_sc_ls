* File: sky130_fd_sc_ls__einvn_8.spice
* Created: Wed Sep  2 11:06:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__einvn_8.pex.spice"
.subckt sky130_fd_sc_ls__einvn_8  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1032 N_A_126_74#_M1032_d N_TE_B_M1032_g N_VGND_M1032_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A_126_74#_M1003_g N_A_293_74#_M1003_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75007 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1003_d N_A_126_74#_M1005_g N_A_293_74#_M1005_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75006.6 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_126_74#_M1015_g N_A_293_74#_M1005_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75006.1 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1015_d N_A_126_74#_M1016_g N_A_293_74#_M1016_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75005.6 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1019_d N_A_126_74#_M1019_g N_A_293_74#_M1016_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75005.2 A=0.111 P=1.78 MULT=1
MM1026 N_VGND_M1019_d N_A_126_74#_M1026_g N_A_293_74#_M1026_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75002.5 SB=75004.7 A=0.111 P=1.78 MULT=1
MM1030 N_VGND_M1030_d N_A_126_74#_M1030_g N_A_293_74#_M1026_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75004.3 A=0.111 P=1.78 MULT=1
MM1033 N_VGND_M1030_d N_A_126_74#_M1033_g N_A_293_74#_M1033_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.4 SB=75003.9 A=0.111 P=1.78 MULT=1
MM1004 N_Z_M1004_d N_A_M1004_g N_A_293_74#_M1033_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.8
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1007 N_Z_M1004_d N_A_M1007_g N_A_293_74#_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.2
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1010 N_Z_M1010_d N_A_M1010_g N_A_293_74#_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.6
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1013 N_Z_M1010_d N_A_M1013_g N_A_293_74#_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75005.1
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1017 N_Z_M1017_d N_A_M1017_g N_A_293_74#_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.6
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1022 N_Z_M1017_d N_A_M1022_g N_A_293_74#_M1022_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1024 N_Z_M1024_d N_A_M1024_g N_A_293_74#_M1022_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75006.4
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1029 N_Z_M1024_d N_A_M1029_g N_A_293_74#_M1029_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.2109 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75007
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_A_126_74#_M1020_d N_TE_B_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.3864 PD=2.83 PS=2.93 NRD=1.7533 NRS=10.5395 M=1
+ R=7.46667 SA=75000.3 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_VPWR_M1000_d N_TE_B_M1000_g N_A_239_368#_M1000_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.3304 PD=1.47 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75007.3 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1000_d N_TE_B_M1002_g N_A_239_368#_M1002_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75006.8 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1008_d N_TE_B_M1008_g N_A_239_368#_M1002_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75006.3 A=0.168 P=2.54 MULT=1
MM1012 N_VPWR_M1008_d N_TE_B_M1012_g N_A_239_368#_M1012_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75005.8 A=0.168 P=2.54 MULT=1
MM1018 N_VPWR_M1018_d N_TE_B_M1018_g N_A_239_368#_M1012_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75005.4 A=0.168 P=2.54 MULT=1
MM1023 N_VPWR_M1018_d N_TE_B_M1023_g N_A_239_368#_M1023_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.6 SB=75004.9 A=0.168 P=2.54 MULT=1
MM1027 N_VPWR_M1027_d N_TE_B_M1027_g N_A_239_368#_M1023_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.1 SB=75004.4 A=0.168 P=2.54 MULT=1
MM1031 N_VPWR_M1027_d N_TE_B_M1031_g N_A_239_368#_M1031_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.6 SB=75003.9 A=0.168 P=2.54 MULT=1
MM1001 N_Z_M1001_d N_A_M1001_g N_A_239_368#_M1031_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.1 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1006 N_Z_M1001_d N_A_M1006_g N_A_239_368#_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.5 SB=75003 A=0.168 P=2.54 MULT=1
MM1009 N_Z_M1009_d N_A_M1009_g N_A_239_368#_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75005 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1011 N_Z_M1009_d N_A_M1011_g N_A_239_368#_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.5 SB=75002 A=0.168 P=2.54 MULT=1
MM1014 N_Z_M1014_d N_A_M1014_g N_A_239_368#_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.9 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1021 N_Z_M1014_d N_A_M1021_g N_A_239_368#_M1021_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.4 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1025 N_Z_M1025_d N_A_M1025_g N_A_239_368#_M1021_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.8 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1028 N_Z_M1025_d N_A_M1028_g N_A_239_368#_M1028_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.3 SB=75000.2 A=0.168 P=2.54 MULT=1
DX34_noxref VNB VPB NWDIODE A=17.67 P=22.72
*
.include "sky130_fd_sc_ls__einvn_8.pxi.spice"
*
.ends
*
*
