* File: sky130_fd_sc_ls__a41o_4.pex.spice
* Created: Wed Sep  2 10:53:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A41O_4%B1 3 5 7 10 12 14 15 19 22
c46 10 0 1.35715e-19 $X=0.92 $Y=0.86
r47 22 23 11.2555 $w=3.64e-07 $l=8.5e-08 $layer=POLY_cond $X=0.92 $Y=1.667
+ $X2=1.005 $Y2=1.667
r48 21 22 54.9533 $w=3.64e-07 $l=4.15e-07 $layer=POLY_cond $X=0.505 $Y=1.667
+ $X2=0.92 $Y2=1.667
r49 20 21 1.98626 $w=3.64e-07 $l=1.5e-08 $layer=POLY_cond $X=0.49 $Y=1.667
+ $X2=0.505 $Y2=1.667
r50 18 20 13.9038 $w=3.64e-07 $l=1.05e-07 $layer=POLY_cond $X=0.385 $Y=1.667
+ $X2=0.49 $Y2=1.667
r51 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.615 $X2=0.385 $Y2=1.615
r52 15 19 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.385 $Y2=1.615
r53 12 23 23.572 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=1.005 $Y=1.885
+ $X2=1.005 $Y2=1.667
r54 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.005 $Y=1.885
+ $X2=1.005 $Y2=2.46
r55 8 22 23.572 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=0.92 $Y=1.45 $X2=0.92
+ $Y2=1.667
r56 8 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.92 $Y=1.45 $X2=0.92
+ $Y2=0.86
r57 5 21 23.572 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=1.667
r58 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.46
r59 1 20 23.572 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=0.49 $Y=1.45 $X2=0.49
+ $Y2=1.667
r60 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.49 $Y=1.45 $X2=0.49
+ $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_4%A_113_98# 1 2 3 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 38 40 47 51 52 53 58 59 72
c146 52 0 6.95417e-20 $X=4.165 $Y=0.34
c147 31 0 1.26721e-19 $X=3.365 $Y=1.765
r148 72 73 57.2541 $w=3.62e-07 $l=4.3e-07 $layer=POLY_cond $X=2.935 $Y=1.552
+ $X2=3.365 $Y2=1.552
r149 71 72 2.66298 $w=3.62e-07 $l=2e-08 $layer=POLY_cond $X=2.915 $Y=1.552
+ $X2=2.935 $Y2=1.552
r150 70 71 54.5912 $w=3.62e-07 $l=4.1e-07 $layer=POLY_cond $X=2.505 $Y=1.552
+ $X2=2.915 $Y2=1.552
r151 69 70 5.32597 $w=3.62e-07 $l=4e-08 $layer=POLY_cond $X=2.465 $Y=1.552
+ $X2=2.505 $Y2=1.552
r152 66 67 11.3177 $w=3.62e-07 $l=8.5e-08 $layer=POLY_cond $X=1.93 $Y=1.552
+ $X2=2.015 $Y2=1.552
r153 59 62 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=4.33 $Y=0.34
+ $X2=4.33 $Y2=0.515
r154 56 57 16.4106 $w=5.65e-07 $l=7.6e-07 $layer=LI1_cond $X=0.882 $Y=0.745
+ $X2=0.882 $Y2=1.505
r155 55 56 2.37522 $w=5.65e-07 $l=2.25386e-07 $layer=LI1_cond $X=0.705 $Y=0.635
+ $X2=0.882 $Y2=0.745
r156 52 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.165 $Y=0.34
+ $X2=4.33 $Y2=0.34
r157 52 53 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.165 $Y=0.34
+ $X2=3.645 $Y2=0.34
r158 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.56 $Y=0.425
+ $X2=3.645 $Y2=0.34
r159 50 51 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.56 $Y=0.425
+ $X2=3.56 $Y2=0.66
r160 48 69 32.6215 $w=3.62e-07 $l=2.45e-07 $layer=POLY_cond $X=2.22 $Y=1.552
+ $X2=2.465 $Y2=1.552
r161 48 67 27.2956 $w=3.62e-07 $l=2.05e-07 $layer=POLY_cond $X=2.22 $Y=1.552
+ $X2=2.015 $Y2=1.552
r162 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.22
+ $Y=1.505 $X2=2.22 $Y2=1.505
r163 45 66 51.9282 $w=3.62e-07 $l=3.9e-07 $layer=POLY_cond $X=1.54 $Y=1.552
+ $X2=1.93 $Y2=1.552
r164 45 64 5.32597 $w=3.62e-07 $l=4e-08 $layer=POLY_cond $X=1.54 $Y=1.552
+ $X2=1.5 $Y2=1.552
r165 44 47 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.54 $Y=1.505
+ $X2=2.22 $Y2=1.505
r166 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.54
+ $Y=1.505 $X2=1.54 $Y2=1.505
r167 42 57 3.88339 $w=3.3e-07 $l=3.43e-07 $layer=LI1_cond $X=1.225 $Y=1.505
+ $X2=0.882 $Y2=1.505
r168 42 44 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.225 $Y=1.505
+ $X2=1.54 $Y2=1.505
r169 41 56 7.93092 $w=1.7e-07 $l=3.43e-07 $layer=LI1_cond $X=1.225 $Y=0.745
+ $X2=0.882 $Y2=0.745
r170 40 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.475 $Y=0.745
+ $X2=3.56 $Y2=0.66
r171 40 41 146.791 $w=1.68e-07 $l=2.25e-06 $layer=LI1_cond $X=3.475 $Y=0.745
+ $X2=1.225 $Y2=0.745
r172 38 57 10.1272 $w=5.65e-07 $l=1.99825e-07 $layer=LI1_cond $X=0.805 $Y=1.67
+ $X2=0.882 $Y2=1.505
r173 38 58 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.805 $Y=1.67
+ $X2=0.805 $Y2=1.95
r174 34 58 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=0.752 $Y=2.087
+ $X2=0.752 $Y2=1.95
r175 34 36 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=0.752 $Y=2.087
+ $X2=0.752 $Y2=2.115
r176 31 73 23.4391 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=3.365 $Y=1.765
+ $X2=3.365 $Y2=1.552
r177 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.365 $Y=1.765
+ $X2=3.365 $Y2=2.4
r178 28 72 23.4391 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=2.935 $Y=1.34
+ $X2=2.935 $Y2=1.552
r179 28 30 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.935 $Y=1.34
+ $X2=2.935 $Y2=0.86
r180 25 71 23.4391 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=2.915 $Y=1.765
+ $X2=2.915 $Y2=1.552
r181 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.915 $Y=1.765
+ $X2=2.915 $Y2=2.4
r182 22 70 23.4391 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=2.505 $Y=1.34
+ $X2=2.505 $Y2=1.552
r183 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.505 $Y=1.34
+ $X2=2.505 $Y2=0.86
r184 19 69 23.4391 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=2.465 $Y=1.765
+ $X2=2.465 $Y2=1.552
r185 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.465 $Y=1.765
+ $X2=2.465 $Y2=2.4
r186 16 67 23.4391 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=2.015 $Y=1.765
+ $X2=2.015 $Y2=1.552
r187 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.015 $Y=1.765
+ $X2=2.015 $Y2=2.4
r188 13 66 23.4391 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=1.93 $Y=1.34
+ $X2=1.93 $Y2=1.552
r189 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.93 $Y=1.34
+ $X2=1.93 $Y2=0.86
r190 10 64 23.4391 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=1.5 $Y=1.34
+ $X2=1.5 $Y2=1.552
r191 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.5 $Y=1.34 $X2=1.5
+ $Y2=0.86
r192 3 36 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.96 $X2=0.78 $Y2=2.115
r193 2 62 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.19
+ $Y=0.37 $X2=4.33 $Y2=0.515
r194 1 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.49 $X2=0.705 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_4%A1 1 3 6 8 10 13 15 16 24
c57 16 0 1.26721e-19 $X=4.08 $Y=1.665
c58 13 0 1.79117e-19 $X=4.545 $Y=0.74
r59 24 25 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=4.53 $Y=1.667
+ $X2=4.545 $Y2=1.667
r60 23 24 53.3413 $w=3.75e-07 $l=4.15e-07 $layer=POLY_cond $X=4.115 $Y=1.667
+ $X2=4.53 $Y2=1.667
r61 21 23 10.9253 $w=3.75e-07 $l=8.5e-08 $layer=POLY_cond $X=4.03 $Y=1.667
+ $X2=4.115 $Y2=1.667
r62 19 21 18.6373 $w=3.75e-07 $l=1.45e-07 $layer=POLY_cond $X=3.885 $Y=1.667
+ $X2=4.03 $Y2=1.667
r63 16 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.03
+ $Y=1.615 $X2=4.03 $Y2=1.615
r64 15 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.6 $Y=1.615
+ $X2=4.03 $Y2=1.615
r65 11 25 24.2915 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=4.545 $Y=1.45
+ $X2=4.545 $Y2=1.667
r66 11 13 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.545 $Y=1.45
+ $X2=4.545 $Y2=0.74
r67 8 24 24.2915 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=4.53 $Y=1.885
+ $X2=4.53 $Y2=1.667
r68 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.53 $Y=1.885
+ $X2=4.53 $Y2=2.46
r69 4 23 24.2915 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=4.115 $Y=1.45
+ $X2=4.115 $Y2=1.667
r70 4 6 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.115 $Y=1.45
+ $X2=4.115 $Y2=0.74
r71 1 19 24.2915 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=3.885 $Y=1.885
+ $X2=3.885 $Y2=1.667
r72 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.885 $Y=1.885
+ $X2=3.885 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_4%A2 3 5 7 10 12 14 15 16 24
r54 24 25 37.8931 $w=3.18e-07 $l=2.5e-07 $layer=POLY_cond $X=5.405 $Y=1.667
+ $X2=5.655 $Y2=1.667
r55 23 24 30.3145 $w=3.18e-07 $l=2e-07 $layer=POLY_cond $X=5.205 $Y=1.667
+ $X2=5.405 $Y2=1.667
r56 21 23 21.2201 $w=3.18e-07 $l=1.4e-07 $layer=POLY_cond $X=5.065 $Y=1.667
+ $X2=5.205 $Y2=1.667
r57 19 21 13.6415 $w=3.18e-07 $l=9e-08 $layer=POLY_cond $X=4.975 $Y=1.667
+ $X2=5.065 $Y2=1.667
r58 15 16 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.615
+ $X2=5.52 $Y2=1.615
r59 15 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.065
+ $Y=1.615 $X2=5.065 $Y2=1.615
r60 12 25 20.3436 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=5.655 $Y=1.885
+ $X2=5.655 $Y2=1.667
r61 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.655 $Y=1.885
+ $X2=5.655 $Y2=2.46
r62 8 24 20.3436 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=5.405 $Y=1.45
+ $X2=5.405 $Y2=1.667
r63 8 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.405 $Y=1.45
+ $X2=5.405 $Y2=0.74
r64 5 23 20.3436 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=5.205 $Y=1.885
+ $X2=5.205 $Y2=1.667
r65 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.205 $Y=1.885
+ $X2=5.205 $Y2=2.46
r66 1 19 20.3436 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=4.975 $Y=1.45
+ $X2=4.975 $Y2=1.667
r67 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.975 $Y=1.45
+ $X2=4.975 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_4%A3 1 3 6 8 10 13 15 16 17 26
c58 6 0 1.25271e-19 $X=6.38 $Y=0.74
r59 26 27 13.3536 $w=3.79e-07 $l=1.05e-07 $layer=POLY_cond $X=6.705 $Y=1.667
+ $X2=6.81 $Y2=1.667
r60 24 26 10.81 $w=3.79e-07 $l=8.5e-08 $layer=POLY_cond $X=6.62 $Y=1.667
+ $X2=6.705 $Y2=1.667
r61 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.62
+ $Y=1.615 $X2=6.62 $Y2=1.615
r62 22 24 30.5224 $w=3.79e-07 $l=2.4e-07 $layer=POLY_cond $X=6.38 $Y=1.667
+ $X2=6.62 $Y2=1.667
r63 21 22 22.2559 $w=3.79e-07 $l=1.75e-07 $layer=POLY_cond $X=6.205 $Y=1.667
+ $X2=6.38 $Y2=1.667
r64 17 25 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.96 $Y=1.615
+ $X2=6.62 $Y2=1.615
r65 16 25 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=6.48 $Y=1.615
+ $X2=6.62 $Y2=1.615
r66 15 16 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6 $Y=1.615 $X2=6.48
+ $Y2=1.615
r67 11 27 24.5487 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=6.81 $Y=1.45
+ $X2=6.81 $Y2=1.667
r68 11 13 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.81 $Y=1.45
+ $X2=6.81 $Y2=0.74
r69 8 26 24.5487 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=6.705 $Y=1.885
+ $X2=6.705 $Y2=1.667
r70 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.705 $Y=1.885
+ $X2=6.705 $Y2=2.46
r71 4 22 24.5487 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=6.38 $Y=1.45
+ $X2=6.38 $Y2=1.667
r72 4 6 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.38 $Y=1.45 $X2=6.38
+ $Y2=0.74
r73 1 21 24.5487 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=6.205 $Y=1.885
+ $X2=6.205 $Y2=1.667
r74 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.205 $Y=1.885
+ $X2=6.205 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_4%A4 1 3 6 8 10 13 15 16 24
r41 24 25 1.85385 $w=3.9e-07 $l=1.5e-08 $layer=POLY_cond $X=7.655 $Y=1.667
+ $X2=7.67 $Y2=1.667
r42 22 24 20.3923 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=7.49 $Y=1.667
+ $X2=7.655 $Y2=1.667
r43 20 22 30.8974 $w=3.9e-07 $l=2.5e-07 $layer=POLY_cond $X=7.24 $Y=1.667
+ $X2=7.49 $Y2=1.667
r44 19 20 4.32564 $w=3.9e-07 $l=3.5e-08 $layer=POLY_cond $X=7.205 $Y=1.667
+ $X2=7.24 $Y2=1.667
r45 15 16 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.615
+ $X2=7.92 $Y2=1.615
r46 15 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.49
+ $Y=1.615 $X2=7.49 $Y2=1.615
r47 11 25 25.2441 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=7.67 $Y=1.45
+ $X2=7.67 $Y2=1.667
r48 11 13 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=7.67 $Y=1.45
+ $X2=7.67 $Y2=0.74
r49 8 24 25.2441 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=7.655 $Y=1.885
+ $X2=7.655 $Y2=1.667
r50 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.655 $Y=1.885
+ $X2=7.655 $Y2=2.46
r51 4 20 25.2441 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=7.24 $Y=1.45
+ $X2=7.24 $Y2=1.667
r52 4 6 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=7.24 $Y=1.45 $X2=7.24
+ $Y2=0.74
r53 1 19 25.2441 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=7.205 $Y=1.885
+ $X2=7.205 $Y2=1.667
r54 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.205 $Y=1.885
+ $X2=7.205 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_4%A_27_392# 1 2 3 4 5 6 21 25 26 29 34 35 37 38
+ 41 45 47 51 53 55 57 59 63 65 67
c135 59 0 1.25754e-19 $X=1.23 $Y=2.375
r136 55 69 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.43 $Y=2.12 $X2=7.43
+ $Y2=2.035
r137 55 57 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=7.43 $Y=2.12
+ $X2=7.43 $Y2=2.815
r138 54 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.595 $Y=2.035
+ $X2=6.43 $Y2=2.035
r139 53 69 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.265 $Y=2.035
+ $X2=7.43 $Y2=2.035
r140 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.265 $Y=2.035
+ $X2=6.595 $Y2=2.035
r141 49 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.43 $Y=2.12
+ $X2=6.43 $Y2=2.035
r142 49 51 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.43 $Y=2.12
+ $X2=6.43 $Y2=2.815
r143 48 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.595 $Y=2.035
+ $X2=5.43 $Y2=2.035
r144 47 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.265 $Y=2.035
+ $X2=6.43 $Y2=2.035
r145 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.265 $Y=2.035
+ $X2=5.595 $Y2=2.035
r146 43 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.43 $Y=2.12
+ $X2=5.43 $Y2=2.035
r147 43 45 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.43 $Y=2.12
+ $X2=5.43 $Y2=2.815
r148 42 61 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.375 $Y=2.035
+ $X2=4.21 $Y2=2.035
r149 41 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.265 $Y=2.035
+ $X2=5.43 $Y2=2.035
r150 41 42 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=5.265 $Y=2.035
+ $X2=4.375 $Y2=2.035
r151 38 63 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.21 $Y=2.29
+ $X2=4.21 $Y2=2.375
r152 37 61 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.21 $Y=2.12 $X2=4.21
+ $Y2=2.035
r153 37 38 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.21 $Y=2.12
+ $X2=4.21 $Y2=2.29
r154 36 59 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=2.375
+ $X2=1.23 $Y2=2.375
r155 35 63 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.045 $Y=2.375
+ $X2=4.21 $Y2=2.375
r156 35 36 172.888 $w=1.68e-07 $l=2.65e-06 $layer=LI1_cond $X=4.045 $Y=2.375
+ $X2=1.395 $Y2=2.375
r157 32 34 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.23 $Y2=2.815
r158 31 59 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.46
+ $X2=1.23 $Y2=2.375
r159 31 34 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.23 $Y=2.46
+ $X2=1.23 $Y2=2.815
r160 27 59 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.29
+ $X2=1.23 $Y2=2.375
r161 27 29 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.23 $Y=2.29
+ $X2=1.23 $Y2=2.105
r162 25 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.065 $Y=2.99
+ $X2=1.23 $Y2=2.905
r163 25 26 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.065 $Y=2.99
+ $X2=0.445 $Y2=2.99
r164 21 24 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115
+ $X2=0.28 $Y2=2.815
r165 19 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r166 19 24 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.28 $Y2=2.815
r167 6 69 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=7.28
+ $Y=1.96 $X2=7.43 $Y2=2.115
r168 6 57 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=7.28
+ $Y=1.96 $X2=7.43 $Y2=2.815
r169 5 67 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.96 $X2=6.43 $Y2=2.115
r170 5 51 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.96 $X2=6.43 $Y2=2.815
r171 4 65 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.96 $X2=5.43 $Y2=2.115
r172 4 45 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.96 $X2=5.43 $Y2=2.815
r173 3 63 300 $w=1.7e-07 $l=6.07268e-07 $layer=licon1_PDIFF $count=2 $X=3.96
+ $Y=1.96 $X2=4.21 $Y2=2.455
r174 3 61 600 $w=1.7e-07 $l=3.18198e-07 $layer=licon1_PDIFF $count=1 $X=3.96
+ $Y=1.96 $X2=4.21 $Y2=2.115
r175 2 34 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.96 $X2=1.23 $Y2=2.815
r176 2 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.96 $X2=1.23 $Y2=2.105
r177 1 24 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r178 1 21 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_4%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 46 48 53
+ 54 55 57 62 67 76 80 85 91 94 97 100 103 107
r107 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r108 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r109 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r110 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r111 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r113 89 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r114 89 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r115 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r116 86 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.095 $Y=3.33
+ $X2=6.93 $Y2=3.33
r117 86 88 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.095 $Y=3.33
+ $X2=7.44 $Y2=3.33
r118 85 106 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.977 $Y2=3.33
r119 85 88 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.44 $Y2=3.33
r120 84 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r121 84 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r122 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r123 81 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.095 $Y=3.33
+ $X2=5.93 $Y2=3.33
r124 81 83 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.095 $Y=3.33
+ $X2=6.48 $Y2=3.33
r125 80 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.765 $Y=3.33
+ $X2=6.93 $Y2=3.33
r126 80 83 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.765 $Y=3.33
+ $X2=6.48 $Y2=3.33
r127 79 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r128 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r129 76 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=5.93 $Y2=3.33
r130 76 78 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=5.52 $Y2=3.33
r131 75 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r132 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r133 72 97 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.775 $Y=3.33
+ $X2=3.6 $Y2=3.33
r134 72 74 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=3.775 $Y=3.33
+ $X2=4.56 $Y2=3.33
r135 71 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r136 71 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r137 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r138 68 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.69 $Y2=3.33
r139 68 70 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.12 $Y2=3.33
r140 67 97 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.6 $Y2=3.33
r141 67 70 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.12 $Y2=3.33
r142 66 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r143 66 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r144 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r145 63 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=1.79 $Y2=3.33
r146 63 65 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=2.16 $Y2=3.33
r147 62 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=2.69 $Y2=3.33
r148 62 65 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=2.16 $Y2=3.33
r149 60 92 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r150 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r151 57 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.625 $Y=3.33
+ $X2=1.79 $Y2=3.33
r152 57 59 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=1.625 $Y=3.33
+ $X2=0.24 $Y2=3.33
r153 55 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r154 55 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r155 53 74 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.635 $Y=3.33
+ $X2=4.56 $Y2=3.33
r156 53 54 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=4.635 $Y=3.33
+ $X2=4.865 $Y2=3.33
r157 52 78 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.095 $Y=3.33
+ $X2=5.52 $Y2=3.33
r158 52 54 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.095 $Y=3.33
+ $X2=4.865 $Y2=3.33
r159 48 51 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=7.92 $Y=2.115
+ $X2=7.92 $Y2=2.815
r160 46 106 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.977 $Y2=3.33
r161 46 51 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=2.815
r162 42 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.93 $Y=3.245
+ $X2=6.93 $Y2=3.33
r163 42 44 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.93 $Y=3.245
+ $X2=6.93 $Y2=2.415
r164 38 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.93 $Y=3.245
+ $X2=5.93 $Y2=3.33
r165 38 40 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.93 $Y=3.245
+ $X2=5.93 $Y2=2.415
r166 34 54 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.865 $Y=3.245
+ $X2=4.865 $Y2=3.33
r167 34 36 22.6215 $w=4.58e-07 $l=8.7e-07 $layer=LI1_cond $X=4.865 $Y=3.245
+ $X2=4.865 $Y2=2.375
r168 30 97 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=3.245 $X2=3.6
+ $Y2=3.33
r169 30 32 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=3.245
+ $X2=3.6 $Y2=2.765
r170 26 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.69 $Y=3.245
+ $X2=2.69 $Y2=3.33
r171 26 28 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.69 $Y=3.245
+ $X2=2.69 $Y2=2.755
r172 22 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=3.245
+ $X2=1.79 $Y2=3.33
r173 22 24 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.79 $Y=3.245
+ $X2=1.79 $Y2=2.755
r174 7 51 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.96 $X2=7.88 $Y2=2.815
r175 7 48 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.96 $X2=7.88 $Y2=2.115
r176 6 44 300 $w=1.7e-07 $l=5.24667e-07 $layer=licon1_PDIFF $count=2 $X=6.78
+ $Y=1.96 $X2=6.93 $Y2=2.415
r177 5 40 300 $w=1.7e-07 $l=5.45917e-07 $layer=licon1_PDIFF $count=2 $X=5.73
+ $Y=1.96 $X2=5.93 $Y2=2.415
r178 4 36 300 $w=1.7e-07 $l=5.29268e-07 $layer=licon1_PDIFF $count=2 $X=4.605
+ $Y=1.96 $X2=4.865 $Y2=2.375
r179 3 32 600 $w=1.7e-07 $l=1.00181e-06 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.84 $X2=3.6 $Y2=2.765
r180 2 28 600 $w=1.7e-07 $l=9.87155e-07 $layer=licon1_PDIFF $count=1 $X=2.54
+ $Y=1.84 $X2=2.69 $Y2=2.755
r181 1 24 600 $w=1.7e-07 $l=9.84835e-07 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=1.84 $X2=1.79 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_4%X 1 2 3 4 13 17 21 24 25 26 30
c41 13 0 1.35715e-19 $X=2.555 $Y=1.085
r42 26 30 2.40606 $w=7.5e-07 $l=1.4e-07 $layer=LI1_cond $X=2.93 $Y=1.98 $X2=2.93
+ $Y2=1.84
r43 25 30 2.79085 $w=7.48e-07 $l=1.75e-07 $layer=LI1_cond $X=2.93 $Y=1.665
+ $X2=2.93 $Y2=1.84
r44 24 25 5.90065 $w=7.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.93 $Y=1.295
+ $X2=2.93 $Y2=1.665
r45 21 24 1.99346 $w=7.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.93 $Y=1.17
+ $X2=2.93 $Y2=1.295
r46 21 23 2.06231 $w=7.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=1.17 $X2=2.93
+ $Y2=1.085
r47 17 26 6.44481 $w=2.8e-07 $l=3.75e-07 $layer=LI1_cond $X=2.555 $Y=1.98
+ $X2=2.93 $Y2=1.98
r48 17 19 12.965 $w=2.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.555 $Y=1.98
+ $X2=2.24 $Y2=1.98
r49 13 23 9.09843 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=2.555 $Y=1.085
+ $X2=2.93 $Y2=1.085
r50 13 15 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.555 $Y=1.085
+ $X2=1.715 $Y2=1.085
r51 4 26 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.84 $X2=3.14 $Y2=2.01
r52 3 19 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=2.09
+ $Y=1.84 $X2=2.24 $Y2=2.02
r53 2 23 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.58
+ $Y=0.49 $X2=2.72 $Y2=1.085
r54 1 15 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.575
+ $Y=0.49 $X2=1.715 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_4%VGND 1 2 3 4 5 16 18 22 26 28 32 36 38 40 45
+ 50 60 61 67 70 73 76
r97 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r98 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r99 71 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r100 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r101 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r102 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r103 61 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r104 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r105 58 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.62 $Y=0 $X2=7.455
+ $Y2=0
r106 58 60 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.62 $Y=0 $X2=7.92
+ $Y2=0
r107 57 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r108 56 57 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r109 54 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r110 53 56 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=6.96
+ $Y2=0
r111 53 54 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r112 51 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.18
+ $Y2=0
r113 51 53 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.6
+ $Y2=0
r114 50 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.29 $Y=0 $X2=7.455
+ $Y2=0
r115 50 56 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.29 $Y=0 $X2=6.96
+ $Y2=0
r116 49 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r117 49 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r118 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r119 46 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.21
+ $Y2=0
r120 46 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0
+ $X2=1.68 $Y2=0
r121 45 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.055 $Y=0 $X2=2.22
+ $Y2=0
r122 45 48 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.055 $Y=0
+ $X2=1.68 $Y2=0
r123 44 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r124 44 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r125 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r126 41 64 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.18
+ $Y2=0
r127 41 43 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.72
+ $Y2=0
r128 40 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.21
+ $Y2=0
r129 40 43 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0
+ $X2=0.72 $Y2=0
r130 38 57 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=6.96 $Y2=0
r131 38 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r132 34 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.455 $Y=0.085
+ $X2=7.455 $Y2=0
r133 34 36 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=7.455 $Y=0.085
+ $X2=7.455 $Y2=0.495
r134 30 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.18 $Y=0.085
+ $X2=3.18 $Y2=0
r135 30 32 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=3.18 $Y=0.085
+ $X2=3.18 $Y2=0.325
r136 29 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.385 $Y=0 $X2=2.22
+ $Y2=0
r137 28 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.055 $Y=0 $X2=3.18
+ $Y2=0
r138 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.055 $Y=0
+ $X2=2.385 $Y2=0
r139 24 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=0.085
+ $X2=2.22 $Y2=0
r140 24 26 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=2.22 $Y=0.085
+ $X2=2.22 $Y2=0.375
r141 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r142 20 22 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.375
r143 16 64 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.235 $Y=0.085
+ $X2=0.18 $Y2=0
r144 16 18 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=0.235 $Y=0.085
+ $X2=0.235 $Y2=0.635
r145 5 36 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=7.315
+ $Y=0.37 $X2=7.455 $Y2=0.495
r146 4 32 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=3.01
+ $Y=0.49 $X2=3.22 $Y2=0.325
r147 3 26 182 $w=1.7e-07 $l=2.66364e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.49 $X2=2.22 $Y2=0.375
r148 2 22 182 $w=1.7e-07 $l=2.66364e-07 $layer=licon1_NDIFF $count=1 $X=0.995
+ $Y=0.49 $X2=1.21 $Y2=0.375
r149 1 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.49 $X2=0.275 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_4%A_751_74# 1 2 3 10 12 13 14 21 27
r40 19 21 2.5834 $w=4.48e-07 $l=8.5e-08 $layer=LI1_cond $X=3.9 $Y=0.925
+ $X2=3.985 $Y2=0.925
r41 15 23 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.845 $Y=0.465
+ $X2=4.76 $Y2=0.465
r42 14 27 3.79804 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.455 $Y=0.465
+ $X2=5.62 $Y2=0.465
r43 14 15 26.0367 $w=2.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.455 $Y=0.465
+ $X2=4.845 $Y2=0.465
r44 13 25 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.76 $Y=0.77 $X2=4.76
+ $Y2=0.96
r45 12 23 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.76 $Y=0.6 $X2=4.76
+ $Y2=0.465
r46 12 13 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.76 $Y=0.6 $X2=4.76
+ $Y2=0.77
r47 10 25 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.675 $Y=0.96
+ $X2=4.76 $Y2=0.96
r48 10 21 20.9259 $w=3.78e-07 $l=6.9e-07 $layer=LI1_cond $X=4.675 $Y=0.96
+ $X2=3.985 $Y2=0.96
r49 3 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.48
+ $Y=0.37 $X2=5.62 $Y2=0.515
r50 2 25 182 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_NDIFF $count=1 $X=4.62
+ $Y=0.37 $X2=4.76 $Y2=0.985
r51 2 23 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.62
+ $Y=0.37 $X2=4.76 $Y2=0.495
r52 1 19 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=3.755
+ $Y=0.37 $X2=3.9 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_4%A_1010_74# 1 2 9 11 12 15
c24 9 0 1.09575e-19 $X=5.19 $Y=0.935
r25 13 15 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.595 $Y=1.11
+ $X2=6.595 $Y2=0.785
r26 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.51 $Y=1.195
+ $X2=6.595 $Y2=1.11
r27 11 12 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=6.51 $Y=1.195
+ $X2=5.285 $Y2=1.195
r28 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.155 $Y=1.11
+ $X2=5.285 $Y2=1.195
r29 7 9 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=5.155 $Y=1.11
+ $X2=5.155 $Y2=0.935
r30 2 15 182 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_NDIFF $count=1 $X=6.455
+ $Y=0.37 $X2=6.595 $Y2=0.785
r31 1 9 182 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_NDIFF $count=1 $X=5.05
+ $Y=0.37 $X2=5.19 $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_LS__A41O_4%A_1205_74# 1 2 3 12 14 15 19 20 21 24
c41 21 0 1.25271e-19 $X=7.11 $Y=1.195
r42 22 24 26.3732 $w=2.58e-07 $l=5.95e-07 $layer=LI1_cond $X=7.92 $Y=1.11
+ $X2=7.92 $Y2=0.515
r43 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.79 $Y=1.195
+ $X2=7.92 $Y2=1.11
r44 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.79 $Y=1.195
+ $X2=7.11 $Y2=1.195
r45 17 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.985 $Y=1.11
+ $X2=7.11 $Y2=1.195
r46 17 19 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=6.985 $Y=1.11
+ $X2=6.985 $Y2=0.515
r47 16 19 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=6.985 $Y=0.425
+ $X2=6.985 $Y2=0.515
r48 14 16 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.86 $Y=0.34
+ $X2=6.985 $Y2=0.425
r49 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.86 $Y=0.34
+ $X2=6.33 $Y2=0.34
r50 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.165 $Y=0.425
+ $X2=6.33 $Y2=0.34
r51 10 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.165 $Y=0.425
+ $X2=6.165 $Y2=0.515
r52 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.745
+ $Y=0.37 $X2=7.885 $Y2=0.515
r53 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.885
+ $Y=0.37 $X2=7.025 $Y2=0.515
r54 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.025
+ $Y=0.37 $X2=6.165 $Y2=0.515
.ends

