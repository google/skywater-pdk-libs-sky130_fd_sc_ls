* File: sky130_fd_sc_ls__o41a_1.pex.spice
* Created: Wed Sep  2 11:23:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O41A_1%A_83_270# 1 2 9 11 13 15 17 19 21 22 25 29
c64 21 0 1.75295e-19 $X=1.75 $Y=2.035
c65 17 0 6.43674e-20 $X=0.62 $Y=1.515
r66 27 29 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=1.915 $Y=2.12
+ $X2=1.915 $Y2=2.13
r67 23 25 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=1.34 $Y=1.11
+ $X2=1.34 $Y2=0.515
r68 21 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.75 $Y=2.035
+ $X2=1.915 $Y2=2.12
r69 21 22 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=1.75 $Y=2.035
+ $X2=0.785 $Y2=2.035
r70 20 31 2.6346 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.785 $Y=1.195
+ $X2=0.62 $Y2=1.195
r71 19 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.175 $Y=1.195
+ $X2=1.34 $Y2=1.11
r72 19 20 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.175 $Y=1.195
+ $X2=0.785 $Y2=1.195
r73 17 31 12.8588 $w=3.3e-07 $l=3.2e-07 $layer=LI1_cond $X=0.62 $Y=1.515
+ $X2=0.62 $Y2=1.195
r74 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.62
+ $Y=1.515 $X2=0.62 $Y2=1.515
r75 15 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.62 $Y=1.95
+ $X2=0.785 $Y2=2.035
r76 15 17 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=0.62 $Y=1.95
+ $X2=0.62 $Y2=1.515
r77 11 18 50.9845 $w=3.31e-07 $l=2.93684e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.6 $Y2=1.515
r78 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r79 7 18 38.6069 $w=3.31e-07 $l=2.11069e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.6 $Y2=1.515
r80 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
r81 2 29 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=1.68
+ $Y=1.985 $X2=1.915 $Y2=2.13
r82 1 25 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.195
+ $Y=0.37 $X2=1.34 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O41A_1%B1 3 5 7 8 12
c36 12 0 1.14234e-20 $X=1.415 $Y=1.615
c37 5 0 6.43674e-20 $X=1.605 $Y=1.91
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.415
+ $Y=1.615 $X2=1.415 $Y2=1.615
r39 8 12 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.415 $Y2=1.615
r40 5 11 55.2309 $w=4.01e-07 $l=3.55331e-07 $layer=POLY_cond $X=1.605 $Y=1.91
+ $X2=1.472 $Y2=1.615
r41 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.605 $Y=1.91
+ $X2=1.605 $Y2=2.405
r42 1 11 39.605 $w=4.01e-07 $l=2.02287e-07 $layer=POLY_cond $X=1.555 $Y=1.45
+ $X2=1.472 $Y2=1.615
r43 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.555 $Y=1.45
+ $X2=1.555 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__O41A_1%A4 3 5 6 7 9 10 14
c47 7 0 1.14234e-20 $X=2.14 $Y=1.765
r48 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.035
+ $Y=1.355 $X2=2.035 $Y2=1.355
r49 10 14 8.82117 $w=4.03e-07 $l=3.1e-07 $layer=LI1_cond $X=2.072 $Y=1.665
+ $X2=2.072 $Y2=1.355
r50 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.14 $Y=1.765
+ $X2=2.14 $Y2=2.4
r51 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.14 $Y=1.675 $X2=2.14
+ $Y2=1.765
r52 5 13 34.0194 $w=3.43e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.14 $Y=1.52
+ $X2=2.05 $Y2=1.355
r53 5 6 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=2.14 $Y=1.52 $X2=2.14
+ $Y2=1.675
r54 1 13 38.7084 $w=3.43e-07 $l=1.67481e-07 $layer=POLY_cond $X=2.055 $Y=1.19
+ $X2=2.05 $Y2=1.355
r55 1 3 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.055 $Y=1.19 $X2=2.055
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__O41A_1%A3 1 3 6 8 9 10 11 18
c39 1 0 1.75295e-19 $X=2.56 $Y=1.765
r40 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.635
+ $Y=1.385 $X2=2.635 $Y2=1.385
r41 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.635 $Y=2.405
+ $X2=2.635 $Y2=2.775
r42 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.635 $Y=2.035
+ $X2=2.635 $Y2=2.405
r43 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.635 $Y=1.665
+ $X2=2.635 $Y2=2.035
r44 8 18 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.635 $Y=1.665
+ $X2=2.635 $Y2=1.385
r45 4 17 38.9026 $w=2.7e-07 $l=1.69926e-07 $layer=POLY_cond $X=2.625 $Y=1.22
+ $X2=2.635 $Y2=1.385
r46 4 6 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.625 $Y=1.22
+ $X2=2.625 $Y2=0.69
r47 1 17 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=2.56 $Y=1.765
+ $X2=2.635 $Y2=1.385
r48 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.56 $Y=1.765
+ $X2=2.56 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O41A_1%A2 3 5 7 8 9 10 11 18
r34 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.205
+ $Y=1.465 $X2=3.205 $Y2=1.465
r35 10 11 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.187 $Y=2.405
+ $X2=3.187 $Y2=2.775
r36 9 10 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.187 $Y=2.035
+ $X2=3.187 $Y2=2.405
r37 8 9 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.187 $Y=1.665
+ $X2=3.187 $Y2=2.035
r38 8 18 6.31476 $w=3.63e-07 $l=2e-07 $layer=LI1_cond $X=3.187 $Y=1.665
+ $X2=3.187 $Y2=1.465
r39 5 17 61.4066 $w=2.86e-07 $l=3.3541e-07 $layer=POLY_cond $X=3.13 $Y=1.765
+ $X2=3.205 $Y2=1.465
r40 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.13 $Y=1.765
+ $X2=3.13 $Y2=2.4
r41 1 17 38.6549 $w=2.86e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.115 $Y=1.3
+ $X2=3.205 $Y2=1.465
r42 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.115 $Y=1.3 $X2=3.115
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__O41A_1%A1 1 3 6 8 9 14
r24 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.775
+ $Y=1.515 $X2=3.775 $Y2=1.515
r25 8 9 7.56494 $w=5.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.902 $Y=1.665
+ $X2=3.902 $Y2=2.035
r26 8 14 3.06687 $w=5.83e-07 $l=1.5e-07 $layer=LI1_cond $X=3.902 $Y=1.665
+ $X2=3.902 $Y2=1.515
r27 4 13 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=3.825 $Y=1.35
+ $X2=3.775 $Y2=1.515
r28 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.825 $Y=1.35
+ $X2=3.825 $Y2=0.69
r29 1 13 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=3.7 $Y=1.765
+ $X2=3.775 $Y2=1.515
r30 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.7 $Y=1.765 $X2=3.7
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O41A_1%X 1 2 9 13 14 15 26 28
r21 14 28 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=0.28 $Y=2.455 $X2=0.28
+ $Y2=2.405
r22 14 28 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=0.28 $Y=2.387
+ $X2=0.28 $Y2=2.405
r23 14 26 6.08745 $w=3.28e-07 $l=9.7e-08 $layer=LI1_cond $X=0.28 $Y=2.387
+ $X2=0.28 $Y2=2.29
r24 14 15 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.28 $Y=2.455
+ $X2=0.28 $Y2=2.775
r25 13 26 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=0.2 $Y=1.13 $X2=0.2
+ $Y2=2.29
r26 7 13 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.245 $Y=1 $X2=0.245
+ $Y2=1.13
r27 7 9 21.4975 $w=2.58e-07 $l=4.85e-07 $layer=LI1_cond $X=0.245 $Y=1 $X2=0.245
+ $Y2=0.515
r28 2 14 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.455
r29 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O41A_1%VPWR 1 2 9 12 14 16 18 23 32 36
r43 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r44 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r45 30 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r46 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r47 27 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 26 29 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r49 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 24 32 15.7083 $w=1.7e-07 $l=4.63e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.077 $Y2=3.33
r51 24 26 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 23 35 5.79967 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=3.76 $Y=3.33 $X2=4.04
+ $Y2=3.33
r53 23 29 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.76 $Y=3.33 $X2=3.6
+ $Y2=3.33
r54 21 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 18 32 15.7083 $w=1.7e-07 $l=4.62e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.077 $Y2=3.33
r57 18 20 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 16 30 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r59 16 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 12 35 2.96198 $w=4.45e-07 $l=1.1025e-07 $layer=LI1_cond $X=3.982 $Y=3.245
+ $X2=4.04 $Y2=3.33
r61 12 14 21.754 $w=4.43e-07 $l=8.4e-07 $layer=LI1_cond $X=3.982 $Y=3.245
+ $X2=3.982 $Y2=2.405
r62 7 32 3.39807 $w=9.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.077 $Y=3.245
+ $X2=1.077 $Y2=3.33
r63 7 9 11.4746 $w=9.23e-07 $l=8.7e-07 $layer=LI1_cond $X=1.077 $Y=3.245
+ $X2=1.077 $Y2=2.375
r64 2 14 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=3.775
+ $Y=1.84 $X2=3.925 $Y2=2.405
r65 1 9 300 $w=1.7e-07 $l=1.02828e-06 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=1.375 $Y2=2.375
r66 1 9 300 $w=1.7e-07 $l=6.27077e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LS__O41A_1%VGND 1 2 3 12 16 20 23 24 25 27 39 45 46 49
+ 52
r56 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r57 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r58 46 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r59 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r60 43 52 11.6921 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.44
+ $Y2=0
r61 43 45 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=4.08
+ $Y2=0
r62 42 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r63 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r64 39 52 11.6921 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.44
+ $Y2=0
r65 39 41 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.12
+ $Y2=0
r66 35 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r67 34 37 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r68 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r69 32 49 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.745
+ $Y2=0
r70 32 34 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r71 30 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r72 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r73 27 49 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.745
+ $Y2=0
r74 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r75 25 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r76 25 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r77 25 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r78 23 37 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.175 $Y=0 $X2=2.16
+ $Y2=0
r79 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=0 $X2=2.34
+ $Y2=0
r80 22 41 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.505 $Y=0 $X2=3.12
+ $Y2=0
r81 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=0 $X2=2.34
+ $Y2=0
r82 18 52 2.222 $w=5.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=0.085 $X2=3.44
+ $Y2=0
r83 18 20 9.70403 $w=5.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.44 $Y=0.085
+ $X2=3.44 $Y2=0.515
r84 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.085
+ $X2=2.34 $Y2=0
r85 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.34 $Y=0.085
+ $X2=2.34 $Y2=0.515
r86 10 49 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0
r87 10 12 11.8125 $w=3.98e-07 $l=4.1e-07 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0.495
r88 3 20 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=3.19
+ $Y=0.37 $X2=3.44 $Y2=0.515
r89 2 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.13
+ $Y=0.37 $X2=2.34 $Y2=0.515
r90 1 12 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LS__O41A_1%A_326_74# 1 2 3 12 14 15 18 20 24 26
r52 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.04 $Y=0.85
+ $X2=4.04 $Y2=0.515
r53 21 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=0.935
+ $X2=2.84 $Y2=0.935
r54 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.875 $Y=0.935
+ $X2=4.04 $Y2=0.85
r55 20 21 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=3.875 $Y=0.935
+ $X2=3.005 $Y2=0.935
r56 16 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=0.85 $X2=2.84
+ $Y2=0.935
r57 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.84 $Y=0.85
+ $X2=2.84 $Y2=0.515
r58 14 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=0.935
+ $X2=2.84 $Y2=0.935
r59 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.675 $Y=0.935
+ $X2=2.005 $Y2=0.935
r60 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.84 $Y=0.85
+ $X2=2.005 $Y2=0.935
r61 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.84 $Y=0.85
+ $X2=1.84 $Y2=0.515
r62 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.9
+ $Y=0.37 $X2=4.04 $Y2=0.515
r63 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.37 $X2=2.84 $Y2=0.515
r64 1 12 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.63
+ $Y=0.37 $X2=1.84 $Y2=0.515
.ends

