* File: sky130_fd_sc_ls__o21bai_1.pxi.spice
* Created: Fri Aug 28 13:46:27 2020
* 
x_PM_SKY130_FD_SC_LS__O21BAI_1%B1_N N_B1_N_M1002_g N_B1_N_c_60_n N_B1_N_M1000_g
+ B1_N N_B1_N_c_61_n PM_SKY130_FD_SC_LS__O21BAI_1%B1_N
x_PM_SKY130_FD_SC_LS__O21BAI_1%A_27_74# N_A_27_74#_M1002_s N_A_27_74#_M1000_s
+ N_A_27_74#_c_91_n N_A_27_74#_c_92_n N_A_27_74#_c_102_n N_A_27_74#_M1007_g
+ N_A_27_74#_M1004_g N_A_27_74#_c_94_n N_A_27_74#_c_95_n N_A_27_74#_c_103_n
+ N_A_27_74#_c_96_n N_A_27_74#_c_97_n N_A_27_74#_c_104_n N_A_27_74#_c_105_n
+ N_A_27_74#_c_98_n N_A_27_74#_c_99_n N_A_27_74#_c_100_n
+ PM_SKY130_FD_SC_LS__O21BAI_1%A_27_74#
x_PM_SKY130_FD_SC_LS__O21BAI_1%A2 N_A2_c_169_n N_A2_M1001_g N_A2_M1005_g A2 A2
+ A2 A2 A2 PM_SKY130_FD_SC_LS__O21BAI_1%A2
x_PM_SKY130_FD_SC_LS__O21BAI_1%A1 N_A1_c_209_n N_A1_M1006_g N_A1_M1003_g A1
+ N_A1_c_211_n PM_SKY130_FD_SC_LS__O21BAI_1%A1
x_PM_SKY130_FD_SC_LS__O21BAI_1%VPWR N_VPWR_M1000_d N_VPWR_M1006_d N_VPWR_c_234_n
+ N_VPWR_c_235_n N_VPWR_c_236_n VPWR N_VPWR_c_237_n N_VPWR_c_238_n
+ N_VPWR_c_239_n N_VPWR_c_233_n PM_SKY130_FD_SC_LS__O21BAI_1%VPWR
x_PM_SKY130_FD_SC_LS__O21BAI_1%Y N_Y_M1004_s N_Y_M1007_d N_Y_c_266_n N_Y_c_267_n
+ Y Y Y Y N_Y_c_268_n PM_SKY130_FD_SC_LS__O21BAI_1%Y
x_PM_SKY130_FD_SC_LS__O21BAI_1%VGND N_VGND_M1002_d N_VGND_M1005_d N_VGND_c_311_n
+ N_VGND_c_312_n VGND N_VGND_c_313_n N_VGND_c_314_n N_VGND_c_315_n
+ N_VGND_c_316_n N_VGND_c_317_n N_VGND_c_318_n PM_SKY130_FD_SC_LS__O21BAI_1%VGND
x_PM_SKY130_FD_SC_LS__O21BAI_1%A_308_74# N_A_308_74#_M1004_d N_A_308_74#_M1003_d
+ N_A_308_74#_c_349_n N_A_308_74#_c_350_n N_A_308_74#_c_351_n
+ N_A_308_74#_c_352_n PM_SKY130_FD_SC_LS__O21BAI_1%A_308_74#
cc_1 VNB N_B1_N_M1002_g 0.0548074f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.645
cc_2 VNB N_B1_N_c_60_n 0.0206119f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.045
cc_3 VNB N_B1_N_c_61_n 0.0105252f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.615
cc_4 VNB N_A_27_74#_c_91_n 0.0183564f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.54
cc_5 VNB N_A_27_74#_c_92_n 0.0102546f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.615
cc_6 VNB N_A_27_74#_M1004_g 0.0258899f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.615
cc_7 VNB N_A_27_74#_c_94_n 0.00625039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_95_n 0.0328912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_96_n 0.00635589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_97_n 0.0100794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_98_n 0.0194928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_99_n 4.49976e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_100_n 0.0361426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_169_n 0.029833f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.45
cc_15 VNB N_A2_M1005_g 0.0218673f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.54
cc_16 VNB A2 0.00676042f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_17 VNB A2 9.9768e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_209_n 0.0601748f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.45
cc_19 VNB N_A1_M1003_g 0.0294024f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.54
cc_20 VNB N_A1_c_211_n 0.00431187f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.615
cc_21 VNB N_VPWR_c_233_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_266_n 0.00782665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_267_n 0.00507195f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_24 VNB N_Y_c_268_n 0.00363505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_311_n 0.014848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_312_n 0.00396562f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_27 VNB N_VGND_c_313_n 0.0172318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_314_n 0.0312347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_315_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_316_n 0.196523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_317_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_318_n 0.00622543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_308_74#_c_349_n 0.00178852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_308_74#_c_350_n 0.0121113f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.615
cc_35 VNB N_A_308_74#_c_351_n 0.0048099f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.615
cc_36 VNB N_A_308_74#_c_352_n 0.0247745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_B1_N_c_60_n 0.0619145f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.045
cc_38 VPB N_B1_N_c_61_n 0.0070275f $X=-0.19 $Y=1.66 $X2=0.4 $Y2=1.615
cc_39 VPB N_A_27_74#_c_92_n 9.32055e-19 $X=-0.19 $Y=1.66 $X2=0.425 $Y2=1.615
cc_40 VPB N_A_27_74#_c_102_n 0.0238006f $X=-0.19 $Y=1.66 $X2=0.4 $Y2=1.615
cc_41 VPB N_A_27_74#_c_103_n 0.035396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_27_74#_c_104_n 0.00680148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_27_74#_c_105_n 0.00956337f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_27_74#_c_99_n 0.00568781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A2_c_169_n 0.0235602f $X=-0.19 $Y=1.66 $X2=0.49 $Y2=1.45
cc_46 VPB A2 0.00309847f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A1_c_209_n 0.0269279f $X=-0.19 $Y=1.66 $X2=0.49 $Y2=1.45
cc_48 VPB N_A1_c_211_n 0.00955428f $X=-0.19 $Y=1.66 $X2=0.4 $Y2=1.615
cc_49 VPB N_VPWR_c_234_n 0.013502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_235_n 0.0103902f $X=-0.19 $Y=1.66 $X2=0.4 $Y2=1.615
cc_51 VPB N_VPWR_c_236_n 0.0498232f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_52 VPB N_VPWR_c_237_n 0.0197879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_238_n 0.0342718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_239_n 0.0128614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_233_n 0.0633384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB Y 0.00945395f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB Y 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_Y_c_268_n 0.00204394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 N_B1_N_M1002_g N_A_27_74#_c_95_n 0.0108396f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_60 N_B1_N_c_60_n N_A_27_74#_c_103_n 0.0178576f $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_61 N_B1_N_M1002_g N_A_27_74#_c_96_n 0.0172243f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_62 N_B1_N_c_60_n N_A_27_74#_c_96_n 0.00212244f $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_63 N_B1_N_c_61_n N_A_27_74#_c_96_n 0.0148079f $X=0.4 $Y=1.615 $X2=0 $Y2=0
cc_64 N_B1_N_c_60_n N_A_27_74#_c_97_n 0.00291196f $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_65 N_B1_N_c_61_n N_A_27_74#_c_97_n 0.0202724f $X=0.4 $Y=1.615 $X2=0 $Y2=0
cc_66 N_B1_N_c_60_n N_A_27_74#_c_104_n 0.0140874f $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_67 N_B1_N_c_61_n N_A_27_74#_c_104_n 0.00710736f $X=0.4 $Y=1.615 $X2=0 $Y2=0
cc_68 N_B1_N_c_60_n N_A_27_74#_c_105_n 0.00967823f $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_69 N_B1_N_c_61_n N_A_27_74#_c_105_n 0.0280174f $X=0.4 $Y=1.615 $X2=0 $Y2=0
cc_70 N_B1_N_M1002_g N_A_27_74#_c_98_n 0.00425012f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_71 N_B1_N_c_60_n N_A_27_74#_c_98_n 6.31941e-19 $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_72 N_B1_N_c_61_n N_A_27_74#_c_98_n 0.014171f $X=0.4 $Y=1.615 $X2=0 $Y2=0
cc_73 N_B1_N_c_60_n N_A_27_74#_c_99_n 0.00705846f $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_74 N_B1_N_c_61_n N_A_27_74#_c_99_n 0.0109803f $X=0.4 $Y=1.615 $X2=0 $Y2=0
cc_75 N_B1_N_M1002_g N_A_27_74#_c_100_n 0.0173988f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_76 N_B1_N_c_61_n N_A_27_74#_c_100_n 2.01862e-19 $X=0.4 $Y=1.615 $X2=0 $Y2=0
cc_77 N_B1_N_c_60_n N_VPWR_c_234_n 0.0187219f $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_78 N_B1_N_c_60_n N_VPWR_c_237_n 0.00445602f $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_79 N_B1_N_c_60_n N_VPWR_c_233_n 0.00865278f $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_80 N_B1_N_M1002_g N_Y_c_266_n 0.0014725f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_81 N_B1_N_M1002_g N_Y_c_267_n 0.00454738f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_82 N_B1_N_c_60_n Y 3.69817e-19 $X=0.525 $Y=2.045 $X2=0 $Y2=0
cc_83 N_B1_N_M1002_g N_VGND_c_311_n 0.018223f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_84 N_B1_N_M1002_g N_VGND_c_313_n 0.00383152f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_85 N_B1_N_M1002_g N_VGND_c_316_n 0.0076118f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_86 N_A_27_74#_c_92_n N_A2_c_169_n 0.00589358f $X=1.45 $Y=1.675 $X2=-0.19
+ $Y2=-0.245
cc_87 N_A_27_74#_c_102_n N_A2_c_169_n 0.0105139f $X=1.45 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_88 N_A_27_74#_c_94_n N_A2_c_169_n 0.0208451f $X=1.45 $Y=1.375 $X2=-0.19
+ $Y2=-0.245
cc_89 N_A_27_74#_M1004_g N_A2_M1005_g 0.0135343f $X=1.465 $Y=0.74 $X2=0 $Y2=0
cc_90 N_A_27_74#_c_94_n A2 0.00121312f $X=1.45 $Y=1.375 $X2=0 $Y2=0
cc_91 N_A_27_74#_c_104_n N_VPWR_M1000_d 0.00188126f $X=0.745 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_92 N_A_27_74#_c_102_n N_VPWR_c_234_n 0.0204823f $X=1.45 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A_27_74#_c_103_n N_VPWR_c_234_n 0.0267702f $X=0.3 $Y=2.265 $X2=0 $Y2=0
cc_94 N_A_27_74#_c_104_n N_VPWR_c_234_n 0.0233603f $X=0.745 $Y=2.035 $X2=0 $Y2=0
cc_95 N_A_27_74#_c_98_n N_VPWR_c_234_n 0.00622181f $X=0.83 $Y=1.63 $X2=0 $Y2=0
cc_96 N_A_27_74#_c_100_n N_VPWR_c_234_n 0.00166955f $X=0.97 $Y=1.375 $X2=0 $Y2=0
cc_97 N_A_27_74#_c_103_n N_VPWR_c_237_n 0.0145938f $X=0.3 $Y=2.265 $X2=0 $Y2=0
cc_98 N_A_27_74#_c_102_n N_VPWR_c_238_n 0.00405947f $X=1.45 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_27_74#_c_102_n N_VPWR_c_233_n 0.00734183f $X=1.45 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A_27_74#_c_103_n N_VPWR_c_233_n 0.0120466f $X=0.3 $Y=2.265 $X2=0 $Y2=0
cc_101 N_A_27_74#_M1004_g N_Y_c_266_n 0.0107219f $X=1.465 $Y=0.74 $X2=0 $Y2=0
cc_102 N_A_27_74#_c_91_n N_Y_c_267_n 0.00697146f $X=1.36 $Y=1.375 $X2=0 $Y2=0
cc_103 N_A_27_74#_M1004_g N_Y_c_267_n 0.00313748f $X=1.465 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A_27_74#_c_98_n N_Y_c_267_n 0.00594309f $X=0.83 $Y=1.63 $X2=0 $Y2=0
cc_105 N_A_27_74#_c_100_n N_Y_c_267_n 3.87822e-19 $X=0.97 $Y=1.375 $X2=0 $Y2=0
cc_106 N_A_27_74#_c_102_n Y 0.013815f $X=1.45 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A_27_74#_c_104_n Y 0.0019861f $X=0.745 $Y=2.035 $X2=0 $Y2=0
cc_108 N_A_27_74#_c_102_n Y 0.0204739f $X=1.45 $Y=1.765 $X2=0 $Y2=0
cc_109 N_A_27_74#_c_104_n Y 0.00448737f $X=0.745 $Y=2.035 $X2=0 $Y2=0
cc_110 N_A_27_74#_c_91_n N_Y_c_268_n 0.00528353f $X=1.36 $Y=1.375 $X2=0 $Y2=0
cc_111 N_A_27_74#_c_92_n N_Y_c_268_n 0.00579483f $X=1.45 $Y=1.675 $X2=0 $Y2=0
cc_112 N_A_27_74#_c_102_n N_Y_c_268_n 0.00594287f $X=1.45 $Y=1.765 $X2=0 $Y2=0
cc_113 N_A_27_74#_M1004_g N_Y_c_268_n 0.00642503f $X=1.465 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A_27_74#_c_94_n N_Y_c_268_n 0.00362444f $X=1.45 $Y=1.375 $X2=0 $Y2=0
cc_115 N_A_27_74#_c_98_n N_Y_c_268_n 0.0326327f $X=0.83 $Y=1.63 $X2=0 $Y2=0
cc_116 N_A_27_74#_c_99_n N_Y_c_268_n 0.0138307f $X=0.83 $Y=1.95 $X2=0 $Y2=0
cc_117 N_A_27_74#_c_100_n N_Y_c_268_n 5.3485e-19 $X=0.97 $Y=1.375 $X2=0 $Y2=0
cc_118 N_A_27_74#_M1004_g N_VGND_c_311_n 0.00394308f $X=1.465 $Y=0.74 $X2=0
+ $Y2=0
cc_119 N_A_27_74#_c_95_n N_VGND_c_311_n 0.0226023f $X=0.275 $Y=0.645 $X2=0 $Y2=0
cc_120 N_A_27_74#_c_96_n N_VGND_c_311_n 0.0169933f $X=0.745 $Y=1.195 $X2=0 $Y2=0
cc_121 N_A_27_74#_c_98_n N_VGND_c_311_n 0.0116183f $X=0.83 $Y=1.63 $X2=0 $Y2=0
cc_122 N_A_27_74#_c_100_n N_VGND_c_311_n 3.25717e-19 $X=0.97 $Y=1.375 $X2=0
+ $Y2=0
cc_123 N_A_27_74#_M1004_g N_VGND_c_312_n 6.23092e-19 $X=1.465 $Y=0.74 $X2=0
+ $Y2=0
cc_124 N_A_27_74#_c_95_n N_VGND_c_313_n 0.011066f $X=0.275 $Y=0.645 $X2=0 $Y2=0
cc_125 N_A_27_74#_M1004_g N_VGND_c_314_n 0.00366292f $X=1.465 $Y=0.74 $X2=0
+ $Y2=0
cc_126 N_A_27_74#_M1004_g N_VGND_c_316_n 0.00606692f $X=1.465 $Y=0.74 $X2=0
+ $Y2=0
cc_127 N_A_27_74#_c_95_n N_VGND_c_316_n 0.00915947f $X=0.275 $Y=0.645 $X2=0
+ $Y2=0
cc_128 N_A_27_74#_M1004_g N_A_308_74#_c_349_n 0.00187536f $X=1.465 $Y=0.74 $X2=0
+ $Y2=0
cc_129 N_A_27_74#_M1004_g N_A_308_74#_c_351_n 6.78975e-19 $X=1.465 $Y=0.74 $X2=0
+ $Y2=0
cc_130 N_A2_c_169_n N_A1_c_209_n 0.0636297f $X=1.9 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_131 A2 N_A1_c_209_n 0.00280484f $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_132 A2 N_A1_c_209_n 0.00819469f $X=2.16 $Y=1.665 $X2=-0.19 $Y2=-0.245
cc_133 N_A2_M1005_g N_A1_M1003_g 0.031308f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A2_c_169_n N_A1_c_211_n 2.28131e-19 $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_135 A2 N_A1_c_211_n 0.0270733f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_136 A2 N_A1_c_211_n 0.0114994f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_137 N_A2_c_169_n N_VPWR_c_238_n 0.00445602f $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_138 A2 N_VPWR_c_238_n 0.00682779f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_139 N_A2_c_169_n N_VPWR_c_233_n 0.00858782f $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_140 A2 N_VPWR_c_233_n 0.00794958f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_141 N_A2_M1005_g N_Y_c_267_n 9.65872e-19 $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A2_c_169_n Y 0.00402647f $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_143 A2 Y 0.0068392f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_144 A2 Y 0.0708234f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_145 N_A2_c_169_n Y 0.0119373f $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A2_c_169_n N_Y_c_268_n 0.00103807f $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_147 A2 N_Y_c_268_n 0.0165956f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_148 A2 N_Y_c_268_n 0.00552603f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_149 A2 A_395_368# 0.0238323f $X=2.16 $Y=1.665 $X2=-0.19 $Y2=-0.245
cc_150 N_A2_M1005_g N_VGND_c_312_n 0.00803907f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A2_M1005_g N_VGND_c_314_n 0.00383152f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A2_M1005_g N_VGND_c_316_n 0.00758084f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A2_M1005_g N_A_308_74#_c_349_n 4.4413e-19 $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A2_c_169_n N_A_308_74#_c_350_n 0.00276992f $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A2_M1005_g N_A_308_74#_c_350_n 0.0125718f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_156 A2 N_A_308_74#_c_350_n 0.0347779f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A2_c_169_n N_A_308_74#_c_351_n 0.00152246f $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_158 A2 N_A_308_74#_c_351_n 0.00548166f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_159 N_A1_c_209_n N_VPWR_c_236_n 0.0119352f $X=2.38 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A1_c_211_n N_VPWR_c_236_n 0.022248f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_161 N_A1_c_209_n N_VPWR_c_238_n 0.00461464f $X=2.38 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A1_c_209_n N_VPWR_c_233_n 0.00912775f $X=2.38 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A1_c_209_n Y 7.27818e-19 $X=2.38 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A1_M1003_g N_VGND_c_312_n 0.0107652f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A1_M1003_g N_VGND_c_315_n 0.00383152f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A1_M1003_g N_VGND_c_316_n 0.00761198f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A1_c_209_n N_A_308_74#_c_350_n 0.00315952f $X=2.38 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A1_M1003_g N_A_308_74#_c_350_n 0.0169051f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A1_c_211_n N_A_308_74#_c_350_n 0.0270164f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_170 N_A1_M1003_g N_A_308_74#_c_352_n 0.00159319f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_171 N_VPWR_M1000_d Y 0.0028151f $X=0.6 $Y=2.12 $X2=0 $Y2=0
cc_172 N_VPWR_c_234_n Y 0.0570768f $X=1.14 $Y=2.455 $X2=0 $Y2=0
cc_173 N_VPWR_c_238_n Y 0.0160091f $X=2.52 $Y=3.33 $X2=0 $Y2=0
cc_174 N_VPWR_c_233_n Y 0.0131029f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_175 N_Y_c_266_n N_VGND_c_311_n 0.0421766f $X=1.25 $Y=0.515 $X2=0 $Y2=0
cc_176 N_Y_c_266_n N_VGND_c_314_n 0.0170618f $X=1.25 $Y=0.515 $X2=0 $Y2=0
cc_177 N_Y_c_266_n N_VGND_c_316_n 0.013925f $X=1.25 $Y=0.515 $X2=0 $Y2=0
cc_178 N_Y_c_266_n N_A_308_74#_c_349_n 0.0455845f $X=1.25 $Y=0.515 $X2=0 $Y2=0
cc_179 N_Y_c_267_n N_A_308_74#_c_351_n 0.0142394f $X=1.28 $Y=1.13 $X2=0 $Y2=0
cc_180 N_VGND_c_312_n N_A_308_74#_c_349_n 0.0125684f $X=2.165 $Y=0.515 $X2=0
+ $Y2=0
cc_181 N_VGND_c_314_n N_A_308_74#_c_349_n 0.00749631f $X=1.995 $Y=0 $X2=0 $Y2=0
cc_182 N_VGND_c_316_n N_A_308_74#_c_349_n 0.0062048f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_183 N_VGND_M1005_d N_A_308_74#_c_350_n 0.00234908f $X=2.02 $Y=0.37 $X2=0
+ $Y2=0
cc_184 N_VGND_c_312_n N_A_308_74#_c_350_n 0.0122946f $X=2.165 $Y=0.515 $X2=0
+ $Y2=0
cc_185 N_VGND_c_312_n N_A_308_74#_c_352_n 0.0126098f $X=2.165 $Y=0.515 $X2=0
+ $Y2=0
cc_186 N_VGND_c_315_n N_A_308_74#_c_352_n 0.011066f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_187 N_VGND_c_316_n N_A_308_74#_c_352_n 0.00915947f $X=2.64 $Y=0 $X2=0 $Y2=0
