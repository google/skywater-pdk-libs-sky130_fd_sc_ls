* File: sky130_fd_sc_ls__or4b_2.spice
* Created: Fri Aug 28 14:00:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__or4b_2.pex.spice"
.subckt sky130_fd_sc_ls__or4b_2  VNB VPB D_N A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_D_N_M1009_g N_A_27_368#_M1009_s VNB NSHORT L=0.15 W=0.55
+ AD=0.109083 AS=0.15675 PD=0.942248 PS=1.67 NRD=18.54 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75003.5 A=0.0825 P=1.4 MULT=1
MM1004 N_X_M1004_d N_A_190_48#_M1004_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.146767 PD=1.02 PS=1.26775 NRD=0 NRS=0.804 M=1 R=4.93333
+ SA=75000.6 SB=75002.7 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1004_d N_A_190_48#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.164409 PD=1.02 PS=1.26551 NRD=0 NRS=18.648 M=1 R=4.93333
+ SA=75001 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1003 N_A_190_48#_M1003_d N_A_M1003_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1408 AS=0.142191 PD=1.08 PS=1.09449 NRD=14.988 NRS=8.436 M=1 R=4.26667
+ SA=75001.7 SB=75002 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_B_M1006_g N_A_190_48#_M1003_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1584 AS=0.1408 PD=1.135 PS=1.08 NRD=17.808 NRS=14.988 M=1 R=4.26667
+ SA=75002.3 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1002 N_A_190_48#_M1002_d N_C_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.64
+ AD=0.104 AS=0.1584 PD=0.965 PS=1.135 NRD=8.436 NRS=22.488 M=1 R=4.26667
+ SA=75002.9 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1010 N_VGND_M1010_d N_A_27_368#_M1010_g N_A_190_48#_M1002_d VNB NSHORT L=0.15
+ W=0.64 AD=0.2272 AS=0.104 PD=1.99 PS=0.965 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75003.4 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_D_N_M1005_g N_A_27_368#_M1005_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.174 AS=0.2478 PD=1.29 PS=2.27 NRD=35.6767 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75003.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1005_d N_A_190_48#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.232 AS=0.168 PD=1.72 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_190_48#_M1011_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.304725 AS=0.168 PD=1.75925 PS=1.42 NRD=22.852 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1012 A_452_392# N_A_M1012_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.272075 PD=1.27 PS=1.57075 NRD=15.7403 NRS=26.5753 M=1 R=6.66667
+ SA=75001.8 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1007 A_536_392# N_B_M1007_g A_452_392# VPB PHIGHVT L=0.15 W=1 AD=0.18 AS=0.135
+ PD=1.36 PS=1.27 NRD=24.6053 NRS=15.7403 M=1 R=6.66667 SA=75002.2 SB=75001.4
+ A=0.15 P=2.3 MULT=1
MM1008 A_638_392# N_C_M1008_g A_536_392# VPB PHIGHVT L=0.15 W=1 AD=0.195 AS=0.18
+ PD=1.39 PS=1.36 NRD=27.5603 NRS=24.6053 M=1 R=6.66667 SA=75002.7 SB=75000.9
+ A=0.15 P=2.3 MULT=1
MM1001 N_A_190_48#_M1001_d N_A_27_368#_M1001_g A_638_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.445 AS=0.195 PD=2.89 PS=1.39 NRD=31.5003 NRS=27.5603 M=1 R=6.66667
+ SA=75003.2 SB=75000.4 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
c_52 VNB 0 1.7764e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__or4b_2.pxi.spice"
*
.ends
*
*
