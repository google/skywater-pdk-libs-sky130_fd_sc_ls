* File: sky130_fd_sc_ls__nor4_1.pxi.spice
* Created: Fri Aug 28 13:39:35 2020
* 
x_PM_SKY130_FD_SC_LS__NOR4_1%A N_A_c_48_n N_A_M1007_g N_A_M1000_g N_A_c_45_n
+ N_A_c_46_n A N_A_c_47_n PM_SKY130_FD_SC_LS__NOR4_1%A
x_PM_SKY130_FD_SC_LS__NOR4_1%B N_B_c_70_n N_B_M1002_g N_B_M1004_g B B B B
+ N_B_c_72_n PM_SKY130_FD_SC_LS__NOR4_1%B
x_PM_SKY130_FD_SC_LS__NOR4_1%C N_C_c_107_n N_C_M1003_g N_C_M1005_g C C
+ N_C_c_109_n PM_SKY130_FD_SC_LS__NOR4_1%C
x_PM_SKY130_FD_SC_LS__NOR4_1%D N_D_M1006_g N_D_c_139_n N_D_M1001_g D N_D_c_140_n
+ PM_SKY130_FD_SC_LS__NOR4_1%D
x_PM_SKY130_FD_SC_LS__NOR4_1%VPWR N_VPWR_M1007_s N_VPWR_c_166_n N_VPWR_c_167_n
+ VPWR N_VPWR_c_168_n N_VPWR_c_165_n PM_SKY130_FD_SC_LS__NOR4_1%VPWR
x_PM_SKY130_FD_SC_LS__NOR4_1%Y N_Y_M1000_d N_Y_M1005_d N_Y_M1001_d N_Y_c_189_n
+ N_Y_c_190_n N_Y_c_191_n N_Y_c_192_n N_Y_c_193_n N_Y_c_194_n N_Y_c_196_n
+ N_Y_c_195_n Y PM_SKY130_FD_SC_LS__NOR4_1%Y
x_PM_SKY130_FD_SC_LS__NOR4_1%VGND N_VGND_M1000_s N_VGND_M1004_d N_VGND_M1006_d
+ N_VGND_c_245_n N_VGND_c_246_n N_VGND_c_247_n N_VGND_c_248_n N_VGND_c_249_n
+ N_VGND_c_250_n N_VGND_c_251_n VGND N_VGND_c_252_n N_VGND_c_253_n
+ PM_SKY130_FD_SC_LS__NOR4_1%VGND
cc_1 VNB N_A_c_45_n 0.0638345f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.385
cc_2 VNB N_A_c_46_n 0.0211013f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.22
cc_3 VNB N_A_c_47_n 0.0240277f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.385
cc_4 VNB N_B_c_70_n 0.0251381f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.765
cc_5 VNB N_B_M1004_g 0.0267613f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=0.74
cc_6 VNB N_B_c_72_n 0.00390329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_C_c_107_n 0.0269867f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.765
cc_8 VNB N_C_M1005_g 0.026814f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=0.74
cc_9 VNB N_C_c_109_n 0.00167078f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.385
cc_10 VNB N_D_M1006_g 0.0264948f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.4
cc_11 VNB N_D_c_139_n 0.0270607f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=0.74
cc_12 VNB N_D_c_140_n 0.00419952f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.385
cc_13 VNB N_VPWR_c_165_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_Y_c_189_n 0.00215184f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.385
cc_15 VNB N_Y_c_190_n 0.0100809f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.385
cc_16 VNB N_Y_c_191_n 0.00906721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_192_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_193_n 0.0227193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_194_n 0.00789082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_195_n 0.0230393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_245_n 0.016404f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_22 VNB N_VGND_c_246_n 0.0351944f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.385
cc_23 VNB N_VGND_c_247_n 0.00900448f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_24 VNB N_VGND_c_248_n 0.0162041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_249_n 0.0323694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_250_n 0.0168561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_251_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_252_n 0.021877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_253_n 0.193176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_A_c_48_n 0.0188098f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.765
cc_31 VPB N_A_c_45_n 0.010078f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=1.385
cc_32 VPB N_B_c_70_n 0.0271179f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.765
cc_33 VPB N_B_c_72_n 0.00202152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_C_c_107_n 0.028714f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.765
cc_35 VPB N_C_c_109_n 0.00186046f $X=-0.19 $Y=1.66 $X2=0.375 $Y2=1.385
cc_36 VPB N_D_c_139_n 0.0327367f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=0.74
cc_37 VPB N_D_c_140_n 0.00647557f $X=-0.19 $Y=1.66 $X2=0.375 $Y2=1.385
cc_38 VPB N_VPWR_c_166_n 0.0164764f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.22
cc_39 VPB N_VPWR_c_167_n 0.0559563f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=0.74
cc_40 VPB N_VPWR_c_168_n 0.0687575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_165_n 0.0929982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_Y_c_196_n 0.0138831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_Y_c_195_n 0.0142968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB Y 0.040652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 N_A_c_48_n N_B_c_70_n 0.0581866f $X=0.645 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_46 N_A_c_45_n N_B_c_70_n 0.0230778f $X=0.555 $Y=1.385 $X2=-0.19 $Y2=-0.245
cc_47 N_A_c_47_n N_B_c_70_n 5.45707e-19 $X=0.375 $Y=1.385 $X2=-0.19 $Y2=-0.245
cc_48 N_A_c_46_n N_B_M1004_g 0.0190702f $X=0.645 $Y=1.22 $X2=0 $Y2=0
cc_49 N_A_c_47_n N_B_M1004_g 5.55714e-19 $X=0.375 $Y=1.385 $X2=0 $Y2=0
cc_50 N_A_c_48_n N_B_c_72_n 0.00419518f $X=0.645 $Y=1.765 $X2=0 $Y2=0
cc_51 N_A_c_45_n N_B_c_72_n 0.00231033f $X=0.555 $Y=1.385 $X2=0 $Y2=0
cc_52 N_A_c_47_n N_B_c_72_n 0.00713992f $X=0.375 $Y=1.385 $X2=0 $Y2=0
cc_53 N_A_c_48_n N_VPWR_c_167_n 0.0237051f $X=0.645 $Y=1.765 $X2=0 $Y2=0
cc_54 N_A_c_45_n N_VPWR_c_167_n 0.00763465f $X=0.555 $Y=1.385 $X2=0 $Y2=0
cc_55 N_A_c_47_n N_VPWR_c_167_n 0.0170992f $X=0.375 $Y=1.385 $X2=0 $Y2=0
cc_56 N_A_c_48_n N_VPWR_c_168_n 0.00413917f $X=0.645 $Y=1.765 $X2=0 $Y2=0
cc_57 N_A_c_48_n N_VPWR_c_165_n 0.00817532f $X=0.645 $Y=1.765 $X2=0 $Y2=0
cc_58 N_A_c_46_n N_Y_c_189_n 4.03226e-19 $X=0.645 $Y=1.22 $X2=0 $Y2=0
cc_59 N_A_c_46_n N_Y_c_191_n 0.00221478f $X=0.645 $Y=1.22 $X2=0 $Y2=0
cc_60 N_A_c_45_n N_VGND_c_246_n 0.00230739f $X=0.555 $Y=1.385 $X2=0 $Y2=0
cc_61 N_A_c_46_n N_VGND_c_246_n 0.0131164f $X=0.645 $Y=1.22 $X2=0 $Y2=0
cc_62 N_A_c_47_n N_VGND_c_246_n 0.0282557f $X=0.375 $Y=1.385 $X2=0 $Y2=0
cc_63 N_A_c_46_n N_VGND_c_250_n 0.00383152f $X=0.645 $Y=1.22 $X2=0 $Y2=0
cc_64 N_A_c_46_n N_VGND_c_253_n 0.00757637f $X=0.645 $Y=1.22 $X2=0 $Y2=0
cc_65 N_B_c_70_n N_C_c_107_n 0.0538351f $X=1.065 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_66 N_B_c_72_n N_C_c_107_n 0.0211023f $X=1.14 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_67 N_B_M1004_g N_C_M1005_g 0.0195058f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_68 N_B_c_70_n N_C_c_109_n 9.13071e-19 $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_69 N_B_c_72_n N_C_c_109_n 0.0412959f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_70 N_B_c_70_n N_VPWR_c_167_n 0.00208978f $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_71 N_B_c_72_n N_VPWR_c_167_n 0.021024f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_72 N_B_c_70_n N_VPWR_c_168_n 0.00303293f $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_73 N_B_c_72_n N_VPWR_c_168_n 0.00941005f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_74 N_B_c_70_n N_VPWR_c_165_n 0.00372936f $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_75 N_B_c_72_n N_VPWR_c_165_n 0.0110375f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_76 N_B_c_72_n A_228_368# 0.0145694f $X=1.14 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_77 N_B_M1004_g N_Y_c_189_n 0.00968448f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_78 N_B_c_70_n N_Y_c_190_n 9.86927e-19 $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_79 N_B_M1004_g N_Y_c_190_n 0.012155f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_80 N_B_c_72_n N_Y_c_190_n 0.0214362f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_81 N_B_c_70_n N_Y_c_191_n 3.05922e-19 $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_82 N_B_M1004_g N_Y_c_191_n 0.00139157f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_83 N_B_c_72_n N_Y_c_191_n 0.0055933f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_84 N_B_M1004_g N_Y_c_192_n 8.51666e-19 $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_85 N_B_M1004_g N_VGND_c_246_n 5.57151e-19 $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_86 N_B_M1004_g N_VGND_c_247_n 0.00543742f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_87 N_B_M1004_g N_VGND_c_250_n 0.00434272f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_88 N_B_M1004_g N_VGND_c_253_n 0.00822072f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_89 N_C_M1005_g N_D_M1006_g 0.0200614f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_90 N_C_c_107_n N_D_c_139_n 0.0576964f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_91 N_C_c_109_n N_D_c_139_n 0.00623452f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_92 N_C_c_107_n N_D_c_140_n 0.00230565f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_93 N_C_c_109_n N_D_c_140_n 0.0349696f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_94 N_C_c_107_n N_VPWR_c_168_n 0.00461464f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_95 N_C_c_107_n N_VPWR_c_165_n 0.00911823f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_96 N_C_c_109_n A_342_368# 0.00880286f $X=1.71 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_97 N_C_M1005_g N_Y_c_189_n 8.12002e-19 $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_98 N_C_c_107_n N_Y_c_190_n 9.67719e-19 $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_99 N_C_M1005_g N_Y_c_190_n 0.012155f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_100 N_C_c_109_n N_Y_c_190_n 0.0205962f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_101 N_C_M1005_g N_Y_c_192_n 0.0111642f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_102 N_C_c_107_n N_Y_c_194_n 3.08675e-19 $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_103 N_C_M1005_g N_Y_c_194_n 0.0015571f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_104 N_C_c_109_n N_Y_c_194_n 0.0055933f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_105 N_C_c_107_n N_Y_c_196_n 0.00387653f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_106 N_C_c_109_n N_Y_c_196_n 0.00847445f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_107 N_C_M1005_g N_VGND_c_247_n 0.00782003f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_108 N_C_M1005_g N_VGND_c_252_n 0.00434272f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_109 N_C_M1005_g N_VGND_c_253_n 0.00823282f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_110 N_D_c_139_n N_VPWR_c_168_n 0.00445602f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_111 N_D_c_139_n N_VPWR_c_165_n 0.00863343f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_112 N_D_M1006_g N_Y_c_192_n 0.01371f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_113 N_D_M1006_g N_Y_c_193_n 0.0129505f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_114 N_D_c_139_n N_Y_c_193_n 0.00126003f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_115 N_D_c_140_n N_Y_c_193_n 0.0229301f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_116 N_D_M1006_g N_Y_c_194_n 0.0015571f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_117 N_D_c_140_n N_Y_c_194_n 0.00829487f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_118 N_D_c_139_n N_Y_c_196_n 0.00517443f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_119 N_D_c_140_n N_Y_c_196_n 0.013098f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_120 N_D_M1006_g N_Y_c_195_n 0.00477786f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_121 N_D_c_139_n N_Y_c_195_n 0.0123296f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_122 N_D_c_140_n N_Y_c_195_n 0.0332226f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_123 N_D_c_139_n Y 0.0164322f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_124 N_D_M1006_g N_VGND_c_249_n 0.00722118f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_125 N_D_M1006_g N_VGND_c_252_n 0.00434272f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_126 N_D_M1006_g N_VGND_c_253_n 0.0082432f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_127 N_VPWR_c_168_n Y 0.0230718f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_128 N_VPWR_c_165_n Y 0.0190639f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_129 N_Y_c_190_n N_VGND_M1004_d 0.00764236f $X=1.81 $Y=1.095 $X2=0 $Y2=0
cc_130 N_Y_c_193_n N_VGND_M1006_d 0.0024352f $X=2.615 $Y=1.095 $X2=0 $Y2=0
cc_131 N_Y_c_189_n N_VGND_c_246_n 0.0262671f $X=0.875 $Y=0.515 $X2=0 $Y2=0
cc_132 N_Y_c_189_n N_VGND_c_247_n 0.0185169f $X=0.875 $Y=0.515 $X2=0 $Y2=0
cc_133 N_Y_c_190_n N_VGND_c_247_n 0.0257907f $X=1.81 $Y=1.095 $X2=0 $Y2=0
cc_134 N_Y_c_192_n N_VGND_c_247_n 0.0267123f $X=1.975 $Y=0.515 $X2=0 $Y2=0
cc_135 N_Y_c_192_n N_VGND_c_249_n 0.0191765f $X=1.975 $Y=0.515 $X2=0 $Y2=0
cc_136 N_Y_c_193_n N_VGND_c_249_n 0.0263592f $X=2.615 $Y=1.095 $X2=0 $Y2=0
cc_137 N_Y_c_189_n N_VGND_c_250_n 0.0114405f $X=0.875 $Y=0.515 $X2=0 $Y2=0
cc_138 N_Y_c_192_n N_VGND_c_252_n 0.0144922f $X=1.975 $Y=0.515 $X2=0 $Y2=0
cc_139 N_Y_c_189_n N_VGND_c_253_n 0.00941304f $X=0.875 $Y=0.515 $X2=0 $Y2=0
cc_140 N_Y_c_192_n N_VGND_c_253_n 0.0118826f $X=1.975 $Y=0.515 $X2=0 $Y2=0
