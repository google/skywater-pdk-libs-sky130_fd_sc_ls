* File: sky130_fd_sc_ls__a2bb2oi_2.spice
* Created: Fri Aug 28 12:56:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a2bb2oi_2.pex.spice"
.subckt sky130_fd_sc_ls__a2bb2oi_2  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1010 N_A_212_102#_M1010_d N_A1_N_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15
+ W=0.64 AD=0.104 AS=0.1696 PD=0.965 PS=1.81 NRD=3.744 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1008_d N_A2_N_M1008_g N_A_212_102#_M1010_d VNB NSHORT L=0.15
+ W=0.64 AD=0.113206 AS=0.104 PD=1.00174 PS=0.965 NRD=11.244 NRS=4.68 M=1
+ R=4.26667 SA=75000.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1004 N_Y_M1004_d N_A_212_102#_M1004_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.130894 PD=1.02 PS=1.15826 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1011 N_Y_M1004_d N_A_212_102#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_B2_M1002_g N_A_615_74#_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1002_d N_B2_M1007_g N_A_615_74#_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1006 N_A_615_74#_M1007_s N_B1_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1014 N_A_615_74#_M1014_d N_B1_M1014_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 A_209_392# N_A1_N_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1 AD=0.12
+ AS=0.275 PD=1.24 PS=2.55 NRD=12.7853 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1013 N_A_212_102#_M1013_d N_A2_N_M1013_g A_209_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.275 AS=0.12 PD=2.55 PS=1.24 NRD=1.9503 NRS=12.7853 M=1 R=6.66667
+ SA=75000.6 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_A_424_368#_M1001_d N_A_212_102#_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1015 N_A_424_368#_M1015_d N_A_212_102#_M1015_g N_Y_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75002 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1003_d N_B2_M1003_g N_A_424_368#_M1015_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1003_d N_B2_M1009_g N_A_424_368#_M1009_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1000 N_A_424_368#_M1009_s N_B1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1012 N_A_424_368#_M1012_d N_B1_M1012_g N_VPWR_M1000_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.4 SB=75000.2 A=0.168 P=2.54 MULT=1
DX16_noxref VNB VPB NWDIODE A=10.5276 P=15.04
c_55 VNB 0 1.56524e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__a2bb2oi_2.pxi.spice"
*
.ends
*
*
