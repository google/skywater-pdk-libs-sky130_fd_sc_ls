# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__o21a_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__o21a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.300000 2.775000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.715000 1.445000 2.275000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.445000 1.435000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.350000 0.365000 1.820000 ;
        RECT 0.115000 1.820000 0.445000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 2.880000 0.085000 ;
        RECT 0.545000  0.085000 0.875000 0.935000 ;
        RECT 2.005000  0.085000 2.335000 0.790000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 2.880000 3.415000 ;
        RECT 0.615000 2.290000 1.180000 3.245000 ;
        RECT 2.435000 1.950000 2.765000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.535000 1.105000 1.395000 1.275000 ;
      RECT 0.535000 1.275000 0.865000 1.550000 ;
      RECT 0.695000 1.550000 0.865000 1.950000 ;
      RECT 0.695000 1.950000 1.690000 2.120000 ;
      RECT 1.145000 0.350000 1.395000 1.105000 ;
      RECT 1.360000 2.120000 1.690000 2.795000 ;
      RECT 1.575000 0.350000 1.825000 0.960000 ;
      RECT 1.575000 0.960000 2.765000 1.130000 ;
      RECT 2.515000 0.350000 2.765000 0.960000 ;
  END
END sky130_fd_sc_ls__o21a_1
