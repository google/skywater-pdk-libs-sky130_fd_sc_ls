* File: sky130_fd_sc_ls__nand2_1.pex.spice
* Created: Wed Sep  2 11:11:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__NAND2_1%B 1 3 4 6 7
r23 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r24 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r25 4 10 38.924 $w=3.61e-07 $l=2.33345e-07 $layer=POLY_cond $X=0.51 $Y=1.22
+ $X2=0.345 $Y2=1.385
r26 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.51 $Y=1.22 $X2=0.51
+ $Y2=0.74
r27 1 10 67.6304 $w=3.61e-07 $l=4.48776e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.345 $Y2=1.385
r28 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__NAND2_1%A 1 3 4 6 7
r23 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.385 $X2=1.17 $Y2=1.385
r24 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.17 $Y=1.295 $X2=1.17
+ $Y2=1.385
r25 4 10 66.5442 $w=3.79e-07 $l=4.4238e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=1.08 $Y2=1.385
r26 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=2.4
r27 1 10 39.2012 $w=3.79e-07 $l=2.49199e-07 $layer=POLY_cond $X=0.9 $Y=1.22
+ $X2=1.08 $Y2=1.385
r28 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.9 $Y=1.22 $X2=0.9
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__NAND2_1%VPWR 1 2 7 9 13 15 19 21 31
r21 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r22 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r23 22 27 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r24 22 24 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r25 21 30 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.222 $Y2=3.33
r26 21 24 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 19 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r28 19 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r29 19 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 15 18 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.17 $Y=1.985
+ $X2=1.17 $Y2=2.815
r31 13 30 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.222 $Y2=3.33
r32 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.815
r33 9 12 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.27 $Y=1.985
+ $X2=0.27 $Y2=2.815
r34 7 27 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r35 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.815
r36 2 18 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=2.815
r37 2 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=1.985
r38 1 12 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.815
r39 1 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__NAND2_1%Y 1 2 9 11 17 18 19 20 21 30 44
r30 20 21 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=2.405
+ $X2=0.72 $Y2=2.775
r31 19 20 21.0446 $w=2.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.72 $Y=1.985
+ $X2=0.72 $Y2=2.405
r32 18 19 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=0.72 $Y2=1.985
r33 17 30 2.15457 $w=2.28e-07 $l=4.3e-08 $layer=LI1_cond $X=0.72 $Y=1.252
+ $X2=0.72 $Y2=1.295
r34 17 44 4.41536 $w=2.28e-07 $l=7.2e-08 $layer=LI1_cond $X=0.72 $Y=1.252
+ $X2=0.72 $Y2=1.18
r35 17 18 16.4348 $w=2.28e-07 $l=3.28e-07 $layer=LI1_cond $X=0.72 $Y=1.337
+ $X2=0.72 $Y2=1.665
r36 17 30 2.10446 $w=2.28e-07 $l=4.2e-08 $layer=LI1_cond $X=0.72 $Y=1.337
+ $X2=0.72 $Y2=1.295
r37 9 13 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.115 $Y=0.925
+ $X2=0.75 $Y2=0.925
r38 9 11 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.115 $Y=0.84
+ $X2=1.115 $Y2=0.515
r39 7 13 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=1.01 $X2=0.75
+ $Y2=0.925
r40 7 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.75 $Y=1.01 $X2=0.75
+ $Y2=1.18
r41 2 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.815
r42 2 19 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=1.985
r43 1 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.975
+ $Y=0.37 $X2=1.115 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__NAND2_1%VGND 1 4 6 8 12 13
r17 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r18 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r19 10 16 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=0 $X2=0.23
+ $Y2=0
r20 10 12 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.46 $Y=0 $X2=1.2
+ $Y2=0
r21 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r22 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r23 4 16 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.23 $Y2=0
r24 4 6 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.295 $Y2=0.515
r25 1 6 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends

