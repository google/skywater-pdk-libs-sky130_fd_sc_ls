* File: sky130_fd_sc_ls__nand4_4.spice
* Created: Wed Sep  2 11:13:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nand4_4.pex.spice"
.subckt sky130_fd_sc_ls__nand4_4  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_D_M1007_g N_A_27_74#_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.7 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1007_d N_D_M1009_g N_A_27_74#_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.7
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_D_M1014_g N_A_27_74#_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2035 AS=0.1295 PD=1.29 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1014_d N_D_M1018_g N_A_27_74#_M1018_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2035 AS=0.1295 PD=1.29 PS=1.09 NRD=32.424 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1001 N_A_554_74#_M1001_d N_C_M1001_g N_A_27_74#_M1018_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75002.4 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1010 N_A_554_74#_M1001_d N_C_M1010_g N_A_27_74#_M1010_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.8 SB=75001 A=0.111 P=1.78 MULT=1
MM1012 N_A_554_74#_M1012_d N_C_M1012_g N_A_27_74#_M1010_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.3 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1019 N_A_554_74#_M1012_d N_C_M1019_g N_A_27_74#_M1019_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.19515 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_923_74#_M1004_d N_B_M1004_g N_A_554_74#_M1004_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1969 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.4 A=0.111 P=1.78 MULT=1
MM1006 N_A_923_74#_M1006_d N_B_M1006_g N_A_554_74#_M1004_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002.9 A=0.111 P=1.78 MULT=1
MM1017 N_A_923_74#_M1006_d N_B_M1017_g N_A_554_74#_M1017_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1021 N_A_923_74#_M1021_d N_B_M1021_g N_A_554_74#_M1017_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g N_A_923_74#_M1021_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1003_d N_A_M1013_g N_A_923_74#_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1015 N_Y_M1015_d N_A_M1015_g N_A_923_74#_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1628 AS=0.1036 PD=1.18 PS=1.02 NRD=12.972 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1023 N_Y_M1015_d N_A_M1023_g N_A_923_74#_M1023_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1628 AS=0.1962 PD=1.18 PS=2.05 NRD=12.972 NRS=0 M=1 R=4.93333 SA=75003.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_D_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12 AD=0.196
+ AS=1.736 PD=1.47 PS=5.34 NRD=1.7533 NRS=2.6201 M=1 R=7.46667 SA=75001.5
+ SB=75006.6 A=0.168 P=2.54 MULT=1
MM1005 N_Y_M1000_d N_D_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.12 AD=0.196
+ AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75006.1 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1011_d N_C_M1011_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3808 AS=0.168 PD=1.8 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.4 SB=75005.6 A=0.168 P=2.54 MULT=1
MM1020 N_Y_M1011_d N_C_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3808 AS=0.4872 PD=1.8 PS=1.99 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.3 SB=75004.8 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1020_s N_B_M1016_g N_Y_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.4872 AS=0.3808 PD=1.99 PS=1.8 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.3 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1022 N_VPWR_M1022_d N_B_M1022_g N_Y_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.9296 AS=0.3808 PD=2.78 PS=1.8 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.1 SB=75003 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1022_d N_A_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.9296 AS=0.4368 PD=2.78 PS=1.9 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.9 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.4368 PD=2.83 PS=1.9 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.8 SB=75000.2 A=0.168 P=2.54 MULT=1
DX24_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_ls__nand4_4.pxi.spice"
*
.ends
*
*
