* File: sky130_fd_sc_ls__decaphe_8.pex.spice
* Created: Wed Sep  2 11:00:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DECAPHE_8%VGND 1 7 13 28 31
r10 30 31 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.6 $Y=0
+ $X2=3.6 $Y2=0
r11 28 30 0.183459 $w=1.33e-06 $l=2e-08 $layer=LI1_cond $X=3.58 $Y=0.757 $X2=3.6
+ $Y2=0.757
r12 23 24 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r13 21 23 4.21955 $w=1.33e-06 $l=4.6e-07 $layer=LI1_cond $X=0.26 $Y=0.757
+ $X2=0.72 $Y2=0.757
r14 19 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r15 18 21 0.183459 $w=1.33e-06 $l=2e-08 $layer=LI1_cond $X=0.24 $Y=0.757
+ $X2=0.26 $Y2=0.757
r16 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r17 16 28 9.67744 $w=1.33e-06 $l=1.055e-06 $layer=LI1_cond $X=2.525 $Y=0.757
+ $X2=3.58 $Y2=0.757
r18 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.525
+ $Y=1.515 $X2=2.525 $Y2=1.515
r19 13 15 18.2029 $w=1.602e-06 $l=6.05e-07 $layer=POLY_cond $X=1.92 $Y=2.287
+ $X2=2.525 $Y2=2.287
r20 11 16 16.1444 $w=1.33e-06 $l=1.76e-06 $layer=LI1_cond $X=0.765 $Y=0.757
+ $X2=2.525 $Y2=0.757
r21 11 23 0.412782 $w=1.33e-06 $l=4.5e-08 $layer=LI1_cond $X=0.765 $Y=0.757
+ $X2=0.72 $Y2=0.757
r22 10 13 34.7509 $w=1.602e-06 $l=1.155e-06 $layer=POLY_cond $X=0.765 $Y=2.287
+ $X2=1.92 $Y2=2.287
r23 10 11 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.765
+ $Y=1.515 $X2=0.765 $Y2=1.515
r24 7 31 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.6
+ $Y2=0
r25 7 24 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=0.72
+ $Y2=0
r26 1 28 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.445
+ $Y=0.235 $X2=3.58 $Y2=0.38
r27 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=3.445
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LS__DECAPHE_8%VPWR 1 7 8 10 11 28 36
r12 28 31 0.136009 $w=1.794e-06 $l=2e-08 $layer=LI1_cond $X=3.58 $Y=2.332
+ $X2=3.6 $Y2=2.332
r13 21 36 0.00397135 $w=3.84e-06 $l=1.22e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.92 $Y2=3.208
r14 21 31 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r15 20 23 0.136009 $w=1.794e-06 $l=2e-08 $layer=LI1_cond $X=0.24 $Y=2.332
+ $X2=0.26 $Y2=2.332
r16 20 21 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r17 18 28 1.19008 $w=1.794e-06 $l=1.75e-07 $layer=LI1_cond $X=3.405 $Y=2.332
+ $X2=3.58 $Y2=2.332
r18 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.405
+ $Y=1.335 $X2=3.405 $Y2=1.335
r19 15 18 11.9688 $w=1.794e-06 $l=1.76e-06 $layer=LI1_cond $X=1.645 $Y=2.332
+ $X2=3.405 $Y2=2.332
r20 15 23 9.41862 $w=1.794e-06 $l=1.385e-06 $layer=LI1_cond $X=1.645 $Y=2.332
+ $X2=0.26 $Y2=2.332
r21 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.645
+ $Y=1.335 $X2=1.645 $Y2=1.335
r22 11 36 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=3.207
+ $X2=1.92 $Y2=3.208
r23 8 14 7.69394 $w=1.205e-06 $l=2.49199e-07 $layer=POLY_cond $X=1.81 $Y=0.622
+ $X2=1.645 $Y2=0.802
r24 8 10 5.46463 $w=1.035e-06 $l=1.1e-07 $layer=POLY_cond $X=1.81 $Y=0.622
+ $X2=1.92 $Y2=0.622
r25 7 17 21.3213 $w=1.201e-06 $l=5.88154e-07 $layer=POLY_cond $X=2.9 $Y=0.622
+ $X2=3.405 $Y2=0.802
r26 7 10 48.6848 $w=1.035e-06 $l=9.8e-07 $layer=POLY_cond $X=2.9 $Y=0.622
+ $X2=1.92 $Y2=0.622
r27 1 28 400 $w=1.7e-07 $l=1.17556e-06 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.84 $X2=3.58 $Y2=2.95
r28 1 28 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.84 $X2=3.58 $Y2=1.985
r29 1 23 400 $w=1.7e-07 $l=1.17083e-06 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.84 $X2=0.26 $Y2=2.95
r30 1 23 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.84 $X2=0.26 $Y2=1.985
.ends

