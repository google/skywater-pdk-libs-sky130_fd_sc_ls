* File: sky130_fd_sc_ls__o21ba_4.pex.spice
* Created: Fri Aug 28 13:46:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O21BA_4%B1_N 1 3 4 6 7
r33 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.385 $X2=0.59 $Y2=1.385
r34 7 11 4.04912 $w=3.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.59 $Y2=1.365
r35 4 10 38.7914 $w=2.76e-07 $l=1.92678e-07 $layer=POLY_cond $X=0.525 $Y=1.22
+ $X2=0.585 $Y2=1.385
r36 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.525 $Y=1.22 $X2=0.525
+ $Y2=0.74
r37 1 10 76.3385 $w=2.76e-07 $l=4.18091e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.585 $Y2=1.385
r38 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_4%A_193_48# 1 2 3 12 14 16 19 21 23 26 28 30
+ 33 35 37 38 47 48 49 50 56 59 60 62 64 66 68 79
c163 50 0 9.42363e-21 $X=3.66 $Y=1.375
c164 33 0 7.8786e-20 $X=2.34 $Y=0.74
c165 12 0 1.76934e-19 $X=1.04 $Y=0.74
r166 79 80 8.11658 $w=3.86e-07 $l=6.5e-08 $layer=POLY_cond $X=2.34 $Y=1.527
+ $X2=2.405 $Y2=1.527
r167 76 77 5.61917 $w=3.86e-07 $l=4.5e-08 $layer=POLY_cond $X=1.91 $Y=1.527
+ $X2=1.955 $Y2=1.527
r168 73 74 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=1.48 $Y=1.527
+ $X2=1.505 $Y2=1.527
r169 72 73 53.0699 $w=3.86e-07 $l=4.25e-07 $layer=POLY_cond $X=1.055 $Y=1.527
+ $X2=1.48 $Y2=1.527
r170 71 72 1.87306 $w=3.86e-07 $l=1.5e-08 $layer=POLY_cond $X=1.04 $Y=1.527
+ $X2=1.055 $Y2=1.527
r171 62 70 5.34211 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.06 $Y=2.3
+ $X2=5.06 $Y2=2.125
r172 62 64 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.06 $Y=2.3 $X2=5.06
+ $Y2=2.57
r173 61 68 0.414005 $w=3.5e-07 $l=3.42491e-07 $layer=LI1_cond $X=3.83 $Y=2.125
+ $X2=3.49 $Y2=2.13
r174 60 70 2.59474 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.975 $Y=2.125
+ $X2=5.06 $Y2=2.125
r175 60 61 37.7014 $w=3.48e-07 $l=1.145e-06 $layer=LI1_cond $X=4.975 $Y=2.125
+ $X2=3.83 $Y2=2.125
r176 59 68 7.71803 $w=2.1e-07 $l=3.33054e-07 $layer=LI1_cond $X=3.745 $Y=1.95
+ $X2=3.49 $Y2=2.13
r177 58 59 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.745 $Y=1.46
+ $X2=3.745 $Y2=1.95
r178 54 56 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.665 $Y=0.425
+ $X2=3.665 $Y2=0.615
r179 51 66 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.98 $Y=1.375
+ $X2=2.895 $Y2=1.455
r180 50 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.66 $Y=1.375
+ $X2=3.745 $Y2=1.46
r181 50 51 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.66 $Y=1.375
+ $X2=2.98 $Y2=1.375
r182 48 54 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.5 $Y=0.34
+ $X2=3.665 $Y2=0.425
r183 48 49 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.5 $Y=0.34
+ $X2=2.98 $Y2=0.34
r184 47 66 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=1.29
+ $X2=2.895 $Y2=1.455
r185 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.895 $Y=0.425
+ $X2=2.98 $Y2=0.34
r186 46 47 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.895 $Y=0.425
+ $X2=2.895 $Y2=1.29
r187 45 79 1.2487 $w=3.86e-07 $l=1e-08 $layer=POLY_cond $X=2.33 $Y=1.527
+ $X2=2.34 $Y2=1.527
r188 45 77 46.8264 $w=3.86e-07 $l=3.75e-07 $layer=POLY_cond $X=2.33 $Y=1.527
+ $X2=1.955 $Y2=1.527
r189 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.33
+ $Y=1.455 $X2=2.33 $Y2=1.455
r190 41 76 32.4663 $w=3.86e-07 $l=2.6e-07 $layer=POLY_cond $X=1.65 $Y=1.527
+ $X2=1.91 $Y2=1.527
r191 41 74 18.1062 $w=3.86e-07 $l=1.45e-07 $layer=POLY_cond $X=1.65 $Y=1.527
+ $X2=1.505 $Y2=1.527
r192 40 44 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.65 $Y=1.455
+ $X2=2.33 $Y2=1.455
r193 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.455 $X2=1.65 $Y2=1.455
r194 38 66 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=1.455
+ $X2=2.895 $Y2=1.455
r195 38 44 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.81 $Y=1.455
+ $X2=2.33 $Y2=1.455
r196 35 80 24.9932 $w=1.5e-07 $l=2.38e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=1.527
r197 35 37 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=2.4
r198 31 79 24.9932 $w=1.5e-07 $l=2.37e-07 $layer=POLY_cond $X=2.34 $Y=1.29
+ $X2=2.34 $Y2=1.527
r199 31 33 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.34 $Y=1.29
+ $X2=2.34 $Y2=0.74
r200 28 77 24.9932 $w=1.5e-07 $l=2.38e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.955 $Y2=1.527
r201 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.955 $Y2=2.4
r202 24 76 24.9932 $w=1.5e-07 $l=2.37e-07 $layer=POLY_cond $X=1.91 $Y=1.29
+ $X2=1.91 $Y2=1.527
r203 24 26 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.91 $Y=1.29
+ $X2=1.91 $Y2=0.74
r204 21 74 24.9932 $w=1.5e-07 $l=2.38e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=1.527
r205 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=2.4
r206 17 73 24.9932 $w=1.5e-07 $l=2.37e-07 $layer=POLY_cond $X=1.48 $Y=1.29
+ $X2=1.48 $Y2=1.527
r207 17 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.48 $Y=1.29
+ $X2=1.48 $Y2=0.74
r208 14 72 24.9932 $w=1.5e-07 $l=2.38e-07 $layer=POLY_cond $X=1.055 $Y=1.765
+ $X2=1.055 $Y2=1.527
r209 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.055 $Y=1.765
+ $X2=1.055 $Y2=2.4
r210 10 71 24.9932 $w=1.5e-07 $l=2.37e-07 $layer=POLY_cond $X=1.04 $Y=1.29
+ $X2=1.04 $Y2=1.527
r211 10 12 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.04 $Y=1.29
+ $X2=1.04 $Y2=0.74
r212 3 70 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.96 $X2=5.06 $Y2=2.115
r213 3 64 600 $w=1.7e-07 $l=6.80882e-07 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.96 $X2=5.06 $Y2=2.57
r214 2 68 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=3.425
+ $Y=2.12 $X2=3.575 $Y2=2.295
r215 1 56 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.525
+ $Y=0.47 $X2=3.665 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_4%A_27_368# 1 2 7 9 12 14 16 19 23 28 31 33 36
+ 37 39 40 41 45 51
c99 23 0 1.76934e-19 $X=0.31 $Y=0.515
r100 51 52 10.9235 $w=3.53e-07 $l=8e-08 $layer=POLY_cond $X=3.8 $Y=1.837
+ $X2=3.88 $Y2=1.837
r101 50 51 47.7904 $w=3.53e-07 $l=3.5e-07 $layer=POLY_cond $X=3.45 $Y=1.837
+ $X2=3.8 $Y2=1.837
r102 49 50 13.6544 $w=3.53e-07 $l=1e-07 $layer=POLY_cond $X=3.35 $Y=1.837
+ $X2=3.45 $Y2=1.837
r103 46 49 3.4136 $w=3.53e-07 $l=2.5e-08 $layer=POLY_cond $X=3.325 $Y=1.837
+ $X2=3.35 $Y2=1.837
r104 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.325
+ $Y=1.795 $X2=3.325 $Y2=1.795
r105 42 45 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.235 $Y=1.795
+ $X2=3.325 $Y2=1.795
r106 39 40 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=1.985
+ $X2=0.265 $Y2=1.82
r107 37 40 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.17 $Y=1.01
+ $X2=0.17 $Y2=1.82
r108 35 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.235 $Y=1.96
+ $X2=3.235 $Y2=1.795
r109 35 36 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.235 $Y=1.96
+ $X2=3.235 $Y2=2.39
r110 34 41 4.14084 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.445 $Y=2.475
+ $X2=0.265 $Y2=2.475
r111 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.15 $Y=2.475
+ $X2=3.235 $Y2=2.39
r112 33 34 176.476 $w=1.68e-07 $l=2.705e-06 $layer=LI1_cond $X=3.15 $Y=2.475
+ $X2=0.445 $Y2=2.475
r113 29 41 2.66603 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.56
+ $X2=0.265 $Y2=2.475
r114 29 31 8.16314 $w=3.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.265 $Y=2.56
+ $X2=0.265 $Y2=2.815
r115 28 41 2.66603 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.39
+ $X2=0.265 $Y2=2.475
r116 27 39 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.265 $Y=2
+ $X2=0.265 $Y2=1.985
r117 27 28 12.4848 $w=3.58e-07 $l=3.9e-07 $layer=LI1_cond $X=0.265 $Y=2
+ $X2=0.265 $Y2=2.39
r118 21 37 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=0.28 $Y=0.815
+ $X2=0.28 $Y2=1.01
r119 21 23 8.86495 $w=3.88e-07 $l=3e-07 $layer=LI1_cond $X=0.28 $Y=0.815
+ $X2=0.28 $Y2=0.515
r120 17 52 22.8335 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.88 $Y=1.63
+ $X2=3.88 $Y2=1.837
r121 17 19 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.88 $Y=1.63
+ $X2=3.88 $Y2=0.79
r122 14 51 22.8335 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.8 $Y=2.045
+ $X2=3.8 $Y2=1.837
r123 14 16 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.8 $Y=2.045
+ $X2=3.8 $Y2=2.54
r124 10 50 22.8335 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.45 $Y=1.63
+ $X2=3.45 $Y2=1.837
r125 10 12 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.45 $Y=1.63
+ $X2=3.45 $Y2=0.79
r126 7 49 22.8335 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.35 $Y=2.045
+ $X2=3.35 $Y2=1.837
r127 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.35 $Y=2.045
+ $X2=3.35 $Y2=2.54
r128 2 39 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r129 2 31 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r130 1 23 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.37 $X2=0.31 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_4%A2 1 3 6 8 10 13 15 16 17 26
c59 13 0 1.44963e-19 $X=5.31 $Y=0.945
c60 6 0 7.82385e-20 $X=4.88 $Y=0.945
r61 26 27 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=5.285 $Y=1.667
+ $X2=5.31 $Y2=1.667
r62 24 26 34.3394 $w=3.86e-07 $l=2.75e-07 $layer=POLY_cond $X=5.01 $Y=1.667
+ $X2=5.285 $Y2=1.667
r63 22 24 16.2332 $w=3.86e-07 $l=1.3e-07 $layer=POLY_cond $X=4.88 $Y=1.667
+ $X2=5.01 $Y2=1.667
r64 21 22 5.61917 $w=3.86e-07 $l=4.5e-08 $layer=POLY_cond $X=4.835 $Y=1.667
+ $X2=4.88 $Y2=1.667
r65 16 17 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.615 $X2=6
+ $Y2=1.615
r66 15 16 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=5.01 $Y=1.615
+ $X2=5.52 $Y2=1.615
r67 15 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.01
+ $Y=1.615 $X2=5.01 $Y2=1.615
r68 11 27 24.9932 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=5.31 $Y=1.45
+ $X2=5.31 $Y2=1.667
r69 11 13 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.31 $Y=1.45
+ $X2=5.31 $Y2=0.945
r70 8 26 24.9932 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=5.285 $Y=1.885
+ $X2=5.285 $Y2=1.667
r71 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.285 $Y=1.885
+ $X2=5.285 $Y2=2.46
r72 4 22 24.9932 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=4.88 $Y=1.45
+ $X2=4.88 $Y2=1.667
r73 4 6 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.88 $Y=1.45 $X2=4.88
+ $Y2=0.945
r74 1 21 24.9932 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=4.835 $Y=1.885
+ $X2=4.835 $Y2=1.667
r75 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.835 $Y=1.885
+ $X2=4.835 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_4%A1 4 5 7 8 9 10 11 12 14 18 20
c70 5 0 9.42363e-21 $X=4.385 $Y=1.885
c71 4 0 4.38187e-20 $X=4.38 $Y=0.945
r72 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.34
+ $Y=1.615 $X2=4.34 $Y2=1.615
r73 20 24 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=4.56 $Y=1.615
+ $X2=4.34 $Y2=1.615
r74 18 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.74 $Y=0.945
+ $X2=5.74 $Y2=1.34
r75 15 18 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.74 $Y=0.255
+ $X2=5.74 $Y2=0.945
r76 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.735 $Y=1.885
+ $X2=5.735 $Y2=2.46
r77 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.735 $Y=1.795
+ $X2=5.735 $Y2=1.885
r78 10 19 36.2738 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.735 $Y=1.43
+ $X2=5.735 $Y2=1.34
r79 10 11 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=5.735 $Y=1.43
+ $X2=5.735 $Y2=1.795
r80 8 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.665 $Y=0.18
+ $X2=5.74 $Y2=0.255
r81 8 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=5.665 $Y=0.18
+ $X2=4.455 $Y2=0.18
r82 5 23 55.8646 $w=2.93e-07 $l=2.91633e-07 $layer=POLY_cond $X=4.385 $Y=1.885
+ $X2=4.34 $Y2=1.615
r83 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.385 $Y=1.885
+ $X2=4.385 $Y2=2.46
r84 2 23 38.5916 $w=2.93e-07 $l=1.83916e-07 $layer=POLY_cond $X=4.38 $Y=1.45
+ $X2=4.34 $Y2=1.615
r85 2 4 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.38 $Y=1.45 $X2=4.38
+ $Y2=0.945
r86 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.38 $Y=0.255
+ $X2=4.455 $Y2=0.18
r87 1 4 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.38 $Y=0.255 $X2=4.38
+ $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_4%VPWR 1 2 3 4 5 18 22 26 28 30 34 36 41 51 56
+ 65 68 72 76 78 82
r78 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r79 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r80 74 76 9.31175 $w=6.83e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=3.072
+ $X2=3.205 $Y2=3.072
r81 71 74 1.39688 $w=6.83e-07 $l=8e-08 $layer=LI1_cond $X=3.04 $Y=3.072 $X2=3.12
+ $Y2=3.072
r82 71 72 17.8676 $w=6.83e-07 $l=5.75e-07 $layer=LI1_cond $X=3.04 $Y=3.072
+ $X2=2.465 $Y2=3.072
r83 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r84 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r85 63 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r86 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r87 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r88 60 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r89 59 62 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=5.52
+ $Y2=3.33
r90 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r91 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.275 $Y=3.33
+ $X2=4.11 $Y2=3.33
r92 57 59 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.275 $Y=3.33
+ $X2=4.56 $Y2=3.33
r93 56 81 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=5.875 $Y=3.33
+ $X2=6.057 $Y2=3.33
r94 56 62 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.875 $Y=3.33
+ $X2=5.52 $Y2=3.33
r95 55 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r96 54 76 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=3.205 $Y2=3.33
r97 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r98 51 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=4.11 $Y2=3.33
r99 51 54 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=3.6 $Y2=3.33
r100 50 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r101 49 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=2.465 $Y2=3.33
r102 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r103 47 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=3.33
+ $X2=1.73 $Y2=3.33
r104 47 49 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.895 $Y=3.33
+ $X2=2.16 $Y2=3.33
r105 45 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r106 45 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r107 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r108 42 65 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=0.805 $Y2=3.33
r109 42 44 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=1.2 $Y2=3.33
r110 41 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.73 $Y2=3.33
r111 41 44 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.2 $Y2=3.33
r112 39 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r114 36 65 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.805 $Y2=3.33
r115 36 38 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r116 34 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r117 34 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r118 34 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r119 30 33 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=6 $Y=2.115 $X2=6
+ $Y2=2.815
r120 28 81 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=6 $Y=3.245
+ $X2=6.057 $Y2=3.33
r121 28 33 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6 $Y=3.245 $X2=6
+ $Y2=2.815
r122 24 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=3.33
r123 24 26 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=2.635
r124 20 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=3.245
+ $X2=1.73 $Y2=3.33
r125 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.73 $Y=3.245
+ $X2=1.73 $Y2=2.815
r126 16 65 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=3.33
r127 16 18 13.0408 $w=3.78e-07 $l=4.3e-07 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=2.815
r128 5 33 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=5.81
+ $Y=1.96 $X2=5.96 $Y2=2.815
r129 5 30 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=5.81
+ $Y=1.96 $X2=5.96 $Y2=2.115
r130 4 26 600 $w=1.7e-07 $l=6.2149e-07 $layer=licon1_PDIFF $count=1 $X=3.875
+ $Y=2.12 $X2=4.11 $Y2=2.635
r131 3 71 300 $w=1.7e-07 $l=1.22337e-06 $layer=licon1_PDIFF $count=2 $X=2.48
+ $Y=1.84 $X2=3.04 $Y2=2.815
r132 2 22 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.73 $Y2=2.815
r133 1 18 600 $w=1.7e-07 $l=1.08167e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.805 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_4%X 1 2 3 4 15 21 23 27 29 30 31 36 38 41
c52 30 0 4.78765e-20 $X=1.115 $Y=1.58
c53 23 0 7.8786e-20 $X=1.96 $Y=1.035
r54 31 36 4.75094 $w=2.3e-07 $l=2e-07 $layer=LI1_cond $X=1.2 $Y=2.02 $X2=1.2
+ $Y2=1.82
r55 30 38 2.15457 $w=2.28e-07 $l=4.3e-08 $layer=LI1_cond $X=1.2 $Y=1.622 $X2=1.2
+ $Y2=1.665
r56 30 41 4.41536 $w=2.28e-07 $l=7.2e-08 $layer=LI1_cond $X=1.2 $Y=1.622 $X2=1.2
+ $Y2=1.55
r57 30 36 5.662 $w=2.28e-07 $l=1.13e-07 $layer=LI1_cond $X=1.2 $Y=1.707 $X2=1.2
+ $Y2=1.82
r58 30 38 2.10446 $w=2.28e-07 $l=4.2e-08 $layer=LI1_cond $X=1.2 $Y=1.707 $X2=1.2
+ $Y2=1.665
r59 25 27 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=2.085 $Y=0.95
+ $X2=2.085 $Y2=0.515
r60 24 29 1.59926 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=1.34 $Y=1.035
+ $X2=1.242 $Y2=1.035
r61 23 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.96 $Y=1.035
+ $X2=2.085 $Y2=0.95
r62 23 24 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.96 $Y=1.035
+ $X2=1.34 $Y2=1.035
r63 19 31 2.73179 $w=4e-07 $l=1.15e-07 $layer=LI1_cond $X=1.315 $Y=2.02 $X2=1.2
+ $Y2=2.02
r64 19 21 24.9216 $w=3.98e-07 $l=8.65e-07 $layer=LI1_cond $X=1.315 $Y=2.02
+ $X2=2.18 $Y2=2.02
r65 17 29 4.86787 $w=1.82e-07 $l=9.0802e-08 $layer=LI1_cond $X=1.23 $Y=1.12
+ $X2=1.242 $Y2=1.035
r66 17 41 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.23 $Y=1.12
+ $X2=1.23 $Y2=1.55
r67 13 29 4.86787 $w=1.82e-07 $l=8.5e-08 $layer=LI1_cond $X=1.242 $Y=0.95
+ $X2=1.242 $Y2=1.035
r68 13 15 24.7413 $w=1.93e-07 $l=4.35e-07 $layer=LI1_cond $X=1.242 $Y=0.95
+ $X2=1.242 $Y2=0.515
r69 4 21 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.84 $X2=2.18 $Y2=2.02
r70 3 31 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.84 $X2=1.28 $Y2=2.02
r71 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.985
+ $Y=0.37 $X2=2.125 $Y2=0.515
r72 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.115
+ $Y=0.37 $X2=1.255 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_4%A_892_392# 1 2 9 11 12 15
r31 15 18 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=5.51 $Y=2.115 $X2=5.51
+ $Y2=2.815
r32 13 18 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.51 $Y=2.905 $X2=5.51
+ $Y2=2.815
r33 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.345 $Y=2.99
+ $X2=5.51 $Y2=2.905
r34 11 12 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.345 $Y=2.99
+ $X2=4.775 $Y2=2.99
r35 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.61 $Y=2.905
+ $X2=4.775 $Y2=2.99
r36 7 9 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=4.61 $Y=2.905 $X2=4.61
+ $Y2=2.635
r37 2 18 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=5.36
+ $Y=1.96 $X2=5.51 $Y2=2.815
r38 2 15 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=5.36
+ $Y=1.96 $X2=5.51 $Y2=2.115
r39 1 9 600 $w=1.7e-07 $l=7.46241e-07 $layer=licon1_PDIFF $count=1 $X=4.46
+ $Y=1.96 $X2=4.61 $Y2=2.635
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_4%VGND 1 2 3 4 5 20 24 28 32 36 39 40 41 43 52
+ 56 63 64 67 70 73 76
r91 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r92 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r93 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r94 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r95 64 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r96 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r97 61 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.61 $Y=0 $X2=5.485
+ $Y2=0
r98 61 63 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=5.61 $Y=0 $X2=6
+ $Y2=0
r99 60 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r100 60 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r101 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r102 57 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.625
+ $Y2=0
r103 57 59 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=5.04
+ $Y2=0
r104 56 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.36 $Y=0 $X2=5.485
+ $Y2=0
r105 56 59 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.36 $Y=0 $X2=5.04
+ $Y2=0
r106 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r107 52 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.5 $Y=0 $X2=4.625
+ $Y2=0
r108 52 54 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=4.5 $Y=0 $X2=2.64
+ $Y2=0
r109 51 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r110 51 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r111 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r112 48 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=1.655
+ $Y2=0
r113 48 50 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=2.16
+ $Y2=0
r114 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r115 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r116 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.81
+ $Y2=0
r118 44 46 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.2
+ $Y2=0
r119 43 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.53 $Y=0 $X2=1.655
+ $Y2=0
r120 43 46 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.53 $Y=0 $X2=1.2
+ $Y2=0
r121 41 74 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=4.56 $Y2=0
r122 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r123 40 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.515 $Y=0 $X2=2.64
+ $Y2=0
r124 39 50 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.16
+ $Y2=0
r125 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.515
+ $Y2=0
r126 34 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.485 $Y=0.085
+ $X2=5.485 $Y2=0
r127 34 36 31.5769 $w=2.48e-07 $l=6.85e-07 $layer=LI1_cond $X=5.485 $Y=0.085
+ $X2=5.485 $Y2=0.77
r128 30 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=0.085
+ $X2=4.625 $Y2=0
r129 30 32 31.5769 $w=2.48e-07 $l=6.85e-07 $layer=LI1_cond $X=4.625 $Y=0.085
+ $X2=4.625 $Y2=0.77
r130 26 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=0.085
+ $X2=2.515 $Y2=0
r131 26 28 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.515 $Y=0.085
+ $X2=2.515 $Y2=0.515
r132 22 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=0.085
+ $X2=1.655 $Y2=0
r133 22 24 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=1.655 $Y=0.085
+ $X2=1.655 $Y2=0.565
r134 18 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=0.085
+ $X2=0.81 $Y2=0
r135 18 20 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.81 $Y=0.085
+ $X2=0.81 $Y2=0.495
r136 5 36 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.385
+ $Y=0.625 $X2=5.525 $Y2=0.77
r137 4 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.455
+ $Y=0.625 $X2=4.665 $Y2=0.77
r138 3 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.415
+ $Y=0.37 $X2=2.555 $Y2=0.515
r139 2 24 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.37 $X2=1.695 $Y2=0.565
r140 1 20 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=0.6
+ $Y=0.37 $X2=0.81 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LS__O21BA_4%A_618_94# 1 2 3 4 15 17 18 19 22 26 28 32 34
+ 37
c61 34 0 7.82385e-20 $X=4.165 $Y=1.035
c62 26 0 1.44963e-19 $X=5.095 $Y=0.77
c63 17 0 4.38187e-20 $X=4 $Y=1.035
r64 34 35 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.165 $Y=1.035
+ $X2=4.165 $Y2=1.195
r65 30 32 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=5.957 $Y=1.11
+ $X2=5.957 $Y2=0.77
r66 29 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.18 $Y=1.195
+ $X2=5.055 $Y2=1.195
r67 28 30 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=5.79 $Y=1.195
+ $X2=5.957 $Y2=1.11
r68 28 29 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.79 $Y=1.195
+ $X2=5.18 $Y2=1.195
r69 24 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=1.11
+ $X2=5.055 $Y2=1.195
r70 24 26 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=5.055 $Y=1.11
+ $X2=5.055 $Y2=0.77
r71 23 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=1.195
+ $X2=4.165 $Y2=1.195
r72 22 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.93 $Y=1.195
+ $X2=5.055 $Y2=1.195
r73 22 23 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.93 $Y=1.195 $X2=4.33
+ $Y2=1.195
r74 19 34 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.165 $Y=0.95
+ $X2=4.165 $Y2=1.035
r75 19 21 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.165 $Y=0.95
+ $X2=4.165 $Y2=0.865
r76 17 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=1.035 $X2=4.165
+ $Y2=1.035
r77 17 18 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4 $Y=1.035 $X2=3.32
+ $Y2=1.035
r78 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.235 $Y=0.95
+ $X2=3.32 $Y2=1.035
r79 13 15 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.235 $Y=0.95
+ $X2=3.235 $Y2=0.855
r80 4 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.815
+ $Y=0.625 $X2=5.955 $Y2=0.77
r81 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.955
+ $Y=0.625 $X2=5.095 $Y2=0.77
r82 2 21 182 $w=1.7e-07 $l=4.88851e-07 $layer=licon1_NDIFF $count=1 $X=3.955
+ $Y=0.47 $X2=4.165 $Y2=0.865
r83 1 15 182 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_NDIFF $count=1 $X=3.09
+ $Y=0.47 $X2=3.235 $Y2=0.855
.ends

