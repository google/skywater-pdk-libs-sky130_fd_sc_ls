* File: sky130_fd_sc_ls__a32o_2.pex.spice
* Created: Wed Sep  2 10:52:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A32O_2%A_45_264# 1 2 7 9 12 14 16 19 22 23 24 26 28
+ 29 30 31 35 40 44 46 50
c110 14 0 1.20518e-19 $X=0.955 $Y=1.765
c111 7 0 3.688e-20 $X=0.505 $Y=1.765
r112 50 51 5.83065 $w=3.72e-07 $l=4.5e-08 $layer=POLY_cond $X=0.955 $Y=1.542
+ $X2=1 $Y2=1.542
r113 49 50 51.1801 $w=3.72e-07 $l=3.95e-07 $layer=POLY_cond $X=0.56 $Y=1.542
+ $X2=0.955 $Y2=1.542
r114 48 49 7.12634 $w=3.72e-07 $l=5.5e-08 $layer=POLY_cond $X=0.505 $Y=1.542
+ $X2=0.56 $Y2=1.542
r115 41 48 14.9005 $w=3.72e-07 $l=1.15e-07 $layer=POLY_cond $X=0.39 $Y=1.542
+ $X2=0.505 $Y2=1.542
r116 40 43 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.39 $Y=1.485
+ $X2=0.39 $Y2=1.65
r117 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.39
+ $Y=1.485 $X2=0.39 $Y2=1.485
r118 33 35 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.94 $Y=1.01
+ $X2=2.94 $Y2=0.515
r119 32 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.275 $Y=2.035
+ $X2=1.19 $Y2=2.035
r120 31 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=2.035
+ $X2=3.54 $Y2=2.035
r121 31 32 137.005 $w=1.68e-07 $l=2.1e-06 $layer=LI1_cond $X=3.375 $Y=2.035
+ $X2=1.275 $Y2=2.035
r122 29 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.775 $Y=1.095
+ $X2=2.94 $Y2=1.01
r123 29 30 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=2.775 $Y=1.095
+ $X2=1.275 $Y2=1.095
r124 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=2.12
+ $X2=1.19 $Y2=2.035
r125 27 28 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.19 $Y=2.12 $X2=1.19
+ $Y2=2.32
r126 26 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=1.95
+ $X2=1.19 $Y2=2.035
r127 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.19 $Y=1.18
+ $X2=1.275 $Y2=1.095
r128 25 26 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.19 $Y=1.18
+ $X2=1.19 $Y2=1.95
r129 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.105 $Y=2.405
+ $X2=1.19 $Y2=2.32
r130 23 24 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.105 $Y=2.405
+ $X2=0.395 $Y2=2.405
r131 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.31 $Y=2.32
+ $X2=0.395 $Y2=2.405
r132 22 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.31 $Y=2.32
+ $X2=0.31 $Y2=1.65
r133 17 51 24.0971 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1 $Y=1.32 $X2=1
+ $Y2=1.542
r134 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1 $Y=1.32 $X2=1
+ $Y2=0.74
r135 14 50 24.0971 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.542
r136 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r137 10 49 24.0971 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.56 $Y=1.32
+ $X2=0.56 $Y2=1.542
r138 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.56 $Y=1.32
+ $X2=0.56 $Y2=0.74
r139 7 48 24.0971 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.542
r140 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r141 2 46 300 $w=1.7e-07 $l=3.09233e-07 $layer=licon1_PDIFF $count=2 $X=3.34
+ $Y=1.84 $X2=3.54 $Y2=2.065
r142 1 35 91 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=2 $X=2.735
+ $Y=0.37 $X2=2.94 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A32O_2%A3 1 3 6 8 12
c31 6 0 1.22536e-19 $X=1.7 $Y=0.74
c32 1 0 1.42058e-19 $X=1.655 $Y=1.765
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.515 $X2=1.61 $Y2=1.515
r34 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.61 $Y=1.665
+ $X2=1.61 $Y2=1.515
r35 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.7 $Y=1.35
+ $X2=1.61 $Y2=1.515
r36 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.7 $Y=1.35 $X2=1.7
+ $Y2=0.74
r37 1 11 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=1.655 $Y=1.765
+ $X2=1.61 $Y2=1.515
r38 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.655 $Y=1.765
+ $X2=1.655 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LS__A32O_2%A2 3 5 7 8 12
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.18
+ $Y=1.515 $X2=2.18 $Y2=1.515
r29 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.18 $Y=1.665
+ $X2=2.18 $Y2=1.515
r30 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.105 $Y=1.765
+ $X2=2.18 $Y2=1.515
r31 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.105 $Y=1.765
+ $X2=2.105 $Y2=2.34
r32 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.09 $Y=1.35
+ $X2=2.18 $Y2=1.515
r33 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.09 $Y=1.35 $X2=2.09
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A32O_2%A1 3 5 7 8 12
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.75
+ $Y=1.515 $X2=2.75 $Y2=1.515
r32 8 12 4.43247 $w=3.88e-07 $l=1.5e-07 $layer=LI1_cond $X=2.72 $Y=1.665
+ $X2=2.72 $Y2=1.515
r33 5 11 52.2586 $w=2.99e-07 $l=2.80624e-07 $layer=POLY_cond $X=2.815 $Y=1.765
+ $X2=2.75 $Y2=1.515
r34 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.815 $Y=1.765
+ $X2=2.815 $Y2=2.34
r35 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.66 $Y=1.35
+ $X2=2.75 $Y2=1.515
r36 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.66 $Y=1.35 $X2=2.66
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A32O_2%B1 3 5 7 8
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.32
+ $Y=1.515 $X2=3.32 $Y2=1.515
r32 8 12 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.32
+ $Y2=1.565
r33 5 11 52.2586 $w=2.99e-07 $l=2.76134e-07 $layer=POLY_cond $X=3.265 $Y=1.765
+ $X2=3.32 $Y2=1.515
r34 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.265 $Y=1.765
+ $X2=3.265 $Y2=2.34
r35 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.23 $Y=1.35
+ $X2=3.32 $Y2=1.515
r36 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.23 $Y=1.35 $X2=3.23
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A32O_2%B2 3 5 7 8 12
r21 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.465 $X2=4.05 $Y2=1.465
r22 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=4.05 $Y=1.665 $X2=4.05
+ $Y2=1.465
r23 5 11 55.8528 $w=4e-07 $l=3.69459e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.97 $Y2=1.465
r24 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=2.34
r25 1 11 39.5853 $w=4e-07 $l=2.38642e-07 $layer=POLY_cond $X=3.8 $Y=1.3 $X2=3.97
+ $Y2=1.465
r26 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.8 $Y=1.3 $X2=3.8
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A32O_2%VPWR 1 2 3 10 12 16 20 22 24 29 36 37 43 46
r55 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r57 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 37 47 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 34 46 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=2.455 $Y2=3.33
r61 34 36 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=4.08 $Y2=3.33
r62 30 43 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.51 $Y=3.33
+ $X2=1.305 $Y2=3.33
r63 30 32 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.51 $Y=3.33
+ $X2=2.16 $Y2=3.33
r64 29 46 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.265 $Y=3.33
+ $X2=2.455 $Y2=3.33
r65 29 32 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.265 $Y=3.33
+ $X2=2.16 $Y2=3.33
r66 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r67 28 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r68 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 25 40 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r70 25 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 24 43 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.1 $Y=3.33
+ $X2=1.305 $Y2=3.33
r72 24 27 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=0.72
+ $Y2=3.33
r73 22 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r74 22 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r75 22 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r76 18 46 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=3.245
+ $X2=2.455 $Y2=3.33
r77 18 20 16.0735 $w=3.78e-07 $l=5.3e-07 $layer=LI1_cond $X=2.455 $Y=3.245
+ $X2=2.455 $Y2=2.715
r78 14 43 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=3.245
+ $X2=1.305 $Y2=3.33
r79 14 16 11.8055 $w=4.08e-07 $l=4.2e-07 $layer=LI1_cond $X=1.305 $Y=3.245
+ $X2=1.305 $Y2=2.825
r80 10 40 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r81 10 12 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.78
r82 3 20 600 $w=1.7e-07 $l=1.0053e-06 $layer=licon1_PDIFF $count=1 $X=2.18
+ $Y=1.84 $X2=2.46 $Y2=2.715
r83 2 16 600 $w=1.7e-07 $l=1.11405e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.305 $Y2=2.825
r84 1 12 600 $w=1.7e-07 $l=1.0099e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_LS__A32O_2%X 1 2 9 13 14 18
c30 18 0 9.33911e-20 $X=0.75 $Y=1.82
c31 14 0 1.1265e-19 $X=0.72 $Y=2.035
c32 13 0 9.54331e-20 $X=0.775 $Y=1.15
r33 14 18 7.2765 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=1.985
+ $X2=0.75 $Y2=1.82
r34 13 18 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=0.83 $Y=1.15
+ $X2=0.83 $Y2=1.82
r35 7 13 7.12386 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=0.775 $Y=0.99
+ $X2=0.775 $Y2=1.15
r36 7 9 17.8269 $w=3.18e-07 $l=4.95e-07 $layer=LI1_cond $X=0.775 $Y=0.99
+ $X2=0.775 $Y2=0.495
r37 2 14 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r38 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.635
+ $Y=0.37 $X2=0.78 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LS__A32O_2%A_346_368# 1 2 3 12 14 15 16 17 20 23
c43 23 0 1.20518e-19 $X=1.88 $Y=2.375
r44 18 20 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=4.04 $Y=2.905
+ $X2=4.04 $Y2=2.065
r45 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.875 $Y=2.99
+ $X2=4.04 $Y2=2.905
r46 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.875 $Y=2.99
+ $X2=3.205 $Y2=2.99
r47 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.04 $Y=2.905
+ $X2=3.205 $Y2=2.99
r48 14 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=2.46 $X2=3.04
+ $Y2=2.375
r49 14 15 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.04 $Y=2.46
+ $X2=3.04 $Y2=2.905
r50 13 23 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=2.375
+ $X2=1.88 $Y2=2.375
r51 12 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=2.375
+ $X2=3.04 $Y2=2.375
r52 12 13 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.875 $Y=2.375
+ $X2=2.045 $Y2=2.375
r53 3 20 300 $w=1.7e-07 $l=2.90474e-07 $layer=licon1_PDIFF $count=2 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.065
r54 2 25 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=2.89
+ $Y=1.84 $X2=3.04 $Y2=2.375
r55 1 23 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=1.73
+ $Y=1.84 $X2=1.88 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LS__A32O_2%VGND 1 2 3 10 12 14 18 20 22 24 26 38 42
r42 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r43 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r45 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r46 33 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r47 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r48 30 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r49 29 32 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r50 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 27 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=0 $X2=1.35
+ $Y2=0
r52 27 29 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=0 $X2=1.68
+ $Y2=0
r53 26 41 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.85 $Y=0 $X2=4.085
+ $Y2=0
r54 26 32 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.85 $Y=0 $X2=3.6
+ $Y2=0
r55 24 33 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r56 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r57 20 41 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=4.015 $Y=0.085
+ $X2=4.085 $Y2=0
r58 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.015 $Y=0.085
+ $X2=4.015 $Y2=0.515
r59 16 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=0.085
+ $X2=1.35 $Y2=0
r60 16 18 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.35 $Y=0.085
+ $X2=1.35 $Y2=0.675
r61 15 35 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r62 14 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.35
+ $Y2=0
r63 14 15 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.185 $Y=0 $X2=0.445
+ $Y2=0
r64 10 35 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r65 10 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.515
r66 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.875
+ $Y=0.37 $X2=4.015 $Y2=0.515
r67 2 18 182 $w=1.7e-07 $l=4.20595e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.37 $X2=1.35 $Y2=0.675
r68 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

