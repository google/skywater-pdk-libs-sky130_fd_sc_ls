* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__maj3_2 A B C VGND VNB VPB VPWR X
X0 X a_87_264# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 VPWR A a_790_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_413_74# B a_87_264# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_793_74# C a_87_264# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 a_577_74# C VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 X a_87_264# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X6 VPWR A a_393_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_87_264# B a_577_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 VGND A a_413_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 a_393_368# B a_87_264# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_584_347# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND A a_793_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 VGND a_87_264# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 a_87_264# B a_584_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VPWR a_87_264# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X15 a_790_368# C a_87_264# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends
