* NGSPICE file created from sky130_fd_sc_ls__einvp_8.ext - technology: sky130A

.subckt sky130_fd_sc_ls__einvp_8 A TE VGND VNB VPB VPWR Z
M1000 a_27_368# A Z VPB phighvt w=1.12e+06u l=150000u
+  ad=3.0016e+12p pd=2.552e+07u as=1.344e+12p ps=1.136e+07u
M1001 a_27_368# a_802_323# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=1.6632e+12p ps=1.417e+07u
M1002 VPWR a_802_323# a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_368# A Z VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_74# TE VGND VNB nshort w=740000u l=150000u
+  ad=2.0276e+12p pd=1.88e+07u as=1.1433e+12p ps=1.049e+07u
M1005 a_27_74# A Z VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=9.842e+11p ps=8.58e+06u
M1006 VPWR a_802_323# a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_802_323# a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_368# a_802_323# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Z A a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Z A a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_368# a_802_323# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_74# TE VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR TE a_802_323# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.192e+11p ps=2.81e+06u
M1014 a_27_74# A Z VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND TE a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Z A a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_74# TE VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_368# A Z VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_802_323# a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_74# A Z VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Z A a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_368# A Z VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Z A a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_74# TE VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Z A a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Z A a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_27_74# A Z VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_27_368# a_802_323# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND TE a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND TE a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Z A a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND TE a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND TE a_802_323# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.146e+11p ps=2.06e+06u
.ends

