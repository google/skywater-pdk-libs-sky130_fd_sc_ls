* NGSPICE file created from sky130_fd_sc_ls__decaphe_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__decaphe_2 VGND VNB VPB VPWR
M1000 VPWR VGND VPWR VPB pshort w=1.255e+06u l=170000u
+  ad=6.526e+11p pd=6.06e+06u as=0p ps=0u
.ends

