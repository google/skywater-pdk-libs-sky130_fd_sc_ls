* NGSPICE file created from sky130_fd_sc_ls__a2bb2oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 Y a_114_392# a_539_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=2.296e+12p ps=1.978e+07u
M1001 a_539_368# B2 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=1.644e+12p ps=1.396e+07u
M1002 VGND a_114_392# Y VNB nshort w=740000u l=150000u
+  ad=1.2654e+12p pd=1.23e+07u as=8.288e+11p ps=8.16e+06u
M1003 Y a_114_392# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A1_N a_114_392# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1005 VPWR A1_N a_29_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=8.5e+11p ps=7.7e+06u
M1006 a_539_368# a_114_392# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B1 a_539_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B2 a_914_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=1.0138e+12p ps=1.014e+07u
M1009 VPWR B1 a_539_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B1 a_914_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_914_74# B2 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_914_74# B2 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_29_392# A1_N VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_114_392# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_539_368# B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR B2 a_539_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_539_368# B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_539_368# B2 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y a_114_392# a_539_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND B1 a_914_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR B2 a_539_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_114_392# A2_N VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y a_114_392# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_539_368# a_114_392# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_914_74# B1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_114_392# A2_N a_29_392# VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1027 a_29_392# A2_N a_114_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_914_74# B1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y B2 a_914_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

