* File: sky130_fd_sc_ls__o211a_4.pxi.spice
* Created: Wed Sep  2 11:17:26 2020
* 
x_PM_SKY130_FD_SC_LS__O211A_4%A_91_48# N_A_91_48#_M1013_s N_A_91_48#_M1003_d
+ N_A_91_48#_M1009_d N_A_91_48#_M1001_d N_A_91_48#_M1007_g N_A_91_48#_c_140_n
+ N_A_91_48#_M1008_g N_A_91_48#_M1015_g N_A_91_48#_c_141_n N_A_91_48#_M1012_g
+ N_A_91_48#_M1016_g N_A_91_48#_c_142_n N_A_91_48#_M1017_g N_A_91_48#_M1023_g
+ N_A_91_48#_c_143_n N_A_91_48#_M1022_g N_A_91_48#_c_134_n N_A_91_48#_c_135_n
+ N_A_91_48#_c_145_n N_A_91_48#_c_208_p N_A_91_48#_c_146_n N_A_91_48#_c_136_n
+ N_A_91_48#_c_137_n N_A_91_48#_c_148_n N_A_91_48#_c_149_n N_A_91_48#_c_138_n
+ N_A_91_48#_c_150_n N_A_91_48#_c_151_n N_A_91_48#_c_139_n
+ PM_SKY130_FD_SC_LS__O211A_4%A_91_48#
x_PM_SKY130_FD_SC_LS__O211A_4%C1 N_C1_c_309_n N_C1_M1004_g N_C1_M1013_g
+ N_C1_c_310_n N_C1_M1009_g N_C1_M1021_g C1 N_C1_c_308_n
+ PM_SKY130_FD_SC_LS__O211A_4%C1
x_PM_SKY130_FD_SC_LS__O211A_4%B1 N_B1_c_358_n N_B1_c_359_n N_B1_c_360_n
+ N_B1_c_366_n N_B1_M1003_g N_B1_c_361_n N_B1_M1011_g N_B1_c_362_n N_B1_c_368_n
+ N_B1_M1010_g N_B1_M1018_g N_B1_c_364_n B1 N_B1_c_365_n
+ PM_SKY130_FD_SC_LS__O211A_4%B1
x_PM_SKY130_FD_SC_LS__O211A_4%A2 N_A2_c_446_n N_A2_M1001_g N_A2_M1002_g
+ N_A2_c_447_n N_A2_M1005_g N_A2_M1019_g A2 A2 N_A2_c_444_n N_A2_c_445_n
+ PM_SKY130_FD_SC_LS__O211A_4%A2
x_PM_SKY130_FD_SC_LS__O211A_4%A1 N_A1_c_493_n N_A1_c_494_n N_A1_c_502_n
+ N_A1_M1000_g N_A1_M1006_g N_A1_c_496_n N_A1_c_497_n N_A1_c_498_n N_A1_M1014_g
+ N_A1_M1020_g A1 PM_SKY130_FD_SC_LS__O211A_4%A1
x_PM_SKY130_FD_SC_LS__O211A_4%VPWR N_VPWR_M1008_d N_VPWR_M1012_d N_VPWR_M1022_d
+ N_VPWR_M1004_s N_VPWR_M1010_s N_VPWR_M1014_s N_VPWR_c_559_n N_VPWR_c_560_n
+ N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_563_n N_VPWR_c_564_n N_VPWR_c_565_n
+ N_VPWR_c_566_n N_VPWR_c_567_n N_VPWR_c_568_n N_VPWR_c_569_n VPWR
+ N_VPWR_c_570_n N_VPWR_c_571_n N_VPWR_c_572_n N_VPWR_c_573_n N_VPWR_c_574_n
+ N_VPWR_c_575_n N_VPWR_c_558_n PM_SKY130_FD_SC_LS__O211A_4%VPWR
x_PM_SKY130_FD_SC_LS__O211A_4%X N_X_M1007_d N_X_M1016_d N_X_M1008_s N_X_M1017_s
+ N_X_c_651_n N_X_c_652_n N_X_c_658_n N_X_c_659_n N_X_c_653_n N_X_c_660_n
+ N_X_c_654_n N_X_c_661_n N_X_c_655_n N_X_c_662_n N_X_c_656_n N_X_c_663_n X X
+ PM_SKY130_FD_SC_LS__O211A_4%X
x_PM_SKY130_FD_SC_LS__O211A_4%A_968_391# N_A_968_391#_M1000_d
+ N_A_968_391#_M1005_s N_A_968_391#_c_734_n N_A_968_391#_c_730_n
+ N_A_968_391#_c_731_n N_A_968_391#_c_732_n
+ PM_SKY130_FD_SC_LS__O211A_4%A_968_391#
x_PM_SKY130_FD_SC_LS__O211A_4%VGND N_VGND_M1007_s N_VGND_M1015_s N_VGND_M1023_s
+ N_VGND_M1006_d N_VGND_M1019_s N_VGND_c_757_n N_VGND_c_758_n N_VGND_c_759_n
+ N_VGND_c_760_n N_VGND_c_761_n N_VGND_c_762_n VGND N_VGND_c_763_n
+ N_VGND_c_764_n N_VGND_c_765_n N_VGND_c_766_n N_VGND_c_767_n N_VGND_c_768_n
+ N_VGND_c_769_n N_VGND_c_770_n N_VGND_c_771_n N_VGND_c_772_n
+ PM_SKY130_FD_SC_LS__O211A_4%VGND
x_PM_SKY130_FD_SC_LS__O211A_4%A_510_125# N_A_510_125#_M1011_d
+ N_A_510_125#_M1018_d N_A_510_125#_M1002_d N_A_510_125#_M1020_s
+ N_A_510_125#_c_845_n N_A_510_125#_c_846_n N_A_510_125#_c_847_n
+ N_A_510_125#_c_848_n N_A_510_125#_c_849_n N_A_510_125#_c_850_n
+ N_A_510_125#_c_851_n N_A_510_125#_c_852_n N_A_510_125#_c_853_n
+ N_A_510_125#_c_854_n PM_SKY130_FD_SC_LS__O211A_4%A_510_125#
x_PM_SKY130_FD_SC_LS__O211A_4%A_597_125# N_A_597_125#_M1011_s
+ N_A_597_125#_M1021_d N_A_597_125#_c_917_n N_A_597_125#_c_918_n
+ N_A_597_125#_c_919_n N_A_597_125#_c_920_n
+ PM_SKY130_FD_SC_LS__O211A_4%A_597_125#
cc_1 VNB N_A_91_48#_M1007_g 0.0225008f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_2 VNB N_A_91_48#_M1015_g 0.0212087f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_3 VNB N_A_91_48#_M1016_g 0.0217869f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=0.74
cc_4 VNB N_A_91_48#_M1023_g 0.0216843f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=0.74
cc_5 VNB N_A_91_48#_c_134_n 0.00579892f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.465
cc_6 VNB N_A_91_48#_c_135_n 4.52924e-19 $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=1.95
cc_7 VNB N_A_91_48#_c_136_n 0.00167683f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=1.195
cc_8 VNB N_A_91_48#_c_137_n 0.00329567f $X=-0.19 $Y=-0.245 $X2=4.035 $Y2=1.95
cc_9 VNB N_A_91_48#_c_138_n 0.00248665f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.105
cc_10 VNB N_A_91_48#_c_139_n 0.111777f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=1.532
cc_11 VNB N_C1_M1013_g 0.0187808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C1_M1021_g 0.018993f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.3
cc_13 VNB C1 9.25683e-19 $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_14 VNB N_C1_c_308_n 0.0246865f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_15 VNB N_B1_c_358_n 0.0589691f $X=-0.19 $Y=-0.245 $X2=2.79 $Y2=1.955
cc_16 VNB N_B1_c_359_n 0.127671f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.955
cc_17 VNB N_B1_c_360_n 0.0123922f $X=-0.19 $Y=-0.245 $X2=5.29 $Y2=1.955
cc_18 VNB N_B1_c_361_n 0.0148688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_362_n 0.00923002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_M1018_g 0.0280602f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_21 VNB N_B1_c_364_n 0.0146186f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_22 VNB N_B1_c_365_n 0.041882f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=0.74
cc_23 VNB N_A2_M1002_g 0.0192298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A2_M1019_g 0.0195968f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.3
cc_25 VNB N_A2_c_444_n 0.00612267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_c_445_n 0.0261941f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.765
cc_27 VNB N_A1_c_493_n 0.0061924f $X=-0.19 $Y=-0.245 $X2=3.415 $Y2=0.625
cc_28 VNB N_A1_c_494_n 0.0141775f $X=-0.19 $Y=-0.245 $X2=2.79 $Y2=1.955
cc_29 VNB N_A1_M1006_g 0.0266069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A1_c_496_n 0.102837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A1_c_497_n 0.00990222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A1_c_498_n 0.0202328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A1_M1020_g 0.0458509f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_34 VNB A1 0.0115553f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.3
cc_35 VNB N_VPWR_c_558_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_651_n 0.00150518f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.3
cc_37 VNB N_X_c_652_n 0.00852127f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_38 VNB N_X_c_653_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_39 VNB N_X_c_654_n 0.00509139f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=1.3
cc_40 VNB N_X_c_655_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=2.4
cc_41 VNB N_X_c_656_n 0.00184578f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.465
cc_42 VNB X 0.0268466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_757_n 0.0117944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_758_n 0.0271311f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_45 VNB N_VGND_c_759_n 0.00495983f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_46 VNB N_VGND_c_760_n 0.0136768f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_47 VNB N_VGND_c_761_n 0.00381151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_762_n 0.0081779f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=1.3
cc_49 VNB N_VGND_c_763_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=1.765
cc_50 VNB N_VGND_c_764_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.465
cc_51 VNB N_VGND_c_765_n 0.0602851f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.465
cc_52 VNB N_VGND_c_766_n 0.0157641f $X=-0.19 $Y=-0.245 $X2=3.105 $Y2=2.035
cc_53 VNB N_VGND_c_767_n 0.0191172f $X=-0.19 $Y=-0.245 $X2=5.325 $Y2=2.035
cc_54 VNB N_VGND_c_768_n 0.351893f $X=-0.19 $Y=-0.245 $X2=4.12 $Y2=2.035
cc_55 VNB N_VGND_c_769_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.105
cc_56 VNB N_VGND_c_770_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_771_n 0.00459433f $X=-0.19 $Y=-0.245 $X2=5.49 $Y2=2.035
cc_58 VNB N_VGND_c_772_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.532
cc_59 VNB N_A_510_125#_c_845_n 0.0136664f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_60 VNB N_A_510_125#_c_846_n 0.0345039f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.765
cc_61 VNB N_A_510_125#_c_847_n 0.0029022f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_62 VNB N_A_510_125#_c_848_n 0.00395785f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_63 VNB N_A_510_125#_c_849_n 0.0042325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_510_125#_c_850_n 0.00458517f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=1.765
cc_65 VNB N_A_510_125#_c_851_n 0.00252813f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=1.3
cc_66 VNB N_A_510_125#_c_852_n 0.0152112f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=0.74
cc_67 VNB N_A_510_125#_c_853_n 0.0230853f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=2.4
cc_68 VNB N_A_510_125#_c_854_n 0.00182475f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=0.74
cc_69 VNB N_A_597_125#_c_917_n 0.00261948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_597_125#_c_918_n 0.00225846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_597_125#_c_919_n 0.0012438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_597_125#_c_920_n 0.00204411f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.3
cc_73 VPB N_A_91_48#_c_140_n 0.0164058f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=1.765
cc_74 VPB N_A_91_48#_c_141_n 0.0159595f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_75 VPB N_A_91_48#_c_142_n 0.0159587f $X=-0.19 $Y=1.66 $X2=1.555 $Y2=1.765
cc_76 VPB N_A_91_48#_c_143_n 0.0165444f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=1.765
cc_77 VPB N_A_91_48#_c_135_n 0.00314843f $X=-0.19 $Y=1.66 $X2=2.2 $Y2=1.95
cc_78 VPB N_A_91_48#_c_145_n 0.0023818f $X=-0.19 $Y=1.66 $X2=2.775 $Y2=2.035
cc_79 VPB N_A_91_48#_c_146_n 0.00565143f $X=-0.19 $Y=1.66 $X2=3.79 $Y2=2.035
cc_80 VPB N_A_91_48#_c_137_n 0.00227956f $X=-0.19 $Y=1.66 $X2=4.035 $Y2=1.95
cc_81 VPB N_A_91_48#_c_148_n 0.0111521f $X=-0.19 $Y=1.66 $X2=5.325 $Y2=2.035
cc_82 VPB N_A_91_48#_c_149_n 0.00884288f $X=-0.19 $Y=1.66 $X2=2.94 $Y2=2.115
cc_83 VPB N_A_91_48#_c_150_n 0.0053021f $X=-0.19 $Y=1.66 $X2=3.955 $Y2=2.115
cc_84 VPB N_A_91_48#_c_151_n 0.00193095f $X=-0.19 $Y=1.66 $X2=5.49 $Y2=2.115
cc_85 VPB N_A_91_48#_c_139_n 0.0270767f $X=-0.19 $Y=1.66 $X2=1.89 $Y2=1.532
cc_86 VPB N_C1_c_309_n 0.0158358f $X=-0.19 $Y=1.66 $X2=3.415 $Y2=0.625
cc_87 VPB N_C1_c_310_n 0.0158113f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_C1_c_308_n 0.0396796f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_89 VPB N_B1_c_366_n 0.0168307f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_B1_c_362_n 0.00704583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_B1_c_368_n 0.0215234f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1.3
cc_92 VPB B1 0.00163858f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_93 VPB N_B1_c_365_n 0.0270013f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=0.74
cc_94 VPB N_A2_c_446_n 0.0151193f $X=-0.19 $Y=1.66 $X2=3.415 $Y2=0.625
cc_95 VPB N_A2_c_447_n 0.0151968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A2_c_444_n 0.00407223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A2_c_445_n 0.0348612f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_98 VPB N_A1_c_494_n 0.00790997f $X=-0.19 $Y=1.66 $X2=2.79 $Y2=1.955
cc_99 VPB N_A1_c_502_n 0.0223404f $X=-0.19 $Y=1.66 $X2=3.805 $Y2=1.955
cc_100 VPB N_A1_c_498_n 0.0408078f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB A1 0.00733815f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.3
cc_102 VPB N_VPWR_c_559_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.4
cc_103 VPB N_VPWR_c_560_n 0.0441676f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_104 VPB N_VPWR_c_561_n 0.00830446f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_105 VPB N_VPWR_c_562_n 0.0186948f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=1.3
cc_106 VPB N_VPWR_c_563_n 0.0153207f $X=-0.19 $Y=1.66 $X2=1.555 $Y2=1.765
cc_107 VPB N_VPWR_c_564_n 0.0237932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_565_n 0.0155827f $X=-0.19 $Y=1.66 $X2=2.115 $Y2=1.465
cc_109 VPB N_VPWR_c_566_n 0.0121872f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_567_n 0.0540269f $X=-0.19 $Y=1.66 $X2=1.8 $Y2=1.465
cc_111 VPB N_VPWR_c_568_n 0.0244965f $X=-0.19 $Y=1.66 $X2=2.285 $Y2=2.035
cc_112 VPB N_VPWR_c_569_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_570_n 0.0186948f $X=-0.19 $Y=1.66 $X2=3.105 $Y2=2.035
cc_114 VPB N_VPWR_c_571_n 0.0209961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_572_n 0.0389417f $X=-0.19 $Y=1.66 $X2=3.555 $Y2=1.105
cc_116 VPB N_VPWR_c_573_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.532
cc_117 VPB N_VPWR_c_574_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.555 $Y2=1.532
cc_118 VPB N_VPWR_c_575_n 0.00631788f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=1.532
cc_119 VPB N_VPWR_c_558_n 0.0977646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_X_c_658_n 0.00173358f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_121 VPB N_X_c_659_n 0.00731501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_X_c_660_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_X_c_661_n 0.00427667f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=0.74
cc_124 VPB N_X_c_662_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_X_c_663_n 0.00183475f $X=-0.19 $Y=1.66 $X2=0.78 $Y2=1.465
cc_126 VPB X 0.00719016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_968_391#_c_730_n 0.00465845f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_968_391#_c_731_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_968_391#_c_732_n 0.00388828f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_130 N_A_91_48#_c_146_n N_C1_c_309_n 0.01419f $X=3.79 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_131 N_A_91_48#_c_149_n N_C1_c_309_n 0.0111444f $X=2.94 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_132 N_A_91_48#_c_150_n N_C1_c_309_n 8.74641e-19 $X=3.955 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_133 N_A_91_48#_c_138_n N_C1_M1013_g 0.00467806f $X=3.555 $Y=1.105 $X2=0 $Y2=0
cc_134 N_A_91_48#_c_146_n N_C1_c_310_n 0.0126656f $X=3.79 $Y=2.035 $X2=0 $Y2=0
cc_135 N_A_91_48#_c_137_n N_C1_c_310_n 0.0014866f $X=4.035 $Y=1.95 $X2=0 $Y2=0
cc_136 N_A_91_48#_c_149_n N_C1_c_310_n 8.66114e-19 $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_137 N_A_91_48#_c_150_n N_C1_c_310_n 0.011429f $X=3.955 $Y=2.115 $X2=0 $Y2=0
cc_138 N_A_91_48#_c_136_n N_C1_M1021_g 0.00999621f $X=3.95 $Y=1.195 $X2=0 $Y2=0
cc_139 N_A_91_48#_c_137_n N_C1_M1021_g 0.00848512f $X=4.035 $Y=1.95 $X2=0 $Y2=0
cc_140 N_A_91_48#_c_138_n N_C1_M1021_g 0.00505149f $X=3.555 $Y=1.105 $X2=0 $Y2=0
cc_141 N_A_91_48#_c_146_n C1 0.0243095f $X=3.79 $Y=2.035 $X2=0 $Y2=0
cc_142 N_A_91_48#_c_136_n C1 0.00423541f $X=3.95 $Y=1.195 $X2=0 $Y2=0
cc_143 N_A_91_48#_c_137_n C1 0.0247996f $X=4.035 $Y=1.95 $X2=0 $Y2=0
cc_144 N_A_91_48#_c_138_n C1 0.0213982f $X=3.555 $Y=1.105 $X2=0 $Y2=0
cc_145 N_A_91_48#_c_146_n N_C1_c_308_n 0.00815181f $X=3.79 $Y=2.035 $X2=0 $Y2=0
cc_146 N_A_91_48#_c_149_n N_C1_c_308_n 4.61094e-19 $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_147 N_A_91_48#_c_138_n N_C1_c_308_n 7.38938e-19 $X=3.555 $Y=1.105 $X2=0 $Y2=0
cc_148 N_A_91_48#_c_150_n N_C1_c_308_n 0.00155734f $X=3.955 $Y=2.115 $X2=0 $Y2=0
cc_149 N_A_91_48#_c_134_n N_B1_c_358_n 0.00639074f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_150 N_A_91_48#_c_139_n N_B1_c_358_n 0.0258648f $X=1.89 $Y=1.532 $X2=0 $Y2=0
cc_151 N_A_91_48#_M1023_g N_B1_c_360_n 0.0209604f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_91_48#_c_143_n N_B1_c_366_n 0.0140662f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A_91_48#_c_135_n N_B1_c_366_n 0.00128099f $X=2.2 $Y=1.95 $X2=0 $Y2=0
cc_154 N_A_91_48#_c_145_n N_B1_c_366_n 0.0128466f $X=2.775 $Y=2.035 $X2=0 $Y2=0
cc_155 N_A_91_48#_c_149_n N_B1_c_366_n 0.0135186f $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_156 N_A_91_48#_c_137_n N_B1_c_362_n 0.0077896f $X=4.035 $Y=1.95 $X2=0 $Y2=0
cc_157 N_A_91_48#_c_137_n N_B1_c_368_n 0.00453113f $X=4.035 $Y=1.95 $X2=0 $Y2=0
cc_158 N_A_91_48#_c_148_n N_B1_c_368_n 0.0172086f $X=5.325 $Y=2.035 $X2=0 $Y2=0
cc_159 N_A_91_48#_c_150_n N_B1_c_368_n 0.0113216f $X=3.955 $Y=2.115 $X2=0 $Y2=0
cc_160 N_A_91_48#_c_136_n N_B1_M1018_g 0.0016974f $X=3.95 $Y=1.195 $X2=0 $Y2=0
cc_161 N_A_91_48#_c_137_n N_B1_M1018_g 0.00136361f $X=4.035 $Y=1.95 $X2=0 $Y2=0
cc_162 N_A_91_48#_c_138_n N_B1_M1018_g 7.49792e-19 $X=3.555 $Y=1.105 $X2=0 $Y2=0
cc_163 N_A_91_48#_c_137_n N_B1_c_364_n 0.00452782f $X=4.035 $Y=1.95 $X2=0 $Y2=0
cc_164 N_A_91_48#_c_148_n N_B1_c_364_n 0.00229403f $X=5.325 $Y=2.035 $X2=0 $Y2=0
cc_165 N_A_91_48#_c_134_n B1 0.013554f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_166 N_A_91_48#_c_135_n B1 0.00932185f $X=2.2 $Y=1.95 $X2=0 $Y2=0
cc_167 N_A_91_48#_c_145_n B1 0.0203389f $X=2.775 $Y=2.035 $X2=0 $Y2=0
cc_168 N_A_91_48#_c_149_n B1 0.00506728f $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_169 N_A_91_48#_c_143_n N_B1_c_365_n 0.00158398f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A_91_48#_c_135_n N_B1_c_365_n 0.00307964f $X=2.2 $Y=1.95 $X2=0 $Y2=0
cc_171 N_A_91_48#_c_145_n N_B1_c_365_n 0.00860676f $X=2.775 $Y=2.035 $X2=0 $Y2=0
cc_172 N_A_91_48#_c_149_n N_B1_c_365_n 0.00602605f $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_173 N_A_91_48#_c_148_n N_A2_c_446_n 0.0150279f $X=5.325 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_174 N_A_91_48#_c_151_n N_A2_c_447_n 0.0091637f $X=5.49 $Y=2.115 $X2=0 $Y2=0
cc_175 N_A_91_48#_c_148_n N_A2_c_444_n 0.0302889f $X=5.325 $Y=2.035 $X2=0 $Y2=0
cc_176 N_A_91_48#_c_151_n N_A2_c_444_n 0.0277622f $X=5.49 $Y=2.115 $X2=0 $Y2=0
cc_177 N_A_91_48#_c_148_n N_A2_c_445_n 0.00132755f $X=5.325 $Y=2.035 $X2=0 $Y2=0
cc_178 N_A_91_48#_c_151_n N_A2_c_445_n 0.00802136f $X=5.49 $Y=2.115 $X2=0 $Y2=0
cc_179 N_A_91_48#_c_137_n N_A1_c_493_n 0.00238486f $X=4.035 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_180 N_A_91_48#_c_137_n N_A1_c_502_n 3.07613e-19 $X=4.035 $Y=1.95 $X2=0 $Y2=0
cc_181 N_A_91_48#_c_148_n N_A1_c_502_n 0.0186244f $X=5.325 $Y=2.035 $X2=0 $Y2=0
cc_182 N_A_91_48#_c_150_n N_A1_c_502_n 8.72518e-19 $X=3.955 $Y=2.115 $X2=0 $Y2=0
cc_183 N_A_91_48#_c_135_n N_VPWR_M1022_d 0.00235241f $X=2.2 $Y=1.95 $X2=0 $Y2=0
cc_184 N_A_91_48#_c_145_n N_VPWR_M1022_d 0.010294f $X=2.775 $Y=2.035 $X2=0 $Y2=0
cc_185 N_A_91_48#_c_208_p N_VPWR_M1022_d 0.00301935f $X=2.285 $Y=2.035 $X2=0
+ $Y2=0
cc_186 N_A_91_48#_c_146_n N_VPWR_M1004_s 0.00368373f $X=3.79 $Y=2.035 $X2=0
+ $Y2=0
cc_187 N_A_91_48#_c_148_n N_VPWR_M1010_s 0.00447846f $X=5.325 $Y=2.035 $X2=0
+ $Y2=0
cc_188 N_A_91_48#_c_140_n N_VPWR_c_560_n 0.0198182f $X=0.555 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_A_91_48#_c_141_n N_VPWR_c_561_n 0.00687925f $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_190 N_A_91_48#_c_142_n N_VPWR_c_561_n 0.00687925f $X=1.555 $Y=1.765 $X2=0
+ $Y2=0
cc_191 N_A_91_48#_c_142_n N_VPWR_c_562_n 0.00445602f $X=1.555 $Y=1.765 $X2=0
+ $Y2=0
cc_192 N_A_91_48#_c_143_n N_VPWR_c_562_n 0.00445602f $X=2.005 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_A_91_48#_c_143_n N_VPWR_c_563_n 0.00939425f $X=2.005 $Y=1.765 $X2=0
+ $Y2=0
cc_194 N_A_91_48#_c_145_n N_VPWR_c_563_n 0.0128995f $X=2.775 $Y=2.035 $X2=0
+ $Y2=0
cc_195 N_A_91_48#_c_208_p N_VPWR_c_563_n 0.0132989f $X=2.285 $Y=2.035 $X2=0
+ $Y2=0
cc_196 N_A_91_48#_c_149_n N_VPWR_c_563_n 0.0245375f $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_197 N_A_91_48#_c_146_n N_VPWR_c_564_n 0.0244889f $X=3.79 $Y=2.035 $X2=0 $Y2=0
cc_198 N_A_91_48#_c_149_n N_VPWR_c_564_n 0.0204897f $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_199 N_A_91_48#_c_150_n N_VPWR_c_564_n 0.0191531f $X=3.955 $Y=2.115 $X2=0
+ $Y2=0
cc_200 N_A_91_48#_c_148_n N_VPWR_c_565_n 0.0249771f $X=5.325 $Y=2.035 $X2=0
+ $Y2=0
cc_201 N_A_91_48#_c_150_n N_VPWR_c_565_n 0.0353168f $X=3.955 $Y=2.115 $X2=0
+ $Y2=0
cc_202 N_A_91_48#_c_149_n N_VPWR_c_568_n 0.00865944f $X=2.94 $Y=2.115 $X2=0
+ $Y2=0
cc_203 N_A_91_48#_c_140_n N_VPWR_c_570_n 0.00445602f $X=0.555 $Y=1.765 $X2=0
+ $Y2=0
cc_204 N_A_91_48#_c_141_n N_VPWR_c_570_n 0.00445602f $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_205 N_A_91_48#_c_150_n N_VPWR_c_571_n 0.00865944f $X=3.955 $Y=2.115 $X2=0
+ $Y2=0
cc_206 N_A_91_48#_c_140_n N_VPWR_c_558_n 0.00860566f $X=0.555 $Y=1.765 $X2=0
+ $Y2=0
cc_207 N_A_91_48#_c_141_n N_VPWR_c_558_n 0.00857797f $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_208 N_A_91_48#_c_142_n N_VPWR_c_558_n 0.00857797f $X=1.555 $Y=1.765 $X2=0
+ $Y2=0
cc_209 N_A_91_48#_c_143_n N_VPWR_c_558_n 0.00861719f $X=2.005 $Y=1.765 $X2=0
+ $Y2=0
cc_210 N_A_91_48#_c_149_n N_VPWR_c_558_n 0.0108276f $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_211 N_A_91_48#_c_150_n N_VPWR_c_558_n 0.0108276f $X=3.955 $Y=2.115 $X2=0
+ $Y2=0
cc_212 N_A_91_48#_M1007_g N_X_c_651_n 0.0143589f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A_91_48#_c_140_n N_X_c_658_n 0.0153702f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_214 N_A_91_48#_c_139_n N_X_c_658_n 8.08947e-19 $X=1.89 $Y=1.532 $X2=0 $Y2=0
cc_215 N_A_91_48#_M1007_g N_X_c_653_n 0.0128625f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A_91_48#_M1015_g N_X_c_653_n 3.97481e-19 $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A_91_48#_c_140_n N_X_c_660_n 0.0165744f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A_91_48#_c_141_n N_X_c_660_n 0.0123916f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A_91_48#_c_142_n N_X_c_660_n 6.94077e-19 $X=1.555 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A_91_48#_M1015_g N_X_c_654_n 0.0128832f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_91_48#_M1016_g N_X_c_654_n 0.0124641f $X=1.46 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A_91_48#_c_134_n N_X_c_654_n 0.0709823f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_223 N_A_91_48#_c_139_n N_X_c_654_n 0.0061855f $X=1.89 $Y=1.532 $X2=0 $Y2=0
cc_224 N_A_91_48#_c_141_n N_X_c_661_n 0.0125195f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_225 N_A_91_48#_c_142_n N_X_c_661_n 0.0134585f $X=1.555 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A_91_48#_c_143_n N_X_c_661_n 0.00237275f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A_91_48#_c_134_n N_X_c_661_n 0.0769703f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_228 N_A_91_48#_c_135_n N_X_c_661_n 0.00779207f $X=2.2 $Y=1.95 $X2=0 $Y2=0
cc_229 N_A_91_48#_c_139_n N_X_c_661_n 0.017972f $X=1.89 $Y=1.532 $X2=0 $Y2=0
cc_230 N_A_91_48#_M1015_g N_X_c_655_n 9.31498e-19 $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A_91_48#_M1016_g N_X_c_655_n 0.00862472f $X=1.46 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A_91_48#_M1023_g N_X_c_655_n 3.97481e-19 $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A_91_48#_c_141_n N_X_c_662_n 6.94077e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A_91_48#_c_142_n N_X_c_662_n 0.0123916f $X=1.555 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A_91_48#_c_143_n N_X_c_662_n 0.0129054f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_236 N_A_91_48#_M1007_g N_X_c_656_n 0.00132316f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A_91_48#_c_134_n N_X_c_656_n 0.0181339f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_238 N_A_91_48#_c_139_n N_X_c_656_n 0.00232957f $X=1.89 $Y=1.532 $X2=0 $Y2=0
cc_239 N_A_91_48#_c_140_n N_X_c_663_n 9.3899e-19 $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_240 N_A_91_48#_c_141_n N_X_c_663_n 9.3899e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A_91_48#_c_134_n N_X_c_663_n 0.0276943f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_242 N_A_91_48#_c_139_n N_X_c_663_n 0.00792231f $X=1.89 $Y=1.532 $X2=0 $Y2=0
cc_243 N_A_91_48#_M1007_g X 0.0109941f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_91_48#_c_140_n X 0.00126693f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_245 N_A_91_48#_c_134_n X 0.0194533f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_246 N_A_91_48#_c_139_n X 0.0105753f $X=1.89 $Y=1.532 $X2=0 $Y2=0
cc_247 N_A_91_48#_c_148_n N_A_968_391#_M1000_d 0.00197722f $X=5.325 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_248 N_A_91_48#_c_148_n N_A_968_391#_c_734_n 0.0171814f $X=5.325 $Y=2.035
+ $X2=0 $Y2=0
cc_249 N_A_91_48#_M1001_d N_A_968_391#_c_730_n 0.00250873f $X=5.29 $Y=1.955
+ $X2=0 $Y2=0
cc_250 N_A_91_48#_c_151_n N_A_968_391#_c_730_n 0.018923f $X=5.49 $Y=2.115 $X2=0
+ $Y2=0
cc_251 N_A_91_48#_c_151_n N_A_968_391#_c_732_n 0.0533133f $X=5.49 $Y=2.115 $X2=0
+ $Y2=0
cc_252 N_A_91_48#_M1007_g N_VGND_c_758_n 0.00409307f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_91_48#_M1007_g N_VGND_c_759_n 5.04273e-19 $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_91_48#_M1015_g N_VGND_c_759_n 0.00935695f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_91_48#_M1016_g N_VGND_c_759_n 0.00397833f $X=1.46 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A_91_48#_M1016_g N_VGND_c_760_n 6.13182e-19 $X=1.46 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A_91_48#_M1023_g N_VGND_c_760_n 0.013465f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A_91_48#_c_134_n N_VGND_c_760_n 0.029036f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_259 N_A_91_48#_c_139_n N_VGND_c_760_n 0.00350673f $X=1.89 $Y=1.532 $X2=0
+ $Y2=0
cc_260 N_A_91_48#_M1007_g N_VGND_c_763_n 0.00434272f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_91_48#_M1015_g N_VGND_c_763_n 0.00383152f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_91_48#_M1016_g N_VGND_c_764_n 0.00434272f $X=1.46 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_91_48#_M1023_g N_VGND_c_764_n 0.00383152f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A_91_48#_M1007_g N_VGND_c_768_n 0.00824056f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A_91_48#_M1015_g N_VGND_c_768_n 0.0075754f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_266 N_A_91_48#_M1016_g N_VGND_c_768_n 0.00820718f $X=1.46 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A_91_48#_M1023_g N_VGND_c_768_n 0.0075754f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A_91_48#_M1023_g N_A_510_125#_c_845_n 4.67658e-19 $X=1.89 $Y=0.74 $X2=0
+ $Y2=0
cc_269 N_A_91_48#_M1023_g N_A_510_125#_c_847_n 2.4306e-19 $X=1.89 $Y=0.74 $X2=0
+ $Y2=0
cc_270 N_A_91_48#_c_148_n N_A_510_125#_c_849_n 0.006809f $X=5.325 $Y=2.035 $X2=0
+ $Y2=0
cc_271 N_A_91_48#_c_136_n N_A_510_125#_c_850_n 0.00537821f $X=3.95 $Y=1.195
+ $X2=0 $Y2=0
cc_272 N_A_91_48#_c_137_n N_A_510_125#_c_850_n 2.47868e-19 $X=4.035 $Y=1.95
+ $X2=0 $Y2=0
cc_273 N_A_91_48#_c_148_n N_A_510_125#_c_850_n 0.00812137f $X=5.325 $Y=2.035
+ $X2=0 $Y2=0
cc_274 N_A_91_48#_c_136_n N_A_597_125#_M1021_d 0.0041638f $X=3.95 $Y=1.195 $X2=0
+ $Y2=0
cc_275 N_A_91_48#_c_146_n N_A_597_125#_c_917_n 0.00298145f $X=3.79 $Y=2.035
+ $X2=0 $Y2=0
cc_276 N_A_91_48#_c_149_n N_A_597_125#_c_917_n 0.00222656f $X=2.94 $Y=2.115
+ $X2=0 $Y2=0
cc_277 N_A_91_48#_c_138_n N_A_597_125#_c_917_n 0.0128711f $X=3.555 $Y=1.105
+ $X2=0 $Y2=0
cc_278 N_A_91_48#_M1013_s N_A_597_125#_c_918_n 0.00169276f $X=3.415 $Y=0.625
+ $X2=0 $Y2=0
cc_279 N_A_91_48#_c_136_n N_A_597_125#_c_918_n 0.0048036f $X=3.95 $Y=1.195 $X2=0
+ $Y2=0
cc_280 N_A_91_48#_c_138_n N_A_597_125#_c_918_n 0.0161743f $X=3.555 $Y=1.105
+ $X2=0 $Y2=0
cc_281 N_A_91_48#_c_136_n N_A_597_125#_c_920_n 0.0182562f $X=3.95 $Y=1.195 $X2=0
+ $Y2=0
cc_282 N_C1_M1013_g N_B1_c_359_n 0.00737859f $X=3.34 $Y=0.945 $X2=0 $Y2=0
cc_283 N_C1_M1021_g N_B1_c_359_n 0.00737859f $X=3.77 $Y=0.945 $X2=0 $Y2=0
cc_284 N_C1_c_309_n N_B1_c_366_n 0.0146597f $X=3.165 $Y=1.88 $X2=0 $Y2=0
cc_285 N_C1_M1013_g N_B1_c_361_n 0.00877012f $X=3.34 $Y=0.945 $X2=0 $Y2=0
cc_286 N_C1_c_308_n N_B1_c_362_n 0.01402f $X=3.73 $Y=1.665 $X2=0 $Y2=0
cc_287 N_C1_c_310_n N_B1_c_368_n 0.0138176f $X=3.73 $Y=1.88 $X2=0 $Y2=0
cc_288 N_C1_M1021_g N_B1_M1018_g 0.0207562f $X=3.77 $Y=0.945 $X2=0 $Y2=0
cc_289 N_C1_M1021_g N_B1_c_364_n 0.01402f $X=3.77 $Y=0.945 $X2=0 $Y2=0
cc_290 C1 N_B1_c_364_n 2.95263e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_291 N_C1_M1013_g B1 0.00140466f $X=3.34 $Y=0.945 $X2=0 $Y2=0
cc_292 C1 B1 0.00858387f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_293 N_C1_c_308_n B1 3.40608e-19 $X=3.73 $Y=1.665 $X2=0 $Y2=0
cc_294 C1 N_B1_c_365_n 0.00107002f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_295 N_C1_c_308_n N_B1_c_365_n 0.0246125f $X=3.73 $Y=1.665 $X2=0 $Y2=0
cc_296 N_C1_c_309_n N_VPWR_c_564_n 0.00653597f $X=3.165 $Y=1.88 $X2=0 $Y2=0
cc_297 N_C1_c_310_n N_VPWR_c_564_n 0.00638017f $X=3.73 $Y=1.88 $X2=0 $Y2=0
cc_298 N_C1_c_309_n N_VPWR_c_568_n 0.00455131f $X=3.165 $Y=1.88 $X2=0 $Y2=0
cc_299 N_C1_c_310_n N_VPWR_c_571_n 0.00455131f $X=3.73 $Y=1.88 $X2=0 $Y2=0
cc_300 N_C1_c_309_n N_VPWR_c_558_n 0.00495025f $X=3.165 $Y=1.88 $X2=0 $Y2=0
cc_301 N_C1_c_310_n N_VPWR_c_558_n 0.00495025f $X=3.73 $Y=1.88 $X2=0 $Y2=0
cc_302 N_C1_M1013_g N_A_510_125#_c_846_n 0.00116683f $X=3.34 $Y=0.945 $X2=0
+ $Y2=0
cc_303 N_C1_M1021_g N_A_510_125#_c_846_n 0.00116683f $X=3.77 $Y=0.945 $X2=0
+ $Y2=0
cc_304 N_C1_M1013_g N_A_597_125#_c_917_n 2.23441e-19 $X=3.34 $Y=0.945 $X2=0
+ $Y2=0
cc_305 N_C1_c_308_n N_A_597_125#_c_917_n 0.00315705f $X=3.73 $Y=1.665 $X2=0
+ $Y2=0
cc_306 N_C1_M1013_g N_A_597_125#_c_918_n 0.0114956f $X=3.34 $Y=0.945 $X2=0 $Y2=0
cc_307 N_C1_M1021_g N_A_597_125#_c_918_n 0.00923977f $X=3.77 $Y=0.945 $X2=0
+ $Y2=0
cc_308 N_C1_M1021_g N_A_597_125#_c_920_n 4.44855e-19 $X=3.77 $Y=0.945 $X2=0
+ $Y2=0
cc_309 N_B1_c_364_n N_A1_c_493_n 0.00605855f $X=4.217 $Y=1.49 $X2=-0.19
+ $Y2=-0.245
cc_310 N_B1_c_362_n N_A1_c_494_n 0.00564817f $X=4.18 $Y=1.79 $X2=0 $Y2=0
cc_311 N_B1_c_368_n N_A1_c_502_n 0.0281668f $X=4.18 $Y=1.88 $X2=0 $Y2=0
cc_312 N_B1_M1018_g N_A1_M1006_g 0.0132251f $X=4.27 $Y=0.945 $X2=0 $Y2=0
cc_313 N_B1_c_359_n N_A1_c_497_n 0.0132251f $X=4.195 $Y=0.18 $X2=0 $Y2=0
cc_314 N_B1_c_366_n N_VPWR_c_563_n 0.00813486f $X=2.715 $Y=1.88 $X2=0 $Y2=0
cc_315 N_B1_c_368_n N_VPWR_c_565_n 0.0082054f $X=4.18 $Y=1.88 $X2=0 $Y2=0
cc_316 N_B1_c_366_n N_VPWR_c_568_n 0.00455131f $X=2.715 $Y=1.88 $X2=0 $Y2=0
cc_317 N_B1_c_368_n N_VPWR_c_571_n 0.00455131f $X=4.18 $Y=1.88 $X2=0 $Y2=0
cc_318 N_B1_c_366_n N_VPWR_c_558_n 0.00495025f $X=2.715 $Y=1.88 $X2=0 $Y2=0
cc_319 N_B1_c_368_n N_VPWR_c_558_n 0.00495025f $X=4.18 $Y=1.88 $X2=0 $Y2=0
cc_320 N_B1_c_366_n N_X_c_662_n 8.83558e-19 $X=2.715 $Y=1.88 $X2=0 $Y2=0
cc_321 N_B1_c_360_n N_VGND_c_760_n 0.0144891f $X=2.475 $Y=0.18 $X2=0 $Y2=0
cc_322 N_B1_c_359_n N_VGND_c_761_n 0.00107466f $X=4.195 $Y=0.18 $X2=0 $Y2=0
cc_323 N_B1_M1018_g N_VGND_c_761_n 2.44756e-19 $X=4.27 $Y=0.945 $X2=0 $Y2=0
cc_324 N_B1_c_360_n N_VGND_c_765_n 0.045518f $X=2.475 $Y=0.18 $X2=0 $Y2=0
cc_325 N_B1_c_359_n N_VGND_c_768_n 0.047086f $X=4.195 $Y=0.18 $X2=0 $Y2=0
cc_326 N_B1_c_360_n N_VGND_c_768_n 0.0114395f $X=2.475 $Y=0.18 $X2=0 $Y2=0
cc_327 N_B1_c_358_n N_A_510_125#_c_845_n 0.0110018f $X=2.4 $Y=1.34 $X2=0 $Y2=0
cc_328 N_B1_c_361_n N_A_510_125#_c_845_n 0.00295702f $X=2.91 $Y=1.34 $X2=0 $Y2=0
cc_329 B1 N_A_510_125#_c_845_n 0.0206962f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_330 N_B1_c_365_n N_A_510_125#_c_845_n 0.00528389f $X=2.715 $Y=1.61 $X2=0
+ $Y2=0
cc_331 N_B1_c_359_n N_A_510_125#_c_846_n 0.023808f $X=4.195 $Y=0.18 $X2=0 $Y2=0
cc_332 N_B1_c_361_n N_A_510_125#_c_846_n 0.00366331f $X=2.91 $Y=1.34 $X2=0 $Y2=0
cc_333 N_B1_M1018_g N_A_510_125#_c_846_n 0.0156653f $X=4.27 $Y=0.945 $X2=0 $Y2=0
cc_334 N_B1_c_358_n N_A_510_125#_c_847_n 0.00198754f $X=2.4 $Y=1.34 $X2=0 $Y2=0
cc_335 N_B1_c_359_n N_A_510_125#_c_847_n 0.00732085f $X=4.195 $Y=0.18 $X2=0
+ $Y2=0
cc_336 N_B1_M1018_g N_A_510_125#_c_848_n 0.0047697f $X=4.27 $Y=0.945 $X2=0 $Y2=0
cc_337 N_B1_M1018_g N_A_510_125#_c_850_n 2.13054e-19 $X=4.27 $Y=0.945 $X2=0
+ $Y2=0
cc_338 N_B1_c_361_n N_A_597_125#_c_917_n 4.5765e-19 $X=2.91 $Y=1.34 $X2=0 $Y2=0
cc_339 N_B1_c_361_n N_A_597_125#_c_919_n 2.90897e-19 $X=2.91 $Y=1.34 $X2=0 $Y2=0
cc_340 N_B1_M1018_g N_A_597_125#_c_920_n 0.00538803f $X=4.27 $Y=0.945 $X2=0
+ $Y2=0
cc_341 N_B1_c_364_n N_A_597_125#_c_920_n 0.00185803f $X=4.217 $Y=1.49 $X2=0
+ $Y2=0
cc_342 N_A2_c_445_n N_A1_c_493_n 0.0157564f $X=5.715 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_343 N_A2_c_444_n N_A1_c_494_n 0.0102979f $X=5.67 $Y=1.615 $X2=0 $Y2=0
cc_344 N_A2_c_445_n N_A1_c_494_n 0.0118237f $X=5.715 $Y=1.665 $X2=0 $Y2=0
cc_345 N_A2_c_446_n N_A1_c_502_n 0.0201905f $X=5.215 $Y=1.88 $X2=0 $Y2=0
cc_346 N_A2_M1002_g N_A1_M1006_g 0.0157564f $X=5.24 $Y=0.945 $X2=0 $Y2=0
cc_347 N_A2_M1002_g N_A1_c_496_n 0.00902758f $X=5.24 $Y=0.945 $X2=0 $Y2=0
cc_348 N_A2_M1019_g N_A1_c_496_n 0.00894529f $X=5.725 $Y=0.945 $X2=0 $Y2=0
cc_349 N_A2_c_447_n N_A1_c_498_n 0.0088506f $X=5.715 $Y=1.88 $X2=0 $Y2=0
cc_350 N_A2_c_444_n N_A1_c_498_n 4.16072e-19 $X=5.67 $Y=1.615 $X2=0 $Y2=0
cc_351 N_A2_c_445_n N_A1_c_498_n 0.0236458f $X=5.715 $Y=1.665 $X2=0 $Y2=0
cc_352 N_A2_M1019_g N_A1_M1020_g 0.0255078f $X=5.725 $Y=0.945 $X2=0 $Y2=0
cc_353 N_A2_c_444_n A1 0.0205984f $X=5.67 $Y=1.615 $X2=0 $Y2=0
cc_354 N_A2_c_445_n A1 4.1393e-19 $X=5.715 $Y=1.665 $X2=0 $Y2=0
cc_355 N_A2_c_446_n N_VPWR_c_572_n 0.00275693f $X=5.215 $Y=1.88 $X2=0 $Y2=0
cc_356 N_A2_c_447_n N_VPWR_c_572_n 0.00275707f $X=5.715 $Y=1.88 $X2=0 $Y2=0
cc_357 N_A2_c_446_n N_VPWR_c_558_n 0.00544287f $X=5.215 $Y=1.88 $X2=0 $Y2=0
cc_358 N_A2_c_447_n N_VPWR_c_558_n 0.00544287f $X=5.715 $Y=1.88 $X2=0 $Y2=0
cc_359 N_A2_c_446_n N_A_968_391#_c_734_n 0.00769156f $X=5.215 $Y=1.88 $X2=0
+ $Y2=0
cc_360 N_A2_c_447_n N_A_968_391#_c_734_n 8.49836e-19 $X=5.715 $Y=1.88 $X2=0
+ $Y2=0
cc_361 N_A2_c_446_n N_A_968_391#_c_730_n 0.0110936f $X=5.215 $Y=1.88 $X2=0 $Y2=0
cc_362 N_A2_c_447_n N_A_968_391#_c_730_n 0.0131124f $X=5.715 $Y=1.88 $X2=0 $Y2=0
cc_363 N_A2_c_446_n N_A_968_391#_c_731_n 0.00177718f $X=5.215 $Y=1.88 $X2=0
+ $Y2=0
cc_364 N_A2_c_447_n N_A_968_391#_c_732_n 0.00631643f $X=5.715 $Y=1.88 $X2=0
+ $Y2=0
cc_365 N_A2_M1002_g N_VGND_c_761_n 0.00684563f $X=5.24 $Y=0.945 $X2=0 $Y2=0
cc_366 N_A2_M1019_g N_VGND_c_761_n 4.05518e-19 $X=5.725 $Y=0.945 $X2=0 $Y2=0
cc_367 N_A2_M1002_g N_VGND_c_762_n 4.23833e-19 $X=5.24 $Y=0.945 $X2=0 $Y2=0
cc_368 N_A2_M1019_g N_VGND_c_762_n 0.00771226f $X=5.725 $Y=0.945 $X2=0 $Y2=0
cc_369 N_A2_M1002_g N_VGND_c_768_n 8.92987e-19 $X=5.24 $Y=0.945 $X2=0 $Y2=0
cc_370 N_A2_M1019_g N_VGND_c_768_n 7.97988e-19 $X=5.725 $Y=0.945 $X2=0 $Y2=0
cc_371 N_A2_M1002_g N_A_510_125#_c_849_n 0.0128053f $X=5.24 $Y=0.945 $X2=0 $Y2=0
cc_372 N_A2_c_444_n N_A_510_125#_c_849_n 0.0319578f $X=5.67 $Y=1.615 $X2=0 $Y2=0
cc_373 N_A2_M1019_g N_A_510_125#_c_852_n 0.0125779f $X=5.725 $Y=0.945 $X2=0
+ $Y2=0
cc_374 N_A2_c_444_n N_A_510_125#_c_852_n 0.0174392f $X=5.67 $Y=1.615 $X2=0 $Y2=0
cc_375 N_A2_c_445_n N_A_510_125#_c_852_n 7.91014e-19 $X=5.715 $Y=1.665 $X2=0
+ $Y2=0
cc_376 N_A2_M1019_g N_A_510_125#_c_853_n 8.30676e-19 $X=5.725 $Y=0.945 $X2=0
+ $Y2=0
cc_377 N_A2_c_444_n N_A_510_125#_c_854_n 0.0210724f $X=5.67 $Y=1.615 $X2=0 $Y2=0
cc_378 N_A2_c_445_n N_A_510_125#_c_854_n 0.00360392f $X=5.715 $Y=1.665 $X2=0
+ $Y2=0
cc_379 N_A1_c_502_n N_VPWR_c_565_n 0.00781719f $X=4.765 $Y=1.88 $X2=0 $Y2=0
cc_380 N_A1_c_498_n N_VPWR_c_567_n 0.0259727f $X=6.165 $Y=1.88 $X2=0 $Y2=0
cc_381 A1 N_VPWR_c_567_n 0.0276867f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_382 N_A1_c_502_n N_VPWR_c_572_n 0.00439231f $X=4.765 $Y=1.88 $X2=0 $Y2=0
cc_383 N_A1_c_498_n N_VPWR_c_572_n 0.00439231f $X=6.165 $Y=1.88 $X2=0 $Y2=0
cc_384 N_A1_c_502_n N_VPWR_c_558_n 0.00544287f $X=4.765 $Y=1.88 $X2=0 $Y2=0
cc_385 N_A1_c_498_n N_VPWR_c_558_n 0.00544287f $X=6.165 $Y=1.88 $X2=0 $Y2=0
cc_386 N_A1_c_502_n N_A_968_391#_c_734_n 0.00623494f $X=4.765 $Y=1.88 $X2=0
+ $Y2=0
cc_387 N_A1_c_498_n N_A_968_391#_c_730_n 0.00324945f $X=6.165 $Y=1.88 $X2=0
+ $Y2=0
cc_388 N_A1_c_502_n N_A_968_391#_c_731_n 0.00324789f $X=4.765 $Y=1.88 $X2=0
+ $Y2=0
cc_389 N_A1_c_498_n N_A_968_391#_c_732_n 0.0101243f $X=6.165 $Y=1.88 $X2=0 $Y2=0
cc_390 A1 N_A_968_391#_c_732_n 0.00238238f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_391 N_A1_M1006_g N_VGND_c_761_n 0.0139844f $X=4.78 $Y=0.945 $X2=0 $Y2=0
cc_392 N_A1_c_496_n N_VGND_c_761_n 0.0185436f $X=6.15 $Y=0.18 $X2=0 $Y2=0
cc_393 N_A1_c_497_n N_VGND_c_761_n 0.00364942f $X=4.855 $Y=0.18 $X2=0 $Y2=0
cc_394 N_A1_c_496_n N_VGND_c_762_n 0.0232456f $X=6.15 $Y=0.18 $X2=0 $Y2=0
cc_395 N_A1_M1020_g N_VGND_c_762_n 0.0151144f $X=6.225 $Y=0.945 $X2=0 $Y2=0
cc_396 N_A1_c_497_n N_VGND_c_765_n 0.00486043f $X=4.855 $Y=0.18 $X2=0 $Y2=0
cc_397 N_A1_c_496_n N_VGND_c_766_n 0.0184168f $X=6.15 $Y=0.18 $X2=0 $Y2=0
cc_398 N_A1_c_496_n N_VGND_c_767_n 0.00730708f $X=6.15 $Y=0.18 $X2=0 $Y2=0
cc_399 N_A1_c_496_n N_VGND_c_768_n 0.0323021f $X=6.15 $Y=0.18 $X2=0 $Y2=0
cc_400 N_A1_c_497_n N_VGND_c_768_n 0.00859636f $X=4.855 $Y=0.18 $X2=0 $Y2=0
cc_401 N_A1_M1006_g N_A_510_125#_c_846_n 0.00157748f $X=4.78 $Y=0.945 $X2=0
+ $Y2=0
cc_402 N_A1_M1006_g N_A_510_125#_c_848_n 0.00421702f $X=4.78 $Y=0.945 $X2=0
+ $Y2=0
cc_403 N_A1_c_493_n N_A_510_125#_c_849_n 0.00105349f $X=4.765 $Y=1.43 $X2=0
+ $Y2=0
cc_404 N_A1_M1006_g N_A_510_125#_c_849_n 0.0167614f $X=4.78 $Y=0.945 $X2=0 $Y2=0
cc_405 N_A1_c_496_n N_A_510_125#_c_851_n 0.00490132f $X=6.15 $Y=0.18 $X2=0 $Y2=0
cc_406 N_A1_c_498_n N_A_510_125#_c_852_n 0.00437819f $X=6.165 $Y=1.88 $X2=0
+ $Y2=0
cc_407 N_A1_M1020_g N_A_510_125#_c_852_n 0.0124988f $X=6.225 $Y=0.945 $X2=0
+ $Y2=0
cc_408 A1 N_A_510_125#_c_852_n 0.0421713f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_409 N_A1_M1020_g N_A_510_125#_c_853_n 0.00759673f $X=6.225 $Y=0.945 $X2=0
+ $Y2=0
cc_410 N_VPWR_M1008_d N_X_c_658_n 7.12223e-19 $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_411 N_VPWR_c_560_n N_X_c_658_n 0.00549591f $X=0.28 $Y=2.305 $X2=0 $Y2=0
cc_412 N_VPWR_M1008_d N_X_c_659_n 0.00362184f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_413 N_VPWR_c_560_n N_X_c_659_n 0.0207257f $X=0.28 $Y=2.305 $X2=0 $Y2=0
cc_414 N_VPWR_c_560_n N_X_c_660_n 0.0323093f $X=0.28 $Y=2.305 $X2=0 $Y2=0
cc_415 N_VPWR_c_561_n N_X_c_660_n 0.0323093f $X=1.28 $Y=2.305 $X2=0 $Y2=0
cc_416 N_VPWR_c_570_n N_X_c_660_n 0.014552f $X=1.115 $Y=3.33 $X2=0 $Y2=0
cc_417 N_VPWR_c_558_n N_X_c_660_n 0.0119791f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_418 N_VPWR_M1012_d N_X_c_661_n 0.00332584f $X=1.08 $Y=1.84 $X2=0 $Y2=0
cc_419 N_VPWR_c_561_n N_X_c_661_n 0.0232685f $X=1.28 $Y=2.305 $X2=0 $Y2=0
cc_420 N_VPWR_c_561_n N_X_c_662_n 0.0323093f $X=1.28 $Y=2.305 $X2=0 $Y2=0
cc_421 N_VPWR_c_562_n N_X_c_662_n 0.014552f $X=2.115 $Y=3.33 $X2=0 $Y2=0
cc_422 N_VPWR_c_563_n N_X_c_662_n 0.0266809f $X=2.28 $Y=2.405 $X2=0 $Y2=0
cc_423 N_VPWR_c_558_n N_X_c_662_n 0.0119791f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_424 N_VPWR_c_567_n N_A_968_391#_c_730_n 0.0121328f $X=6.44 $Y=2.115 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_572_n N_A_968_391#_c_730_n 0.0620441f $X=6.275 $Y=3.33 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_558_n N_A_968_391#_c_730_n 0.0346602f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_565_n N_A_968_391#_c_731_n 0.0121328f $X=4.49 $Y=2.41 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_572_n N_A_968_391#_c_731_n 0.0235512f $X=6.275 $Y=3.33 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_558_n N_A_968_391#_c_731_n 0.0126924f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_567_n N_A_968_391#_c_732_n 0.0344717f $X=6.44 $Y=2.115 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_567_n N_A_510_125#_c_852_n 3.21367e-19 $X=6.44 $Y=2.115 $X2=0
+ $Y2=0
cc_432 N_X_c_651_n N_VGND_M1007_s 4.46468e-19 $X=0.58 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_433 N_X_c_652_n N_VGND_M1007_s 0.00291902f $X=0.355 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_434 N_X_c_654_n N_VGND_M1015_s 0.00250873f $X=1.51 $Y=1.045 $X2=0 $Y2=0
cc_435 N_X_c_651_n N_VGND_c_758_n 0.00346194f $X=0.58 $Y=1.045 $X2=0 $Y2=0
cc_436 N_X_c_652_n N_VGND_c_758_n 0.0184602f $X=0.355 $Y=1.045 $X2=0 $Y2=0
cc_437 N_X_c_653_n N_VGND_c_758_n 0.0158413f $X=0.745 $Y=0.515 $X2=0 $Y2=0
cc_438 N_X_c_653_n N_VGND_c_759_n 0.0164981f $X=0.745 $Y=0.515 $X2=0 $Y2=0
cc_439 N_X_c_654_n N_VGND_c_759_n 0.0210288f $X=1.51 $Y=1.045 $X2=0 $Y2=0
cc_440 N_X_c_655_n N_VGND_c_759_n 0.0166127f $X=1.675 $Y=0.515 $X2=0 $Y2=0
cc_441 N_X_c_654_n N_VGND_c_760_n 0.00697079f $X=1.51 $Y=1.045 $X2=0 $Y2=0
cc_442 N_X_c_655_n N_VGND_c_760_n 0.0225912f $X=1.675 $Y=0.515 $X2=0 $Y2=0
cc_443 N_X_c_653_n N_VGND_c_763_n 0.0109942f $X=0.745 $Y=0.515 $X2=0 $Y2=0
cc_444 N_X_c_655_n N_VGND_c_764_n 0.0109942f $X=1.675 $Y=0.515 $X2=0 $Y2=0
cc_445 N_X_c_653_n N_VGND_c_768_n 0.00904371f $X=0.745 $Y=0.515 $X2=0 $Y2=0
cc_446 N_X_c_655_n N_VGND_c_768_n 0.00904371f $X=1.675 $Y=0.515 $X2=0 $Y2=0
cc_447 N_A_968_391#_c_732_n N_A_510_125#_c_852_n 0.00707466f $X=5.94 $Y=2.115
+ $X2=0 $Y2=0
cc_448 N_VGND_c_760_n N_A_510_125#_c_845_n 0.0426691f $X=2.105 $Y=0.515 $X2=0
+ $Y2=0
cc_449 N_VGND_c_761_n N_A_510_125#_c_846_n 0.0137357f $X=5 $Y=0.77 $X2=0 $Y2=0
cc_450 N_VGND_c_765_n N_A_510_125#_c_846_n 0.121756f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_451 N_VGND_c_768_n N_A_510_125#_c_846_n 0.0642692f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_452 N_VGND_c_760_n N_A_510_125#_c_847_n 0.011157f $X=2.105 $Y=0.515 $X2=0
+ $Y2=0
cc_453 N_VGND_c_765_n N_A_510_125#_c_847_n 0.0170431f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_454 N_VGND_c_768_n N_A_510_125#_c_847_n 0.00857552f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_455 N_VGND_c_761_n N_A_510_125#_c_848_n 0.0259901f $X=5 $Y=0.77 $X2=0 $Y2=0
cc_456 N_VGND_M1006_d N_A_510_125#_c_849_n 0.00210887f $X=4.855 $Y=0.625 $X2=0
+ $Y2=0
cc_457 N_VGND_c_761_n N_A_510_125#_c_849_n 0.0179772f $X=5 $Y=0.77 $X2=0 $Y2=0
cc_458 N_VGND_c_761_n N_A_510_125#_c_851_n 0.0132249f $X=5 $Y=0.77 $X2=0 $Y2=0
cc_459 N_VGND_c_762_n N_A_510_125#_c_851_n 0.0127348f $X=5.94 $Y=0.77 $X2=0
+ $Y2=0
cc_460 N_VGND_c_766_n N_A_510_125#_c_851_n 0.00533975f $X=5.775 $Y=0 $X2=0 $Y2=0
cc_461 N_VGND_c_768_n N_A_510_125#_c_851_n 0.00671154f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_462 N_VGND_M1019_s N_A_510_125#_c_852_n 0.00250873f $X=5.8 $Y=0.625 $X2=0
+ $Y2=0
cc_463 N_VGND_c_762_n N_A_510_125#_c_852_n 0.0209867f $X=5.94 $Y=0.77 $X2=0
+ $Y2=0
cc_464 N_VGND_c_762_n N_A_510_125#_c_853_n 0.0133605f $X=5.94 $Y=0.77 $X2=0
+ $Y2=0
cc_465 N_VGND_c_767_n N_A_510_125#_c_853_n 0.00701744f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_466 N_VGND_c_768_n N_A_510_125#_c_853_n 0.0100487f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_467 N_A_510_125#_c_846_n N_A_597_125#_c_918_n 0.0471472f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_468 N_A_510_125#_c_845_n N_A_597_125#_c_919_n 0.00186525f $X=2.695 $Y=0.76
+ $X2=0 $Y2=0
cc_469 N_A_510_125#_c_846_n N_A_597_125#_c_919_n 0.0134458f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_470 N_A_510_125#_c_846_n N_A_597_125#_c_920_n 0.0244253f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_471 N_A_510_125#_c_848_n N_A_597_125#_c_920_n 0.0134764f $X=4.485 $Y=0.77
+ $X2=0 $Y2=0
