* File: sky130_fd_sc_ls__dlrbn_2.pxi.spice
* Created: Fri Aug 28 13:18:03 2020
* 
x_PM_SKY130_FD_SC_LS__DLRBN_2%D N_D_c_176_n N_D_M1009_g N_D_c_181_n N_D_M1013_g
+ D N_D_c_179_n PM_SKY130_FD_SC_LS__DLRBN_2%D
x_PM_SKY130_FD_SC_LS__DLRBN_2%GATE_N N_GATE_N_M1007_g N_GATE_N_c_215_n
+ N_GATE_N_M1006_g N_GATE_N_c_212_n GATE_N N_GATE_N_c_213_n N_GATE_N_c_214_n
+ PM_SKY130_FD_SC_LS__DLRBN_2%GATE_N
x_PM_SKY130_FD_SC_LS__DLRBN_2%A_230_74# N_A_230_74#_M1007_d N_A_230_74#_M1006_d
+ N_A_230_74#_M1019_g N_A_230_74#_c_249_n N_A_230_74#_c_261_n
+ N_A_230_74#_M1022_g N_A_230_74#_M1001_g N_A_230_74#_c_262_n
+ N_A_230_74#_M1000_g N_A_230_74#_c_250_n N_A_230_74#_c_264_n
+ N_A_230_74#_c_251_n N_A_230_74#_c_252_n N_A_230_74#_c_385_p
+ N_A_230_74#_c_253_n N_A_230_74#_c_267_n N_A_230_74#_c_268_n
+ N_A_230_74#_c_269_n N_A_230_74#_c_254_n N_A_230_74#_c_270_n
+ N_A_230_74#_c_255_n N_A_230_74#_c_256_n N_A_230_74#_c_316_p
+ N_A_230_74#_c_257_n N_A_230_74#_c_258_n N_A_230_74#_c_259_n
+ PM_SKY130_FD_SC_LS__DLRBN_2%A_230_74#
x_PM_SKY130_FD_SC_LS__DLRBN_2%A_27_112# N_A_27_112#_M1009_s N_A_27_112#_M1013_s
+ N_A_27_112#_M1002_g N_A_27_112#_c_399_n N_A_27_112#_M1016_g
+ N_A_27_112#_c_400_n N_A_27_112#_c_401_n N_A_27_112#_c_406_n
+ N_A_27_112#_c_418_n N_A_27_112#_c_407_n N_A_27_112#_c_429_n
+ N_A_27_112#_c_451_n N_A_27_112#_c_408_n N_A_27_112#_c_402_n
+ N_A_27_112#_c_409_n N_A_27_112#_c_410_n N_A_27_112#_c_403_n
+ PM_SKY130_FD_SC_LS__DLRBN_2%A_27_112#
x_PM_SKY130_FD_SC_LS__DLRBN_2%A_363_74# N_A_363_74#_M1019_s N_A_363_74#_M1022_s
+ N_A_363_74#_c_509_n N_A_363_74#_M1003_g N_A_363_74#_c_510_n
+ N_A_363_74#_c_511_n N_A_363_74#_M1010_g N_A_363_74#_c_502_n
+ N_A_363_74#_c_503_n N_A_363_74#_c_504_n N_A_363_74#_c_505_n
+ N_A_363_74#_c_506_n N_A_363_74#_c_513_n N_A_363_74#_c_507_n
+ N_A_363_74#_c_508_n PM_SKY130_FD_SC_LS__DLRBN_2%A_363_74#
x_PM_SKY130_FD_SC_LS__DLRBN_2%A_838_48# N_A_838_48#_M1025_s N_A_838_48#_M1015_d
+ N_A_838_48#_c_605_n N_A_838_48#_M1020_g N_A_838_48#_c_606_n
+ N_A_838_48#_c_619_n N_A_838_48#_M1021_g N_A_838_48#_c_607_n
+ N_A_838_48#_c_621_n N_A_838_48#_M1004_g N_A_838_48#_M1012_g
+ N_A_838_48#_c_609_n N_A_838_48#_c_622_n N_A_838_48#_M1023_g
+ N_A_838_48#_M1027_g N_A_838_48#_c_623_n N_A_838_48#_M1005_g
+ N_A_838_48#_M1011_g N_A_838_48#_c_612_n N_A_838_48#_c_613_n
+ N_A_838_48#_c_624_n N_A_838_48#_c_614_n N_A_838_48#_c_626_n
+ N_A_838_48#_c_627_n N_A_838_48#_c_685_p N_A_838_48#_c_628_n
+ N_A_838_48#_c_615_n N_A_838_48#_c_616_n N_A_838_48#_c_617_n
+ PM_SKY130_FD_SC_LS__DLRBN_2%A_838_48#
x_PM_SKY130_FD_SC_LS__DLRBN_2%A_670_74# N_A_670_74#_M1001_d N_A_670_74#_M1003_d
+ N_A_670_74#_c_781_n N_A_670_74#_M1015_g N_A_670_74#_M1025_g
+ N_A_670_74#_c_774_n N_A_670_74#_c_775_n N_A_670_74#_c_776_n
+ N_A_670_74#_c_784_n N_A_670_74#_c_785_n N_A_670_74#_c_777_n
+ N_A_670_74#_c_778_n N_A_670_74#_c_787_n N_A_670_74#_c_779_n
+ N_A_670_74#_c_797_n N_A_670_74#_c_789_n N_A_670_74#_c_780_n
+ N_A_670_74#_c_790_n PM_SKY130_FD_SC_LS__DLRBN_2%A_670_74#
x_PM_SKY130_FD_SC_LS__DLRBN_2%RESET_B N_RESET_B_c_882_n N_RESET_B_M1026_g
+ N_RESET_B_c_883_n N_RESET_B_M1017_g RESET_B
+ PM_SKY130_FD_SC_LS__DLRBN_2%RESET_B
x_PM_SKY130_FD_SC_LS__DLRBN_2%A_1446_368# N_A_1446_368#_M1011_d
+ N_A_1446_368#_M1005_d N_A_1446_368#_c_918_n N_A_1446_368#_M1014_g
+ N_A_1446_368#_c_919_n N_A_1446_368#_M1008_g N_A_1446_368#_c_920_n
+ N_A_1446_368#_c_921_n N_A_1446_368#_c_930_n N_A_1446_368#_M1018_g
+ N_A_1446_368#_c_922_n N_A_1446_368#_M1024_g N_A_1446_368#_c_923_n
+ N_A_1446_368#_c_924_n N_A_1446_368#_c_925_n N_A_1446_368#_c_926_n
+ N_A_1446_368#_c_927_n N_A_1446_368#_c_941_n
+ PM_SKY130_FD_SC_LS__DLRBN_2%A_1446_368#
x_PM_SKY130_FD_SC_LS__DLRBN_2%VPWR N_VPWR_M1013_d N_VPWR_M1022_d N_VPWR_M1021_d
+ N_VPWR_M1017_d N_VPWR_M1023_d N_VPWR_M1008_s N_VPWR_M1018_s N_VPWR_c_988_n
+ N_VPWR_c_989_n N_VPWR_c_990_n N_VPWR_c_991_n N_VPWR_c_992_n N_VPWR_c_993_n
+ N_VPWR_c_994_n N_VPWR_c_995_n N_VPWR_c_996_n VPWR N_VPWR_c_997_n
+ N_VPWR_c_998_n N_VPWR_c_999_n N_VPWR_c_1000_n N_VPWR_c_1001_n N_VPWR_c_1002_n
+ N_VPWR_c_1003_n N_VPWR_c_1004_n N_VPWR_c_1005_n N_VPWR_c_1006_n N_VPWR_c_987_n
+ PM_SKY130_FD_SC_LS__DLRBN_2%VPWR
x_PM_SKY130_FD_SC_LS__DLRBN_2%Q N_Q_M1012_s N_Q_M1004_s N_Q_c_1111_n
+ N_Q_c_1109_n Q PM_SKY130_FD_SC_LS__DLRBN_2%Q
x_PM_SKY130_FD_SC_LS__DLRBN_2%Q_N N_Q_N_M1014_s N_Q_N_M1008_d N_Q_N_c_1145_n Q_N
+ Q_N Q_N Q_N N_Q_N_c_1141_n PM_SKY130_FD_SC_LS__DLRBN_2%Q_N
x_PM_SKY130_FD_SC_LS__DLRBN_2%VGND N_VGND_M1009_d N_VGND_M1019_d N_VGND_M1020_d
+ N_VGND_M1026_d N_VGND_M1027_d N_VGND_M1014_d N_VGND_M1024_d N_VGND_c_1167_n
+ N_VGND_c_1168_n N_VGND_c_1169_n N_VGND_c_1170_n N_VGND_c_1171_n
+ N_VGND_c_1172_n N_VGND_c_1173_n N_VGND_c_1174_n N_VGND_c_1175_n VGND
+ N_VGND_c_1176_n N_VGND_c_1177_n N_VGND_c_1178_n N_VGND_c_1179_n
+ N_VGND_c_1180_n N_VGND_c_1181_n N_VGND_c_1182_n N_VGND_c_1183_n
+ N_VGND_c_1184_n N_VGND_c_1185_n N_VGND_c_1186_n N_VGND_c_1187_n
+ PM_SKY130_FD_SC_LS__DLRBN_2%VGND
cc_1 VNB N_D_c_176_n 0.0161132f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.76
cc_2 VNB N_D_M1009_g 0.0253508f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_3 VNB D 0.00288429f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_D_c_179_n 0.0185146f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.425
cc_5 VNB N_GATE_N_M1007_g 0.025295f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.26
cc_6 VNB N_GATE_N_c_212_n 0.0176964f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_7 VNB N_GATE_N_c_213_n 0.0178601f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.425
cc_8 VNB N_GATE_N_c_214_n 0.00223122f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.26
cc_9 VNB N_A_230_74#_c_249_n 0.00267921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_230_74#_c_250_n 0.00969645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_230_74#_c_251_n 6.76447e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_230_74#_c_252_n 0.0222345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_230_74#_c_253_n 0.00368107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_230_74#_c_254_n 0.0154535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_230_74#_c_255_n 0.00580321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_230_74#_c_256_n 0.0354769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_230_74#_c_257_n 0.0305451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_230_74#_c_258_n 0.0228564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_230_74#_c_259_n 0.0189144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_112#_M1002_g 0.0368093f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_21 VNB N_A_27_112#_c_399_n 0.0198227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_112#_c_400_n 0.0185219f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.425
cc_23 VNB N_A_27_112#_c_401_n 0.0266292f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.595
cc_24 VNB N_A_27_112#_c_402_n 0.00710642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_112#_c_403_n 0.00162179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_363_74#_M1010_g 0.0358196f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.425
cc_27 VNB N_A_363_74#_c_502_n 0.00629876f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.595
cc_28 VNB N_A_363_74#_c_503_n 0.00990916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_363_74#_c_504_n 0.00402727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_363_74#_c_505_n 0.0027542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_363_74#_c_506_n 0.00153707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_363_74#_c_507_n 0.00530228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_363_74#_c_508_n 0.038505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_838_48#_c_605_n 0.0163494f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.045
cc_35 VNB N_A_838_48#_c_606_n 0.0350078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_838_48#_c_607_n 0.00912119f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.595
cc_37 VNB N_A_838_48#_M1012_g 0.0230556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_838_48#_c_609_n 0.0091229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_838_48#_M1027_g 0.0230016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_838_48#_M1011_g 0.0320384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_838_48#_c_612_n 0.0223826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_838_48#_c_613_n 0.00731011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_838_48#_c_614_n 0.0037738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_838_48#_c_615_n 0.0142822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_838_48#_c_616_n 0.00201541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_838_48#_c_617_n 0.0513367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_670_74#_M1025_g 0.0266948f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.425
cc_48 VNB N_A_670_74#_c_774_n 0.0303389f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.425
cc_49 VNB N_A_670_74#_c_775_n 0.0104774f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.26
cc_50 VNB N_A_670_74#_c_776_n 0.00594597f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.595
cc_51 VNB N_A_670_74#_c_777_n 8.83266e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_670_74#_c_778_n 0.00488861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_670_74#_c_779_n 0.00740554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_670_74#_c_780_n 0.00458916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_RESET_B_c_882_n 0.017547f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.43
cc_56 VNB N_RESET_B_c_883_n 0.0354835f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_57 VNB RESET_B 0.0173431f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.045
cc_58 VNB N_A_1446_368#_c_918_n 0.0193826f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.045
cc_59 VNB N_A_1446_368#_c_919_n 0.0160298f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_60 VNB N_A_1446_368#_c_920_n 0.0112701f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.425
cc_61 VNB N_A_1446_368#_c_921_n 0.0160627f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.595
cc_62 VNB N_A_1446_368#_c_922_n 0.0204036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1446_368#_c_923_n 0.0621023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1446_368#_c_924_n 0.0186247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1446_368#_c_925_n 0.0114111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1446_368#_c_926_n 0.00155823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1446_368#_c_927_n 0.00222672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VPWR_c_987_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_Q_c_1109_n 0.00244275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB Q 0.00387264f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.425
cc_71 VNB N_Q_N_c_1141_n 0.00320587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1167_n 0.0168478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1168_n 0.0131928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1169_n 0.006605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1170_n 0.0112424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1171_n 0.0157081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1172_n 0.0108703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1173_n 0.0513343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1174_n 0.0291058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1175_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1176_n 0.020108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1177_n 0.036157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1178_n 0.0425683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1179_n 0.0241211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1180_n 0.0206041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1181_n 0.02253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1182_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1183_n 0.0189263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1184_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1185_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1186_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1187_n 0.520754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VPB N_D_c_176_n 0.031681f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.76
cc_94 VPB N_D_c_181_n 0.0221378f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_95 VPB D 0.00209841f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_96 VPB N_GATE_N_c_215_n 0.0213417f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.835
cc_97 VPB N_GATE_N_c_212_n 0.03364f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_98 VPB N_GATE_N_c_214_n 0.00148103f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.26
cc_99 VPB N_A_230_74#_c_249_n 0.0108612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_230_74#_c_261_n 0.025597f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.425
cc_101 VPB N_A_230_74#_c_262_n 0.063867f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.595
cc_102 VPB N_A_230_74#_c_250_n 0.0123488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_230_74#_c_264_n 0.00961418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_230_74#_c_251_n 0.00195002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_230_74#_c_253_n 0.00241401f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_230_74#_c_267_n 0.00632058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_230_74#_c_268_n 0.00211104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_230_74#_c_269_n 0.00407213f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_230_74#_c_270_n 0.0103296f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_27_112#_c_399_n 0.0363734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_27_112#_c_401_n 0.0207356f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.595
cc_112 VPB N_A_27_112#_c_406_n 0.00798527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_27_112#_c_407_n 0.00714322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_27_112#_c_408_n 0.00104736f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_112#_c_409_n 0.0450025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_27_112#_c_410_n 0.00502212f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_363_74#_c_509_n 0.0146907f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_118 VPB N_A_363_74#_c_510_n 0.0309149f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_119 VPB N_A_363_74#_c_511_n 0.01f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_363_74#_c_503_n 0.00382545f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_363_74#_c_513_n 0.00971474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_363_74#_c_508_n 0.00879292f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_838_48#_c_606_n 0.0273201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_838_48#_c_619_n 0.0570552f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.425
cc_125 VPB N_A_838_48#_c_607_n 7.38289e-19 $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.595
cc_126 VPB N_A_838_48#_c_621_n 0.0209486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_838_48#_c_622_n 0.0168214f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_838_48#_c_623_n 0.0172751f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_838_48#_c_624_n 0.00579102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_838_48#_c_614_n 0.00157737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_838_48#_c_626_n 0.00732891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_838_48#_c_627_n 0.00265926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_838_48#_c_628_n 0.00264805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_838_48#_c_617_n 0.0148614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_670_74#_c_781_n 0.017589f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_136 VPB N_A_670_74#_c_774_n 0.0129544f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.425
cc_137 VPB N_A_670_74#_c_775_n 0.00663917f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.26
cc_138 VPB N_A_670_74#_c_784_n 0.0139502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_670_74#_c_785_n 2.40333e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_670_74#_c_778_n 5.47069e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_670_74#_c_787_n 0.010915f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_670_74#_c_779_n 3.3123e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_670_74#_c_789_n 0.00315717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_670_74#_c_790_n 0.00301383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_RESET_B_c_883_n 0.0235413f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.835
cc_146 VPB N_A_1446_368#_c_919_n 0.0246718f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_147 VPB N_A_1446_368#_c_921_n 0.00111912f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.595
cc_148 VPB N_A_1446_368#_c_930_n 0.0258516f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_1446_368#_c_926_n 0.015382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_988_n 0.0082415f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_989_n 0.0137119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_990_n 0.00514606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_991_n 0.010436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_992_n 0.0249297f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_993_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_994_n 0.0645677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_995_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_996_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_997_n 0.0437096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_998_n 0.0446611f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_999_n 0.0187066f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_1000_n 0.0213015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1001_n 0.0204479f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_1002_n 0.0231158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_1003_n 0.00631708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1004_n 0.0204849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_1005_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1006_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_987_n 0.12856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_Q_c_1111_n 0.00365896f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_171 VPB N_Q_c_1109_n 0.00137598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB Q_N 0.00404267f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.425
cc_173 VPB Q_N 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_Q_N_c_1141_n 0.00151138f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 N_D_M1009_g N_GATE_N_M1007_g 0.0178869f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_176 N_D_c_181_n N_GATE_N_c_215_n 0.0143522f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_177 N_D_c_176_n N_GATE_N_c_212_n 0.0244018f $X=0.585 $Y=1.76 $X2=0 $Y2=0
cc_178 D N_GATE_N_c_213_n 0.00389099f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_179 N_D_c_179_n N_GATE_N_c_213_n 0.0208612f $X=0.59 $Y=1.425 $X2=0 $Y2=0
cc_180 D N_GATE_N_c_214_n 0.0534095f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_181 N_D_c_179_n N_GATE_N_c_214_n 7.38266e-19 $X=0.59 $Y=1.425 $X2=0 $Y2=0
cc_182 N_D_M1009_g N_A_27_112#_c_400_n 0.00590244f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_183 N_D_M1009_g N_A_27_112#_c_401_n 0.00411368f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_184 D N_A_27_112#_c_401_n 0.0509214f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_185 N_D_c_179_n N_A_27_112#_c_401_n 0.0193371f $X=0.59 $Y=1.425 $X2=0 $Y2=0
cc_186 N_D_c_176_n N_A_27_112#_c_406_n 0.00460733f $X=0.585 $Y=1.76 $X2=0 $Y2=0
cc_187 N_D_c_181_n N_A_27_112#_c_406_n 0.0129287f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_188 D N_A_27_112#_c_406_n 0.028288f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_189 N_D_c_181_n N_A_27_112#_c_418_n 0.00160792f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_190 N_D_M1009_g N_A_27_112#_c_402_n 0.00408614f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_191 D N_A_27_112#_c_402_n 0.00157312f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_192 N_D_c_176_n N_A_27_112#_c_409_n 7.04954e-19 $X=0.585 $Y=1.76 $X2=0 $Y2=0
cc_193 N_D_c_181_n N_A_27_112#_c_409_n 0.0134076f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_194 D N_A_27_112#_c_409_n 0.00170517f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_195 N_D_c_181_n N_VPWR_c_988_n 0.0056519f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_196 N_D_c_181_n N_VPWR_c_1002_n 0.00445602f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_197 N_D_c_181_n N_VPWR_c_987_n 0.00862861f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_198 N_D_M1009_g N_VGND_c_1167_n 0.00658895f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_199 D N_VGND_c_1167_n 0.0157345f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_200 N_D_c_179_n N_VGND_c_1167_n 0.00346007f $X=0.59 $Y=1.425 $X2=0 $Y2=0
cc_201 N_D_M1009_g N_VGND_c_1176_n 0.0043356f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_202 N_D_M1009_g N_VGND_c_1187_n 0.00487769f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_203 N_GATE_N_M1007_g N_A_230_74#_c_250_n 0.00471659f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_204 N_GATE_N_c_215_n N_A_230_74#_c_250_n 0.00181649f $X=1.185 $Y=2.045 $X2=0
+ $Y2=0
cc_205 N_GATE_N_c_212_n N_A_230_74#_c_250_n 0.00397658f $X=1.13 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_GATE_N_c_213_n N_A_230_74#_c_250_n 0.0151579f $X=1.13 $Y=1.425 $X2=0
+ $Y2=0
cc_207 N_GATE_N_c_214_n N_A_230_74#_c_250_n 0.0500404f $X=1.13 $Y=1.425 $X2=0
+ $Y2=0
cc_208 N_GATE_N_M1007_g N_A_230_74#_c_254_n 0.00910897f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_209 N_GATE_N_c_213_n N_A_230_74#_c_254_n 0.00140316f $X=1.13 $Y=1.425 $X2=0
+ $Y2=0
cc_210 N_GATE_N_c_214_n N_A_230_74#_c_254_n 0.0111169f $X=1.13 $Y=1.425 $X2=0
+ $Y2=0
cc_211 N_GATE_N_c_215_n N_A_230_74#_c_270_n 0.00164325f $X=1.185 $Y=2.045 $X2=0
+ $Y2=0
cc_212 N_GATE_N_c_215_n N_A_27_112#_c_406_n 0.00578906f $X=1.185 $Y=2.045 $X2=0
+ $Y2=0
cc_213 N_GATE_N_c_212_n N_A_27_112#_c_406_n 0.00184207f $X=1.13 $Y=1.765 $X2=0
+ $Y2=0
cc_214 N_GATE_N_c_214_n N_A_27_112#_c_406_n 0.015685f $X=1.13 $Y=1.425 $X2=0
+ $Y2=0
cc_215 N_GATE_N_c_215_n N_A_27_112#_c_418_n 0.0107332f $X=1.185 $Y=2.045 $X2=0
+ $Y2=0
cc_216 N_GATE_N_c_215_n N_A_27_112#_c_407_n 0.0118423f $X=1.185 $Y=2.045 $X2=0
+ $Y2=0
cc_217 N_GATE_N_c_215_n N_A_27_112#_c_429_n 0.0034142f $X=1.185 $Y=2.045 $X2=0
+ $Y2=0
cc_218 N_GATE_N_c_215_n N_A_27_112#_c_409_n 2.16358e-19 $X=1.185 $Y=2.045 $X2=0
+ $Y2=0
cc_219 N_GATE_N_c_215_n N_A_27_112#_c_410_n 0.00292174f $X=1.185 $Y=2.045 $X2=0
+ $Y2=0
cc_220 N_GATE_N_M1007_g N_A_363_74#_c_502_n 5.41378e-19 $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_221 N_GATE_N_c_215_n N_VPWR_c_988_n 0.00637675f $X=1.185 $Y=2.045 $X2=0 $Y2=0
cc_222 N_GATE_N_c_215_n N_VPWR_c_997_n 0.00311972f $X=1.185 $Y=2.045 $X2=0 $Y2=0
cc_223 N_GATE_N_c_215_n N_VPWR_c_987_n 0.00392193f $X=1.185 $Y=2.045 $X2=0 $Y2=0
cc_224 N_GATE_N_M1007_g N_VGND_c_1167_n 0.0103395f $X=1.075 $Y=0.74 $X2=0 $Y2=0
cc_225 N_GATE_N_M1007_g N_VGND_c_1177_n 0.00434272f $X=1.075 $Y=0.74 $X2=0 $Y2=0
cc_226 N_GATE_N_M1007_g N_VGND_c_1187_n 0.00830058f $X=1.075 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A_230_74#_c_252_n N_A_27_112#_M1002_g 0.014698f $X=3.155 $Y=1.215 $X2=0
+ $Y2=0
cc_228 N_A_230_74#_c_255_n N_A_27_112#_M1002_g 0.00358507f $X=2.305 $Y=1.215
+ $X2=0 $Y2=0
cc_229 N_A_230_74#_c_256_n N_A_27_112#_M1002_g 0.00767944f $X=2.285 $Y=1.385
+ $X2=0 $Y2=0
cc_230 N_A_230_74#_c_258_n N_A_27_112#_M1002_g 0.0178599f $X=2.275 $Y=1.22 $X2=0
+ $Y2=0
cc_231 N_A_230_74#_c_259_n N_A_27_112#_M1002_g 0.065042f $X=3.365 $Y=1.12 $X2=0
+ $Y2=0
cc_232 N_A_230_74#_c_249_n N_A_27_112#_c_399_n 0.0102232f $X=2.28 $Y=1.795 $X2=0
+ $Y2=0
cc_233 N_A_230_74#_c_261_n N_A_27_112#_c_399_n 0.0244726f $X=2.28 $Y=1.885 $X2=0
+ $Y2=0
cc_234 N_A_230_74#_c_264_n N_A_27_112#_c_399_n 5.39985e-19 $X=2.305 $Y=2.225
+ $X2=0 $Y2=0
cc_235 N_A_230_74#_c_251_n N_A_27_112#_c_399_n 8.59566e-19 $X=2.39 $Y=2.14 $X2=0
+ $Y2=0
cc_236 N_A_230_74#_c_252_n N_A_27_112#_c_399_n 0.00144981f $X=3.155 $Y=1.215
+ $X2=0 $Y2=0
cc_237 N_A_230_74#_c_253_n N_A_27_112#_c_399_n 0.00668225f $X=3.24 $Y=1.97 $X2=0
+ $Y2=0
cc_238 N_A_230_74#_c_268_n N_A_27_112#_c_399_n 0.00131424f $X=3.18 $Y=2.99 $X2=0
+ $Y2=0
cc_239 N_A_230_74#_c_255_n N_A_27_112#_c_399_n 0.00203002f $X=2.305 $Y=1.215
+ $X2=0 $Y2=0
cc_240 N_A_230_74#_c_256_n N_A_27_112#_c_399_n 0.0050142f $X=2.285 $Y=1.385
+ $X2=0 $Y2=0
cc_241 N_A_230_74#_c_270_n N_A_27_112#_c_406_n 0.0145981f $X=1.625 $Y=2.29 $X2=0
+ $Y2=0
cc_242 N_A_230_74#_c_270_n N_A_27_112#_c_418_n 0.0155954f $X=1.625 $Y=2.29 $X2=0
+ $Y2=0
cc_243 N_A_230_74#_M1006_d N_A_27_112#_c_407_n 0.00734801f $X=1.26 $Y=2.12 $X2=0
+ $Y2=0
cc_244 N_A_230_74#_c_264_n N_A_27_112#_c_407_n 0.00790193f $X=2.305 $Y=2.225
+ $X2=0 $Y2=0
cc_245 N_A_230_74#_c_270_n N_A_27_112#_c_407_n 0.022752f $X=1.625 $Y=2.29 $X2=0
+ $Y2=0
cc_246 N_A_230_74#_c_261_n N_A_27_112#_c_451_n 0.0135857f $X=2.28 $Y=1.885 $X2=0
+ $Y2=0
cc_247 N_A_230_74#_c_264_n N_A_27_112#_c_451_n 0.0288493f $X=2.305 $Y=2.225
+ $X2=0 $Y2=0
cc_248 N_A_230_74#_c_261_n N_A_27_112#_c_408_n 0.00465064f $X=2.28 $Y=1.885
+ $X2=0 $Y2=0
cc_249 N_A_230_74#_c_264_n N_A_27_112#_c_408_n 0.0129839f $X=2.305 $Y=2.225
+ $X2=0 $Y2=0
cc_250 N_A_230_74#_c_251_n N_A_27_112#_c_408_n 0.0235411f $X=2.39 $Y=2.14 $X2=0
+ $Y2=0
cc_251 N_A_230_74#_c_253_n N_A_27_112#_c_408_n 0.00745183f $X=3.24 $Y=1.97 $X2=0
+ $Y2=0
cc_252 N_A_230_74#_c_261_n N_A_27_112#_c_410_n 0.00610769f $X=2.28 $Y=1.885
+ $X2=0 $Y2=0
cc_253 N_A_230_74#_c_264_n N_A_27_112#_c_410_n 0.0130148f $X=2.305 $Y=2.225
+ $X2=0 $Y2=0
cc_254 N_A_230_74#_c_249_n N_A_27_112#_c_403_n 2.68674e-19 $X=2.28 $Y=1.795
+ $X2=0 $Y2=0
cc_255 N_A_230_74#_c_252_n N_A_27_112#_c_403_n 0.0245759f $X=3.155 $Y=1.215
+ $X2=0 $Y2=0
cc_256 N_A_230_74#_c_253_n N_A_27_112#_c_403_n 0.0247726f $X=3.24 $Y=1.97 $X2=0
+ $Y2=0
cc_257 N_A_230_74#_c_255_n N_A_27_112#_c_403_n 0.0235411f $X=2.305 $Y=1.215
+ $X2=0 $Y2=0
cc_258 N_A_230_74#_c_264_n N_A_363_74#_M1022_s 0.008749f $X=2.305 $Y=2.225 $X2=0
+ $Y2=0
cc_259 N_A_230_74#_c_262_n N_A_363_74#_c_509_n 0.0209658f $X=3.84 $Y=2.465 $X2=0
+ $Y2=0
cc_260 N_A_230_74#_c_253_n N_A_363_74#_c_509_n 0.00204355f $X=3.24 $Y=1.97 $X2=0
+ $Y2=0
cc_261 N_A_230_74#_c_267_n N_A_363_74#_c_509_n 0.013189f $X=3.835 $Y=2.99 $X2=0
+ $Y2=0
cc_262 N_A_230_74#_c_269_n N_A_363_74#_c_509_n 5.06441e-19 $X=4 $Y=2.215 $X2=0
+ $Y2=0
cc_263 N_A_230_74#_c_316_p N_A_363_74#_c_509_n 0.00916584f $X=3.24 $Y=2.055
+ $X2=0 $Y2=0
cc_264 N_A_230_74#_c_262_n N_A_363_74#_c_510_n 0.0130722f $X=3.84 $Y=2.465 $X2=0
+ $Y2=0
cc_265 N_A_230_74#_c_252_n N_A_363_74#_c_511_n 0.00125752f $X=3.155 $Y=1.215
+ $X2=0 $Y2=0
cc_266 N_A_230_74#_c_253_n N_A_363_74#_c_511_n 0.00722355f $X=3.24 $Y=1.97 $X2=0
+ $Y2=0
cc_267 N_A_230_74#_c_257_n N_A_363_74#_c_511_n 0.0175343f $X=3.365 $Y=1.285
+ $X2=0 $Y2=0
cc_268 N_A_230_74#_c_257_n N_A_363_74#_M1010_g 0.0149209f $X=3.365 $Y=1.285
+ $X2=0 $Y2=0
cc_269 N_A_230_74#_c_259_n N_A_363_74#_M1010_g 0.022907f $X=3.365 $Y=1.12 $X2=0
+ $Y2=0
cc_270 N_A_230_74#_c_254_n N_A_363_74#_c_502_n 0.0369241f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_271 N_A_230_74#_c_258_n N_A_363_74#_c_502_n 0.00725643f $X=2.275 $Y=1.22
+ $X2=0 $Y2=0
cc_272 N_A_230_74#_c_249_n N_A_363_74#_c_503_n 0.00343183f $X=2.28 $Y=1.795
+ $X2=0 $Y2=0
cc_273 N_A_230_74#_c_251_n N_A_363_74#_c_503_n 0.00724105f $X=2.39 $Y=2.14 $X2=0
+ $Y2=0
cc_274 N_A_230_74#_c_254_n N_A_363_74#_c_503_n 0.0580213f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_275 N_A_230_74#_c_255_n N_A_363_74#_c_503_n 0.0315988f $X=2.305 $Y=1.215
+ $X2=0 $Y2=0
cc_276 N_A_230_74#_c_258_n N_A_363_74#_c_503_n 0.0136738f $X=2.275 $Y=1.22 $X2=0
+ $Y2=0
cc_277 N_A_230_74#_c_252_n N_A_363_74#_c_504_n 0.0675138f $X=3.155 $Y=1.215
+ $X2=0 $Y2=0
cc_278 N_A_230_74#_c_255_n N_A_363_74#_c_504_n 0.0236679f $X=2.305 $Y=1.215
+ $X2=0 $Y2=0
cc_279 N_A_230_74#_c_256_n N_A_363_74#_c_504_n 9.91944e-19 $X=2.285 $Y=1.385
+ $X2=0 $Y2=0
cc_280 N_A_230_74#_c_257_n N_A_363_74#_c_504_n 0.00113748f $X=3.365 $Y=1.285
+ $X2=0 $Y2=0
cc_281 N_A_230_74#_c_258_n N_A_363_74#_c_504_n 0.00981853f $X=2.275 $Y=1.22
+ $X2=0 $Y2=0
cc_282 N_A_230_74#_c_259_n N_A_363_74#_c_504_n 0.0119591f $X=3.365 $Y=1.12 $X2=0
+ $Y2=0
cc_283 N_A_230_74#_c_252_n N_A_363_74#_c_505_n 0.00747745f $X=3.155 $Y=1.215
+ $X2=0 $Y2=0
cc_284 N_A_230_74#_c_257_n N_A_363_74#_c_505_n 6.36324e-19 $X=3.365 $Y=1.285
+ $X2=0 $Y2=0
cc_285 N_A_230_74#_c_259_n N_A_363_74#_c_505_n 0.00297915f $X=3.365 $Y=1.12
+ $X2=0 $Y2=0
cc_286 N_A_230_74#_c_254_n N_A_363_74#_c_506_n 0.0163625f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_287 N_A_230_74#_c_258_n N_A_363_74#_c_506_n 0.00173383f $X=2.275 $Y=1.22
+ $X2=0 $Y2=0
cc_288 N_A_230_74#_c_249_n N_A_363_74#_c_513_n 0.0037919f $X=2.28 $Y=1.795 $X2=0
+ $Y2=0
cc_289 N_A_230_74#_c_261_n N_A_363_74#_c_513_n 0.00183029f $X=2.28 $Y=1.885
+ $X2=0 $Y2=0
cc_290 N_A_230_74#_c_250_n N_A_363_74#_c_513_n 0.0198009f $X=1.54 $Y=2.1 $X2=0
+ $Y2=0
cc_291 N_A_230_74#_c_264_n N_A_363_74#_c_513_n 0.025473f $X=2.305 $Y=2.225 $X2=0
+ $Y2=0
cc_292 N_A_230_74#_c_251_n N_A_363_74#_c_513_n 0.0187806f $X=2.39 $Y=2.14 $X2=0
+ $Y2=0
cc_293 N_A_230_74#_c_256_n N_A_363_74#_c_513_n 0.0015091f $X=2.285 $Y=1.385
+ $X2=0 $Y2=0
cc_294 N_A_230_74#_c_252_n N_A_363_74#_c_507_n 0.0171782f $X=3.155 $Y=1.215
+ $X2=0 $Y2=0
cc_295 N_A_230_74#_c_253_n N_A_363_74#_c_507_n 0.00403635f $X=3.24 $Y=1.97 $X2=0
+ $Y2=0
cc_296 N_A_230_74#_c_257_n N_A_363_74#_c_507_n 0.00147537f $X=3.365 $Y=1.285
+ $X2=0 $Y2=0
cc_297 N_A_230_74#_c_262_n N_A_363_74#_c_508_n 0.0033105f $X=3.84 $Y=2.465 $X2=0
+ $Y2=0
cc_298 N_A_230_74#_c_252_n N_A_363_74#_c_508_n 2.45285e-19 $X=3.155 $Y=1.215
+ $X2=0 $Y2=0
cc_299 N_A_230_74#_c_253_n N_A_363_74#_c_508_n 0.00423603f $X=3.24 $Y=1.97 $X2=0
+ $Y2=0
cc_300 N_A_230_74#_c_262_n N_A_838_48#_c_619_n 0.0349741f $X=3.84 $Y=2.465 $X2=0
+ $Y2=0
cc_301 N_A_230_74#_c_267_n N_A_838_48#_c_619_n 0.001726f $X=3.835 $Y=2.99 $X2=0
+ $Y2=0
cc_302 N_A_230_74#_c_269_n N_A_838_48#_c_619_n 0.00940072f $X=4 $Y=2.215 $X2=0
+ $Y2=0
cc_303 N_A_230_74#_c_262_n N_A_838_48#_c_624_n 0.00108139f $X=3.84 $Y=2.465
+ $X2=0 $Y2=0
cc_304 N_A_230_74#_c_269_n N_A_838_48#_c_624_n 0.0200695f $X=4 $Y=2.215 $X2=0
+ $Y2=0
cc_305 N_A_230_74#_c_267_n N_A_670_74#_M1003_d 0.00437091f $X=3.835 $Y=2.99
+ $X2=0 $Y2=0
cc_306 N_A_230_74#_c_259_n N_A_670_74#_c_776_n 0.00887218f $X=3.365 $Y=1.12
+ $X2=0 $Y2=0
cc_307 N_A_230_74#_c_262_n N_A_670_74#_c_784_n 0.00304809f $X=3.84 $Y=2.465
+ $X2=0 $Y2=0
cc_308 N_A_230_74#_c_269_n N_A_670_74#_c_784_n 0.0262124f $X=4 $Y=2.215 $X2=0
+ $Y2=0
cc_309 N_A_230_74#_c_252_n N_A_670_74#_c_785_n 0.00193642f $X=3.155 $Y=1.215
+ $X2=0 $Y2=0
cc_310 N_A_230_74#_c_253_n N_A_670_74#_c_785_n 0.0131299f $X=3.24 $Y=1.97 $X2=0
+ $Y2=0
cc_311 N_A_230_74#_c_262_n N_A_670_74#_c_797_n 0.00219249f $X=3.84 $Y=2.465
+ $X2=0 $Y2=0
cc_312 N_A_230_74#_c_267_n N_A_670_74#_c_797_n 0.0190351f $X=3.835 $Y=2.99 $X2=0
+ $Y2=0
cc_313 N_A_230_74#_c_262_n N_A_670_74#_c_789_n 0.00373541f $X=3.84 $Y=2.465
+ $X2=0 $Y2=0
cc_314 N_A_230_74#_c_253_n N_A_670_74#_c_789_n 0.00635216f $X=3.24 $Y=1.97 $X2=0
+ $Y2=0
cc_315 N_A_230_74#_c_269_n N_A_670_74#_c_789_n 0.0516627f $X=4 $Y=2.215 $X2=0
+ $Y2=0
cc_316 N_A_230_74#_c_316_p N_A_670_74#_c_789_n 0.0124226f $X=3.24 $Y=2.055 $X2=0
+ $Y2=0
cc_317 N_A_230_74#_c_264_n N_VPWR_M1022_d 0.00232895f $X=2.305 $Y=2.225 $X2=0
+ $Y2=0
cc_318 N_A_230_74#_c_251_n N_VPWR_M1022_d 0.00165969f $X=2.39 $Y=2.14 $X2=0
+ $Y2=0
cc_319 N_A_230_74#_c_261_n N_VPWR_c_989_n 0.00317424f $X=2.28 $Y=1.885 $X2=0
+ $Y2=0
cc_320 N_A_230_74#_c_268_n N_VPWR_c_989_n 0.00925116f $X=3.18 $Y=2.99 $X2=0
+ $Y2=0
cc_321 N_A_230_74#_c_261_n N_VPWR_c_997_n 0.0036399f $X=2.28 $Y=1.885 $X2=0
+ $Y2=0
cc_322 N_A_230_74#_c_262_n N_VPWR_c_998_n 0.00278193f $X=3.84 $Y=2.465 $X2=0
+ $Y2=0
cc_323 N_A_230_74#_c_267_n N_VPWR_c_998_n 0.064841f $X=3.835 $Y=2.99 $X2=0 $Y2=0
cc_324 N_A_230_74#_c_268_n N_VPWR_c_998_n 0.0121867f $X=3.18 $Y=2.99 $X2=0 $Y2=0
cc_325 N_A_230_74#_c_262_n N_VPWR_c_1004_n 4.07803e-19 $X=3.84 $Y=2.465 $X2=0
+ $Y2=0
cc_326 N_A_230_74#_c_267_n N_VPWR_c_1004_n 0.00844737f $X=3.835 $Y=2.99 $X2=0
+ $Y2=0
cc_327 N_A_230_74#_c_269_n N_VPWR_c_1004_n 0.0116264f $X=4 $Y=2.215 $X2=0 $Y2=0
cc_328 N_A_230_74#_c_261_n N_VPWR_c_987_n 0.0049649f $X=2.28 $Y=1.885 $X2=0
+ $Y2=0
cc_329 N_A_230_74#_c_262_n N_VPWR_c_987_n 0.00356158f $X=3.84 $Y=2.465 $X2=0
+ $Y2=0
cc_330 N_A_230_74#_c_267_n N_VPWR_c_987_n 0.0360768f $X=3.835 $Y=2.99 $X2=0
+ $Y2=0
cc_331 N_A_230_74#_c_268_n N_VPWR_c_987_n 0.00660921f $X=3.18 $Y=2.99 $X2=0
+ $Y2=0
cc_332 N_A_230_74#_c_385_p A_595_392# 0.00326441f $X=3.095 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_333 N_A_230_74#_c_316_p A_595_392# 0.00283134f $X=3.24 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_334 N_A_230_74#_c_267_n A_783_508# 8.83155e-19 $X=3.835 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_335 N_A_230_74#_c_269_n A_783_508# 0.00570902f $X=4 $Y=2.215 $X2=-0.19
+ $Y2=-0.245
cc_336 N_A_230_74#_c_254_n N_VGND_c_1167_n 0.0303788f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_337 N_A_230_74#_c_254_n N_VGND_c_1177_n 0.0221495f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_338 N_A_230_74#_c_258_n N_VGND_c_1177_n 0.00434272f $X=2.275 $Y=1.22 $X2=0
+ $Y2=0
cc_339 N_A_230_74#_c_259_n N_VGND_c_1178_n 0.00433387f $X=3.365 $Y=1.12 $X2=0
+ $Y2=0
cc_340 N_A_230_74#_c_258_n N_VGND_c_1183_n 0.00563529f $X=2.275 $Y=1.22 $X2=0
+ $Y2=0
cc_341 N_A_230_74#_c_259_n N_VGND_c_1183_n 0.00128674f $X=3.365 $Y=1.12 $X2=0
+ $Y2=0
cc_342 N_A_230_74#_c_254_n N_VGND_c_1187_n 0.018277f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_343 N_A_230_74#_c_258_n N_VGND_c_1187_n 0.00439489f $X=2.275 $Y=1.22 $X2=0
+ $Y2=0
cc_344 N_A_230_74#_c_259_n N_VGND_c_1187_n 0.00435873f $X=3.365 $Y=1.12 $X2=0
+ $Y2=0
cc_345 N_A_27_112#_c_451_n N_A_363_74#_M1022_s 0.00635501f $X=2.66 $Y=2.565
+ $X2=0 $Y2=0
cc_346 N_A_27_112#_c_410_n N_A_363_74#_M1022_s 0.00623236f $X=1.88 $Y=2.565
+ $X2=0 $Y2=0
cc_347 N_A_27_112#_c_399_n N_A_363_74#_c_509_n 0.0547826f $X=2.9 $Y=1.885 $X2=0
+ $Y2=0
cc_348 N_A_27_112#_c_408_n N_A_363_74#_c_509_n 3.16254e-19 $X=2.745 $Y=2.48
+ $X2=0 $Y2=0
cc_349 N_A_27_112#_c_399_n N_A_363_74#_c_511_n 0.0119877f $X=2.9 $Y=1.885 $X2=0
+ $Y2=0
cc_350 N_A_27_112#_M1002_g N_A_363_74#_c_502_n 9.02769e-19 $X=2.885 $Y=0.69
+ $X2=0 $Y2=0
cc_351 N_A_27_112#_M1002_g N_A_363_74#_c_504_n 0.0124067f $X=2.885 $Y=0.69 $X2=0
+ $Y2=0
cc_352 N_A_27_112#_M1002_g N_A_670_74#_c_776_n 7.17942e-19 $X=2.885 $Y=0.69
+ $X2=0 $Y2=0
cc_353 N_A_27_112#_c_406_n N_VPWR_M1013_d 0.0100177f $X=0.985 $Y=2.185 $X2=-0.19
+ $Y2=-0.245
cc_354 N_A_27_112#_c_418_n N_VPWR_M1013_d 0.00429376f $X=1.07 $Y=2.65 $X2=-0.19
+ $Y2=-0.245
cc_355 N_A_27_112#_c_429_n N_VPWR_M1013_d 0.00267641f $X=1.155 $Y=2.735
+ $X2=-0.19 $Y2=-0.245
cc_356 N_A_27_112#_c_451_n N_VPWR_M1022_d 0.0125866f $X=2.66 $Y=2.565 $X2=0
+ $Y2=0
cc_357 N_A_27_112#_c_408_n N_VPWR_M1022_d 0.00536652f $X=2.745 $Y=2.48 $X2=0
+ $Y2=0
cc_358 N_A_27_112#_c_406_n N_VPWR_c_988_n 0.0136682f $X=0.985 $Y=2.185 $X2=0
+ $Y2=0
cc_359 N_A_27_112#_c_418_n N_VPWR_c_988_n 0.0152166f $X=1.07 $Y=2.65 $X2=0 $Y2=0
cc_360 N_A_27_112#_c_429_n N_VPWR_c_988_n 0.0138309f $X=1.155 $Y=2.735 $X2=0
+ $Y2=0
cc_361 N_A_27_112#_c_409_n N_VPWR_c_988_n 0.0354398f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_362 N_A_27_112#_c_399_n N_VPWR_c_989_n 0.005161f $X=2.9 $Y=1.885 $X2=0 $Y2=0
cc_363 N_A_27_112#_c_451_n N_VPWR_c_989_n 0.0260645f $X=2.66 $Y=2.565 $X2=0
+ $Y2=0
cc_364 N_A_27_112#_c_407_n N_VPWR_c_997_n 0.0145908f $X=1.795 $Y=2.735 $X2=0
+ $Y2=0
cc_365 N_A_27_112#_c_429_n N_VPWR_c_997_n 0.00366075f $X=1.155 $Y=2.735 $X2=0
+ $Y2=0
cc_366 N_A_27_112#_c_451_n N_VPWR_c_997_n 0.00629534f $X=2.66 $Y=2.565 $X2=0
+ $Y2=0
cc_367 N_A_27_112#_c_410_n N_VPWR_c_997_n 0.00430904f $X=1.88 $Y=2.565 $X2=0
+ $Y2=0
cc_368 N_A_27_112#_c_399_n N_VPWR_c_998_n 0.00457111f $X=2.9 $Y=1.885 $X2=0
+ $Y2=0
cc_369 N_A_27_112#_c_451_n N_VPWR_c_998_n 7.90126e-19 $X=2.66 $Y=2.565 $X2=0
+ $Y2=0
cc_370 N_A_27_112#_c_409_n N_VPWR_c_1002_n 0.0159324f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_371 N_A_27_112#_c_399_n N_VPWR_c_987_n 0.00897215f $X=2.9 $Y=1.885 $X2=0
+ $Y2=0
cc_372 N_A_27_112#_c_407_n N_VPWR_c_987_n 0.0196082f $X=1.795 $Y=2.735 $X2=0
+ $Y2=0
cc_373 N_A_27_112#_c_429_n N_VPWR_c_987_n 0.00543326f $X=1.155 $Y=2.735 $X2=0
+ $Y2=0
cc_374 N_A_27_112#_c_451_n N_VPWR_c_987_n 0.0161828f $X=2.66 $Y=2.565 $X2=0
+ $Y2=0
cc_375 N_A_27_112#_c_409_n N_VPWR_c_987_n 0.0131546f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_376 N_A_27_112#_c_410_n N_VPWR_c_987_n 0.00542643f $X=1.88 $Y=2.565 $X2=0
+ $Y2=0
cc_377 N_A_27_112#_c_400_n N_VGND_c_1167_n 0.0206999f $X=0.265 $Y=0.91 $X2=0
+ $Y2=0
cc_378 N_A_27_112#_c_400_n N_VGND_c_1176_n 0.00882793f $X=0.265 $Y=0.91 $X2=0
+ $Y2=0
cc_379 N_A_27_112#_M1002_g N_VGND_c_1178_n 0.00384553f $X=2.885 $Y=0.69 $X2=0
+ $Y2=0
cc_380 N_A_27_112#_M1002_g N_VGND_c_1183_n 0.0135587f $X=2.885 $Y=0.69 $X2=0
+ $Y2=0
cc_381 N_A_27_112#_M1002_g N_VGND_c_1187_n 0.00371083f $X=2.885 $Y=0.69 $X2=0
+ $Y2=0
cc_382 N_A_27_112#_c_400_n N_VGND_c_1187_n 0.0115594f $X=0.265 $Y=0.91 $X2=0
+ $Y2=0
cc_383 N_A_363_74#_M1010_g N_A_838_48#_c_605_n 0.0401136f $X=3.875 $Y=0.58 $X2=0
+ $Y2=0
cc_384 N_A_363_74#_M1010_g N_A_838_48#_c_606_n 0.00486351f $X=3.875 $Y=0.58
+ $X2=0 $Y2=0
cc_385 N_A_363_74#_c_505_n N_A_838_48#_c_606_n 2.07695e-19 $X=3.8 $Y=1.225 $X2=0
+ $Y2=0
cc_386 N_A_363_74#_c_507_n N_A_838_48#_c_606_n 3.47742e-19 $X=3.965 $Y=1.39
+ $X2=0 $Y2=0
cc_387 N_A_363_74#_c_508_n N_A_838_48#_c_606_n 0.0246062f $X=3.965 $Y=1.39 $X2=0
+ $Y2=0
cc_388 N_A_363_74#_c_504_n N_A_670_74#_M1001_d 0.00785398f $X=3.715 $Y=0.865
+ $X2=-0.19 $Y2=-0.245
cc_389 N_A_363_74#_M1010_g N_A_670_74#_c_776_n 0.0146888f $X=3.875 $Y=0.58 $X2=0
+ $Y2=0
cc_390 N_A_363_74#_c_504_n N_A_670_74#_c_776_n 0.0324151f $X=3.715 $Y=0.865
+ $X2=0 $Y2=0
cc_391 N_A_363_74#_c_507_n N_A_670_74#_c_776_n 0.00370667f $X=3.965 $Y=1.39
+ $X2=0 $Y2=0
cc_392 N_A_363_74#_c_508_n N_A_670_74#_c_776_n 0.00150024f $X=3.965 $Y=1.39
+ $X2=0 $Y2=0
cc_393 N_A_363_74#_c_510_n N_A_670_74#_c_784_n 0.00522521f $X=3.8 $Y=1.765 $X2=0
+ $Y2=0
cc_394 N_A_363_74#_c_507_n N_A_670_74#_c_784_n 0.0305111f $X=3.965 $Y=1.39 $X2=0
+ $Y2=0
cc_395 N_A_363_74#_c_508_n N_A_670_74#_c_784_n 0.00796518f $X=3.965 $Y=1.39
+ $X2=0 $Y2=0
cc_396 N_A_363_74#_c_510_n N_A_670_74#_c_785_n 0.0140898f $X=3.8 $Y=1.765 $X2=0
+ $Y2=0
cc_397 N_A_363_74#_c_511_n N_A_670_74#_c_785_n 8.84976e-19 $X=3.38 $Y=1.765
+ $X2=0 $Y2=0
cc_398 N_A_363_74#_M1010_g N_A_670_74#_c_777_n 0.00431645f $X=3.875 $Y=0.58
+ $X2=0 $Y2=0
cc_399 N_A_363_74#_c_504_n N_A_670_74#_c_777_n 0.00837739f $X=3.715 $Y=0.865
+ $X2=0 $Y2=0
cc_400 N_A_363_74#_M1010_g N_A_670_74#_c_778_n 0.00117587f $X=3.875 $Y=0.58
+ $X2=0 $Y2=0
cc_401 N_A_363_74#_c_505_n N_A_670_74#_c_778_n 0.00623713f $X=3.8 $Y=1.225 $X2=0
+ $Y2=0
cc_402 N_A_363_74#_c_507_n N_A_670_74#_c_778_n 0.0240592f $X=3.965 $Y=1.39 $X2=0
+ $Y2=0
cc_403 N_A_363_74#_c_508_n N_A_670_74#_c_778_n 0.00405396f $X=3.965 $Y=1.39
+ $X2=0 $Y2=0
cc_404 N_A_363_74#_c_509_n N_A_670_74#_c_797_n 0.0038846f $X=3.29 $Y=1.885 $X2=0
+ $Y2=0
cc_405 N_A_363_74#_c_510_n N_A_670_74#_c_797_n 0.00225716f $X=3.8 $Y=1.765 $X2=0
+ $Y2=0
cc_406 N_A_363_74#_c_509_n N_A_670_74#_c_789_n 0.0061512f $X=3.29 $Y=1.885 $X2=0
+ $Y2=0
cc_407 N_A_363_74#_M1010_g N_A_670_74#_c_780_n 0.00115459f $X=3.875 $Y=0.58
+ $X2=0 $Y2=0
cc_408 N_A_363_74#_c_504_n N_A_670_74#_c_780_n 0.00549096f $X=3.715 $Y=0.865
+ $X2=0 $Y2=0
cc_409 N_A_363_74#_c_505_n N_A_670_74#_c_780_n 0.00800927f $X=3.8 $Y=1.225 $X2=0
+ $Y2=0
cc_410 N_A_363_74#_c_507_n N_A_670_74#_c_780_n 0.00561677f $X=3.965 $Y=1.39
+ $X2=0 $Y2=0
cc_411 N_A_363_74#_c_508_n N_A_670_74#_c_780_n 0.00168154f $X=3.965 $Y=1.39
+ $X2=0 $Y2=0
cc_412 N_A_363_74#_c_509_n N_VPWR_c_998_n 0.00278271f $X=3.29 $Y=1.885 $X2=0
+ $Y2=0
cc_413 N_A_363_74#_c_509_n N_VPWR_c_987_n 0.00354243f $X=3.29 $Y=1.885 $X2=0
+ $Y2=0
cc_414 N_A_363_74#_c_504_n N_VGND_M1019_d 0.0110774f $X=3.715 $Y=0.865 $X2=0
+ $Y2=0
cc_415 N_A_363_74#_c_502_n N_VGND_c_1177_n 0.0145091f $X=1.96 $Y=0.515 $X2=0
+ $Y2=0
cc_416 N_A_363_74#_M1010_g N_VGND_c_1178_n 0.00292999f $X=3.875 $Y=0.58 $X2=0
+ $Y2=0
cc_417 N_A_363_74#_c_502_n N_VGND_c_1183_n 0.0102322f $X=1.96 $Y=0.515 $X2=0
+ $Y2=0
cc_418 N_A_363_74#_c_504_n N_VGND_c_1183_n 0.0353648f $X=3.715 $Y=0.865 $X2=0
+ $Y2=0
cc_419 N_A_363_74#_M1010_g N_VGND_c_1187_n 0.00361394f $X=3.875 $Y=0.58 $X2=0
+ $Y2=0
cc_420 N_A_363_74#_c_502_n N_VGND_c_1187_n 0.0119768f $X=1.96 $Y=0.515 $X2=0
+ $Y2=0
cc_421 N_A_363_74#_c_504_n N_VGND_c_1187_n 0.0238967f $X=3.715 $Y=0.865 $X2=0
+ $Y2=0
cc_422 N_A_363_74#_c_504_n A_592_74# 0.00377716f $X=3.715 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_423 N_A_838_48#_c_606_n N_A_670_74#_c_781_n 0.00489279f $X=4.45 $Y=2.035
+ $X2=0 $Y2=0
cc_424 N_A_838_48#_c_619_n N_A_670_74#_c_781_n 0.0194673f $X=4.465 $Y=2.465
+ $X2=0 $Y2=0
cc_425 N_A_838_48#_c_624_n N_A_670_74#_c_781_n 0.0128279f $X=5.23 $Y=2.2 $X2=0
+ $Y2=0
cc_426 N_A_838_48#_c_614_n N_A_670_74#_c_781_n 0.00111494f $X=5.315 $Y=1.82
+ $X2=0 $Y2=0
cc_427 N_A_838_48#_c_626_n N_A_670_74#_c_781_n 0.0183157f $X=5.475 $Y=2.41 $X2=0
+ $Y2=0
cc_428 N_A_838_48#_c_627_n N_A_670_74#_c_781_n 0.0135904f $X=5.475 $Y=2.815
+ $X2=0 $Y2=0
cc_429 N_A_838_48#_c_612_n N_A_670_74#_M1025_g 0.00674246f $X=4.45 $Y=0.94 $X2=0
+ $Y2=0
cc_430 N_A_838_48#_c_614_n N_A_670_74#_M1025_g 0.0110443f $X=5.315 $Y=1.82 $X2=0
+ $Y2=0
cc_431 N_A_838_48#_c_615_n N_A_670_74#_M1025_g 0.020219f $X=5.04 $Y=0.515 $X2=0
+ $Y2=0
cc_432 N_A_838_48#_c_606_n N_A_670_74#_c_774_n 0.0201372f $X=4.45 $Y=2.035 $X2=0
+ $Y2=0
cc_433 N_A_838_48#_c_624_n N_A_670_74#_c_774_n 0.00373089f $X=5.23 $Y=2.2 $X2=0
+ $Y2=0
cc_434 N_A_838_48#_c_615_n N_A_670_74#_c_774_n 0.006551f $X=5.04 $Y=0.515 $X2=0
+ $Y2=0
cc_435 N_A_838_48#_c_606_n N_A_670_74#_c_775_n 9.42097e-19 $X=4.45 $Y=2.035
+ $X2=0 $Y2=0
cc_436 N_A_838_48#_c_614_n N_A_670_74#_c_775_n 0.011331f $X=5.315 $Y=1.82 $X2=0
+ $Y2=0
cc_437 N_A_838_48#_c_605_n N_A_670_74#_c_776_n 0.00576439f $X=4.265 $Y=0.865
+ $X2=0 $Y2=0
cc_438 N_A_838_48#_c_612_n N_A_670_74#_c_784_n 4.98229e-19 $X=4.45 $Y=0.94 $X2=0
+ $Y2=0
cc_439 N_A_838_48#_c_605_n N_A_670_74#_c_777_n 0.00610868f $X=4.265 $Y=0.865
+ $X2=0 $Y2=0
cc_440 N_A_838_48#_c_612_n N_A_670_74#_c_777_n 7.55125e-19 $X=4.45 $Y=0.94 $X2=0
+ $Y2=0
cc_441 N_A_838_48#_c_615_n N_A_670_74#_c_777_n 0.00484459f $X=5.04 $Y=0.515
+ $X2=0 $Y2=0
cc_442 N_A_838_48#_c_606_n N_A_670_74#_c_778_n 0.0225477f $X=4.45 $Y=2.035 $X2=0
+ $Y2=0
cc_443 N_A_838_48#_c_612_n N_A_670_74#_c_778_n 7.62906e-19 $X=4.45 $Y=0.94 $X2=0
+ $Y2=0
cc_444 N_A_838_48#_c_615_n N_A_670_74#_c_778_n 0.00309878f $X=5.04 $Y=0.515
+ $X2=0 $Y2=0
cc_445 N_A_838_48#_c_606_n N_A_670_74#_c_787_n 0.00716452f $X=4.45 $Y=2.035
+ $X2=0 $Y2=0
cc_446 N_A_838_48#_c_619_n N_A_670_74#_c_787_n 0.00418655f $X=4.465 $Y=2.465
+ $X2=0 $Y2=0
cc_447 N_A_838_48#_c_624_n N_A_670_74#_c_787_n 0.0471087f $X=5.23 $Y=2.2 $X2=0
+ $Y2=0
cc_448 N_A_838_48#_c_614_n N_A_670_74#_c_787_n 0.00880617f $X=5.315 $Y=1.82
+ $X2=0 $Y2=0
cc_449 N_A_838_48#_c_626_n N_A_670_74#_c_787_n 0.00509089f $X=5.475 $Y=2.41
+ $X2=0 $Y2=0
cc_450 N_A_838_48#_c_606_n N_A_670_74#_c_779_n 0.00132925f $X=4.45 $Y=2.035
+ $X2=0 $Y2=0
cc_451 N_A_838_48#_c_614_n N_A_670_74#_c_779_n 0.0257578f $X=5.315 $Y=1.82 $X2=0
+ $Y2=0
cc_452 N_A_838_48#_c_615_n N_A_670_74#_c_779_n 0.0131945f $X=5.04 $Y=0.515 $X2=0
+ $Y2=0
cc_453 N_A_838_48#_c_606_n N_A_670_74#_c_780_n 0.00163074f $X=4.45 $Y=2.035
+ $X2=0 $Y2=0
cc_454 N_A_838_48#_c_612_n N_A_670_74#_c_780_n 0.0161253f $X=4.45 $Y=0.94 $X2=0
+ $Y2=0
cc_455 N_A_838_48#_c_615_n N_A_670_74#_c_780_n 0.00735291f $X=5.04 $Y=0.515
+ $X2=0 $Y2=0
cc_456 N_A_838_48#_c_606_n N_A_670_74#_c_790_n 0.0059317f $X=4.45 $Y=2.035 $X2=0
+ $Y2=0
cc_457 N_A_838_48#_c_624_n N_A_670_74#_c_790_n 0.00753145f $X=5.23 $Y=2.2 $X2=0
+ $Y2=0
cc_458 N_A_838_48#_M1012_g N_RESET_B_c_882_n 0.013193f $X=6.235 $Y=0.74
+ $X2=-0.19 $Y2=-0.245
cc_459 N_A_838_48#_c_614_n N_RESET_B_c_882_n 0.00111087f $X=5.315 $Y=1.82
+ $X2=-0.19 $Y2=-0.245
cc_460 N_A_838_48#_c_615_n N_RESET_B_c_882_n 0.00906715f $X=5.04 $Y=0.515
+ $X2=-0.19 $Y2=-0.245
cc_461 N_A_838_48#_c_607_n N_RESET_B_c_883_n 0.00886509f $X=6.2 $Y=1.675 $X2=0
+ $Y2=0
cc_462 N_A_838_48#_c_621_n N_RESET_B_c_883_n 0.036562f $X=6.2 $Y=1.765 $X2=0
+ $Y2=0
cc_463 N_A_838_48#_M1012_g N_RESET_B_c_883_n 0.00440952f $X=6.235 $Y=0.74 $X2=0
+ $Y2=0
cc_464 N_A_838_48#_c_613_n N_RESET_B_c_883_n 0.0149211f $X=6.21 $Y=1.395 $X2=0
+ $Y2=0
cc_465 N_A_838_48#_c_614_n N_RESET_B_c_883_n 0.00532382f $X=5.315 $Y=1.82 $X2=0
+ $Y2=0
cc_466 N_A_838_48#_c_626_n N_RESET_B_c_883_n 0.0106712f $X=5.475 $Y=2.41 $X2=0
+ $Y2=0
cc_467 N_A_838_48#_c_627_n N_RESET_B_c_883_n 0.00765005f $X=5.475 $Y=2.815 $X2=0
+ $Y2=0
cc_468 N_A_838_48#_c_685_p N_RESET_B_c_883_n 0.0183068f $X=6.785 $Y=2.325 $X2=0
+ $Y2=0
cc_469 N_A_838_48#_c_607_n RESET_B 0.002008f $X=6.2 $Y=1.675 $X2=0 $Y2=0
cc_470 N_A_838_48#_M1012_g RESET_B 0.00116016f $X=6.235 $Y=0.74 $X2=0 $Y2=0
cc_471 N_A_838_48#_c_613_n RESET_B 0.00368677f $X=6.21 $Y=1.395 $X2=0 $Y2=0
cc_472 N_A_838_48#_c_614_n RESET_B 0.0288549f $X=5.315 $Y=1.82 $X2=0 $Y2=0
cc_473 N_A_838_48#_c_626_n RESET_B 0.00414357f $X=5.475 $Y=2.41 $X2=0 $Y2=0
cc_474 N_A_838_48#_M1011_g N_A_1446_368#_c_923_n 0.00380849f $X=7.165 $Y=0.69
+ $X2=0 $Y2=0
cc_475 N_A_838_48#_c_617_n N_A_1446_368#_c_923_n 0.00904455f $X=7.155 $Y=1.542
+ $X2=0 $Y2=0
cc_476 N_A_838_48#_M1027_g N_A_1446_368#_c_925_n 7.6339e-19 $X=6.665 $Y=0.74
+ $X2=0 $Y2=0
cc_477 N_A_838_48#_M1011_g N_A_1446_368#_c_925_n 0.015226f $X=7.165 $Y=0.69
+ $X2=0 $Y2=0
cc_478 N_A_838_48#_c_622_n N_A_1446_368#_c_926_n 8.65463e-19 $X=6.65 $Y=1.765
+ $X2=0 $Y2=0
cc_479 N_A_838_48#_c_623_n N_A_1446_368#_c_926_n 0.01541f $X=7.155 $Y=1.765
+ $X2=0 $Y2=0
cc_480 N_A_838_48#_c_685_p N_A_1446_368#_c_926_n 0.010126f $X=6.785 $Y=2.325
+ $X2=0 $Y2=0
cc_481 N_A_838_48#_c_616_n N_A_1446_368#_c_926_n 0.0369366f $X=6.79 $Y=1.485
+ $X2=0 $Y2=0
cc_482 N_A_838_48#_c_617_n N_A_1446_368#_c_926_n 0.00825057f $X=7.155 $Y=1.542
+ $X2=0 $Y2=0
cc_483 N_A_838_48#_M1027_g N_A_1446_368#_c_941_n 4.64054e-19 $X=6.665 $Y=0.74
+ $X2=0 $Y2=0
cc_484 N_A_838_48#_M1011_g N_A_1446_368#_c_941_n 0.00336549f $X=7.165 $Y=0.69
+ $X2=0 $Y2=0
cc_485 N_A_838_48#_c_616_n N_A_1446_368#_c_941_n 0.0130535f $X=6.79 $Y=1.485
+ $X2=0 $Y2=0
cc_486 N_A_838_48#_c_617_n N_A_1446_368#_c_941_n 0.00799528f $X=7.155 $Y=1.542
+ $X2=0 $Y2=0
cc_487 N_A_838_48#_c_624_n N_VPWR_M1021_d 0.00649248f $X=5.23 $Y=2.2 $X2=0 $Y2=0
cc_488 N_A_838_48#_c_685_p N_VPWR_M1017_d 0.0101418f $X=6.785 $Y=2.325 $X2=0
+ $Y2=0
cc_489 N_A_838_48#_c_685_p N_VPWR_M1023_d 0.00406293f $X=6.785 $Y=2.325 $X2=0
+ $Y2=0
cc_490 N_A_838_48#_c_628_n N_VPWR_M1023_d 0.0102704f $X=6.87 $Y=2.24 $X2=0 $Y2=0
cc_491 N_A_838_48#_c_621_n N_VPWR_c_990_n 0.0110436f $X=6.2 $Y=1.765 $X2=0 $Y2=0
cc_492 N_A_838_48#_c_622_n N_VPWR_c_990_n 0.0015077f $X=6.65 $Y=1.765 $X2=0
+ $Y2=0
cc_493 N_A_838_48#_c_627_n N_VPWR_c_990_n 0.0157994f $X=5.475 $Y=2.815 $X2=0
+ $Y2=0
cc_494 N_A_838_48#_c_685_p N_VPWR_c_990_n 0.0202671f $X=6.785 $Y=2.325 $X2=0
+ $Y2=0
cc_495 N_A_838_48#_c_621_n N_VPWR_c_991_n 0.0015077f $X=6.2 $Y=1.765 $X2=0 $Y2=0
cc_496 N_A_838_48#_c_622_n N_VPWR_c_991_n 0.0130128f $X=6.65 $Y=1.765 $X2=0
+ $Y2=0
cc_497 N_A_838_48#_c_623_n N_VPWR_c_991_n 0.00470488f $X=7.155 $Y=1.765 $X2=0
+ $Y2=0
cc_498 N_A_838_48#_c_685_p N_VPWR_c_991_n 0.0163963f $X=6.785 $Y=2.325 $X2=0
+ $Y2=0
cc_499 N_A_838_48#_c_623_n N_VPWR_c_992_n 0.00441756f $X=7.155 $Y=1.765 $X2=0
+ $Y2=0
cc_500 N_A_838_48#_c_621_n N_VPWR_c_995_n 0.00413917f $X=6.2 $Y=1.765 $X2=0
+ $Y2=0
cc_501 N_A_838_48#_c_622_n N_VPWR_c_995_n 0.00413917f $X=6.65 $Y=1.765 $X2=0
+ $Y2=0
cc_502 N_A_838_48#_c_619_n N_VPWR_c_998_n 0.00415318f $X=4.465 $Y=2.465 $X2=0
+ $Y2=0
cc_503 N_A_838_48#_c_627_n N_VPWR_c_999_n 0.0145819f $X=5.475 $Y=2.815 $X2=0
+ $Y2=0
cc_504 N_A_838_48#_c_623_n N_VPWR_c_1000_n 0.00481995f $X=7.155 $Y=1.765 $X2=0
+ $Y2=0
cc_505 N_A_838_48#_c_619_n N_VPWR_c_1004_n 0.0185817f $X=4.465 $Y=2.465 $X2=0
+ $Y2=0
cc_506 N_A_838_48#_c_624_n N_VPWR_c_1004_n 0.0305033f $X=5.23 $Y=2.2 $X2=0 $Y2=0
cc_507 N_A_838_48#_c_627_n N_VPWR_c_1004_n 0.0132508f $X=5.475 $Y=2.815 $X2=0
+ $Y2=0
cc_508 N_A_838_48#_c_619_n N_VPWR_c_987_n 0.00856988f $X=4.465 $Y=2.465 $X2=0
+ $Y2=0
cc_509 N_A_838_48#_c_621_n N_VPWR_c_987_n 0.00817726f $X=6.2 $Y=1.765 $X2=0
+ $Y2=0
cc_510 N_A_838_48#_c_622_n N_VPWR_c_987_n 0.00817726f $X=6.65 $Y=1.765 $X2=0
+ $Y2=0
cc_511 N_A_838_48#_c_623_n N_VPWR_c_987_n 0.00508379f $X=7.155 $Y=1.765 $X2=0
+ $Y2=0
cc_512 N_A_838_48#_c_627_n N_VPWR_c_987_n 0.0120273f $X=5.475 $Y=2.815 $X2=0
+ $Y2=0
cc_513 N_A_838_48#_c_685_p N_Q_M1004_s 0.00907415f $X=6.785 $Y=2.325 $X2=0 $Y2=0
cc_514 N_A_838_48#_c_621_n N_Q_c_1111_n 0.00619743f $X=6.2 $Y=1.765 $X2=0 $Y2=0
cc_515 N_A_838_48#_c_609_n N_Q_c_1111_n 4.44921e-19 $X=6.56 $Y=1.395 $X2=0 $Y2=0
cc_516 N_A_838_48#_c_622_n N_Q_c_1111_n 0.00360318f $X=6.65 $Y=1.765 $X2=0 $Y2=0
cc_517 N_A_838_48#_c_626_n N_Q_c_1111_n 0.00655226f $X=5.475 $Y=2.41 $X2=0 $Y2=0
cc_518 N_A_838_48#_c_685_p N_Q_c_1111_n 0.0166367f $X=6.785 $Y=2.325 $X2=0 $Y2=0
cc_519 N_A_838_48#_c_628_n N_Q_c_1111_n 0.0166315f $X=6.87 $Y=2.24 $X2=0 $Y2=0
cc_520 N_A_838_48#_c_617_n N_Q_c_1111_n 7.34584e-19 $X=7.155 $Y=1.542 $X2=0
+ $Y2=0
cc_521 N_A_838_48#_c_607_n N_Q_c_1109_n 0.00462704f $X=6.2 $Y=1.675 $X2=0 $Y2=0
cc_522 N_A_838_48#_c_621_n N_Q_c_1109_n 0.00396515f $X=6.2 $Y=1.765 $X2=0 $Y2=0
cc_523 N_A_838_48#_M1012_g N_Q_c_1109_n 0.00410571f $X=6.235 $Y=0.74 $X2=0 $Y2=0
cc_524 N_A_838_48#_c_609_n N_Q_c_1109_n 0.00703306f $X=6.56 $Y=1.395 $X2=0 $Y2=0
cc_525 N_A_838_48#_M1027_g N_Q_c_1109_n 0.00301876f $X=6.665 $Y=0.74 $X2=0 $Y2=0
cc_526 N_A_838_48#_c_613_n N_Q_c_1109_n 0.00224562f $X=6.21 $Y=1.395 $X2=0 $Y2=0
cc_527 N_A_838_48#_c_628_n N_Q_c_1109_n 0.00566705f $X=6.87 $Y=2.24 $X2=0 $Y2=0
cc_528 N_A_838_48#_c_616_n N_Q_c_1109_n 0.0242389f $X=6.79 $Y=1.485 $X2=0 $Y2=0
cc_529 N_A_838_48#_c_617_n N_Q_c_1109_n 0.00234865f $X=7.155 $Y=1.542 $X2=0
+ $Y2=0
cc_530 N_A_838_48#_M1012_g Q 0.00628447f $X=6.235 $Y=0.74 $X2=0 $Y2=0
cc_531 N_A_838_48#_c_609_n Q 0.00186821f $X=6.56 $Y=1.395 $X2=0 $Y2=0
cc_532 N_A_838_48#_M1027_g Q 0.00629995f $X=6.665 $Y=0.74 $X2=0 $Y2=0
cc_533 N_A_838_48#_M1011_g Q 3.11727e-19 $X=7.165 $Y=0.69 $X2=0 $Y2=0
cc_534 N_A_838_48#_c_605_n N_VGND_c_1168_n 0.00506215f $X=4.265 $Y=0.865 $X2=0
+ $Y2=0
cc_535 N_A_838_48#_c_612_n N_VGND_c_1168_n 0.00478042f $X=4.45 $Y=0.94 $X2=0
+ $Y2=0
cc_536 N_A_838_48#_c_615_n N_VGND_c_1168_n 0.0249954f $X=5.04 $Y=0.515 $X2=0
+ $Y2=0
cc_537 N_A_838_48#_M1012_g N_VGND_c_1169_n 0.016125f $X=6.235 $Y=0.74 $X2=0
+ $Y2=0
cc_538 N_A_838_48#_c_615_n N_VGND_c_1169_n 0.0348801f $X=5.04 $Y=0.515 $X2=0
+ $Y2=0
cc_539 N_A_838_48#_M1027_g N_VGND_c_1170_n 0.00348163f $X=6.665 $Y=0.74 $X2=0
+ $Y2=0
cc_540 N_A_838_48#_M1011_g N_VGND_c_1170_n 0.00679159f $X=7.165 $Y=0.69 $X2=0
+ $Y2=0
cc_541 N_A_838_48#_c_616_n N_VGND_c_1170_n 0.00991353f $X=6.79 $Y=1.485 $X2=0
+ $Y2=0
cc_542 N_A_838_48#_c_617_n N_VGND_c_1170_n 0.00276433f $X=7.155 $Y=1.542 $X2=0
+ $Y2=0
cc_543 N_A_838_48#_M1011_g N_VGND_c_1171_n 0.00393759f $X=7.165 $Y=0.69 $X2=0
+ $Y2=0
cc_544 N_A_838_48#_c_615_n N_VGND_c_1174_n 0.0228884f $X=5.04 $Y=0.515 $X2=0
+ $Y2=0
cc_545 N_A_838_48#_c_605_n N_VGND_c_1178_n 0.00422124f $X=4.265 $Y=0.865 $X2=0
+ $Y2=0
cc_546 N_A_838_48#_M1012_g N_VGND_c_1179_n 0.00461464f $X=6.235 $Y=0.74 $X2=0
+ $Y2=0
cc_547 N_A_838_48#_M1027_g N_VGND_c_1179_n 0.00461464f $X=6.665 $Y=0.74 $X2=0
+ $Y2=0
cc_548 N_A_838_48#_M1011_g N_VGND_c_1180_n 0.00434272f $X=7.165 $Y=0.69 $X2=0
+ $Y2=0
cc_549 N_A_838_48#_c_605_n N_VGND_c_1187_n 0.00784892f $X=4.265 $Y=0.865 $X2=0
+ $Y2=0
cc_550 N_A_838_48#_M1012_g N_VGND_c_1187_n 0.00836717f $X=6.235 $Y=0.74 $X2=0
+ $Y2=0
cc_551 N_A_838_48#_M1027_g N_VGND_c_1187_n 0.0083477f $X=6.665 $Y=0.74 $X2=0
+ $Y2=0
cc_552 N_A_838_48#_M1011_g N_VGND_c_1187_n 0.00825717f $X=7.165 $Y=0.69 $X2=0
+ $Y2=0
cc_553 N_A_838_48#_c_612_n N_VGND_c_1187_n 0.00123274f $X=4.45 $Y=0.94 $X2=0
+ $Y2=0
cc_554 N_A_838_48#_c_615_n N_VGND_c_1187_n 0.0185926f $X=5.04 $Y=0.515 $X2=0
+ $Y2=0
cc_555 N_A_838_48#_c_615_n A_1066_74# 0.00827328f $X=5.04 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_556 N_A_670_74#_M1025_g N_RESET_B_c_882_n 0.0336962f $X=5.255 $Y=0.74
+ $X2=-0.19 $Y2=-0.245
cc_557 N_A_670_74#_c_781_n N_RESET_B_c_883_n 0.0095821f $X=5.24 $Y=1.765 $X2=0
+ $Y2=0
cc_558 N_A_670_74#_c_775_n N_RESET_B_c_883_n 0.0426444f $X=5.24 $Y=1.557 $X2=0
+ $Y2=0
cc_559 N_A_670_74#_M1025_g RESET_B 4.04852e-19 $X=5.255 $Y=0.74 $X2=0 $Y2=0
cc_560 N_A_670_74#_c_787_n N_VPWR_M1021_d 0.00222541f $X=4.735 $Y=1.795 $X2=0
+ $Y2=0
cc_561 N_A_670_74#_c_781_n N_VPWR_c_999_n 0.00456932f $X=5.24 $Y=1.765 $X2=0
+ $Y2=0
cc_562 N_A_670_74#_c_781_n N_VPWR_c_1004_n 0.00523396f $X=5.24 $Y=1.765 $X2=0
+ $Y2=0
cc_563 N_A_670_74#_c_781_n N_VPWR_c_987_n 0.00892062f $X=5.24 $Y=1.765 $X2=0
+ $Y2=0
cc_564 N_A_670_74#_M1025_g N_VGND_c_1168_n 0.0032926f $X=5.255 $Y=0.74 $X2=0
+ $Y2=0
cc_565 N_A_670_74#_c_776_n N_VGND_c_1168_n 0.0108916f $X=4.055 $Y=0.485 $X2=0
+ $Y2=0
cc_566 N_A_670_74#_c_780_n N_VGND_c_1168_n 0.005796f $X=4.385 $Y=0.97 $X2=0
+ $Y2=0
cc_567 N_A_670_74#_M1025_g N_VGND_c_1169_n 0.00119755f $X=5.255 $Y=0.74 $X2=0
+ $Y2=0
cc_568 N_A_670_74#_M1025_g N_VGND_c_1174_n 0.00291513f $X=5.255 $Y=0.74 $X2=0
+ $Y2=0
cc_569 N_A_670_74#_c_776_n N_VGND_c_1178_n 0.0356621f $X=4.055 $Y=0.485 $X2=0
+ $Y2=0
cc_570 N_A_670_74#_c_776_n N_VGND_c_1183_n 0.00832678f $X=4.055 $Y=0.485 $X2=0
+ $Y2=0
cc_571 N_A_670_74#_M1025_g N_VGND_c_1187_n 0.00363725f $X=5.255 $Y=0.74 $X2=0
+ $Y2=0
cc_572 N_A_670_74#_c_776_n N_VGND_c_1187_n 0.0310952f $X=4.055 $Y=0.485 $X2=0
+ $Y2=0
cc_573 N_A_670_74#_c_776_n A_790_74# 8.31311e-19 $X=4.055 $Y=0.485 $X2=-0.19
+ $Y2=-0.245
cc_574 N_A_670_74#_c_777_n A_790_74# 0.00197162f $X=4.14 $Y=0.885 $X2=-0.19
+ $Y2=-0.245
cc_575 N_RESET_B_c_883_n N_VPWR_c_990_n 0.00393828f $X=5.7 $Y=1.765 $X2=0 $Y2=0
cc_576 N_RESET_B_c_883_n N_VPWR_c_999_n 0.00445602f $X=5.7 $Y=1.765 $X2=0 $Y2=0
cc_577 N_RESET_B_c_883_n N_VPWR_c_987_n 0.00857605f $X=5.7 $Y=1.765 $X2=0 $Y2=0
cc_578 N_RESET_B_c_883_n N_Q_c_1111_n 7.58301e-19 $X=5.7 $Y=1.765 $X2=0 $Y2=0
cc_579 N_RESET_B_c_883_n N_Q_c_1109_n 0.00119389f $X=5.7 $Y=1.765 $X2=0 $Y2=0
cc_580 RESET_B N_Q_c_1109_n 0.028017f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_581 N_RESET_B_c_882_n Q 5.33099e-19 $X=5.645 $Y=1.22 $X2=0 $Y2=0
cc_582 N_RESET_B_c_882_n N_VGND_c_1169_n 0.0130957f $X=5.645 $Y=1.22 $X2=0 $Y2=0
cc_583 N_RESET_B_c_883_n N_VGND_c_1169_n 0.00111502f $X=5.7 $Y=1.765 $X2=0 $Y2=0
cc_584 RESET_B N_VGND_c_1169_n 0.025907f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_585 N_RESET_B_c_882_n N_VGND_c_1174_n 0.00383152f $X=5.645 $Y=1.22 $X2=0
+ $Y2=0
cc_586 N_RESET_B_c_882_n N_VGND_c_1187_n 0.0075725f $X=5.645 $Y=1.22 $X2=0 $Y2=0
cc_587 N_A_1446_368#_c_926_n N_VPWR_c_991_n 0.0110392f $X=7.38 $Y=1.985 $X2=0
+ $Y2=0
cc_588 N_A_1446_368#_c_919_n N_VPWR_c_992_n 0.0100916f $X=8.165 $Y=1.765 $X2=0
+ $Y2=0
cc_589 N_A_1446_368#_c_923_n N_VPWR_c_992_n 0.00546342f $X=8.075 $Y=1.385 $X2=0
+ $Y2=0
cc_590 N_A_1446_368#_c_926_n N_VPWR_c_992_n 0.0686723f $X=7.38 $Y=1.985 $X2=0
+ $Y2=0
cc_591 N_A_1446_368#_c_927_n N_VPWR_c_992_n 0.0148177f $X=8.065 $Y=1.385 $X2=0
+ $Y2=0
cc_592 N_A_1446_368#_c_930_n N_VPWR_c_994_n 0.00972643f $X=8.615 $Y=1.765 $X2=0
+ $Y2=0
cc_593 N_A_1446_368#_c_926_n N_VPWR_c_1000_n 0.0097982f $X=7.38 $Y=1.985 $X2=0
+ $Y2=0
cc_594 N_A_1446_368#_c_919_n N_VPWR_c_1001_n 0.00445602f $X=8.165 $Y=1.765 $X2=0
+ $Y2=0
cc_595 N_A_1446_368#_c_930_n N_VPWR_c_1001_n 0.00422942f $X=8.615 $Y=1.765 $X2=0
+ $Y2=0
cc_596 N_A_1446_368#_c_919_n N_VPWR_c_987_n 0.00862391f $X=8.165 $Y=1.765 $X2=0
+ $Y2=0
cc_597 N_A_1446_368#_c_930_n N_VPWR_c_987_n 0.0078771f $X=8.615 $Y=1.765 $X2=0
+ $Y2=0
cc_598 N_A_1446_368#_c_926_n N_VPWR_c_987_n 0.0111907f $X=7.38 $Y=1.985 $X2=0
+ $Y2=0
cc_599 N_A_1446_368#_c_925_n Q 0.00211465f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_600 N_A_1446_368#_c_918_n N_Q_N_c_1145_n 0.00315047f $X=8.155 $Y=1.22 $X2=0
+ $Y2=0
cc_601 N_A_1446_368#_c_920_n N_Q_N_c_1145_n 0.0032084f $X=8.525 $Y=1.295 $X2=0
+ $Y2=0
cc_602 N_A_1446_368#_c_922_n N_Q_N_c_1145_n 0.00289446f $X=8.625 $Y=1.22 $X2=0
+ $Y2=0
cc_603 N_A_1446_368#_c_927_n N_Q_N_c_1145_n 0.00175142f $X=8.065 $Y=1.385 $X2=0
+ $Y2=0
cc_604 N_A_1446_368#_c_919_n Q_N 0.00328275f $X=8.165 $Y=1.765 $X2=0 $Y2=0
cc_605 N_A_1446_368#_c_920_n Q_N 0.00260132f $X=8.525 $Y=1.295 $X2=0 $Y2=0
cc_606 N_A_1446_368#_c_930_n Q_N 0.00227136f $X=8.615 $Y=1.765 $X2=0 $Y2=0
cc_607 N_A_1446_368#_c_919_n Q_N 0.0115887f $X=8.165 $Y=1.765 $X2=0 $Y2=0
cc_608 N_A_1446_368#_c_930_n Q_N 0.0126237f $X=8.615 $Y=1.765 $X2=0 $Y2=0
cc_609 N_A_1446_368#_c_918_n N_Q_N_c_1141_n 0.0033377f $X=8.155 $Y=1.22 $X2=0
+ $Y2=0
cc_610 N_A_1446_368#_c_919_n N_Q_N_c_1141_n 0.00626192f $X=8.165 $Y=1.765 $X2=0
+ $Y2=0
cc_611 N_A_1446_368#_c_920_n N_Q_N_c_1141_n 0.0053896f $X=8.525 $Y=1.295 $X2=0
+ $Y2=0
cc_612 N_A_1446_368#_c_921_n N_Q_N_c_1141_n 0.0105594f $X=8.615 $Y=1.675 $X2=0
+ $Y2=0
cc_613 N_A_1446_368#_c_930_n N_Q_N_c_1141_n 0.00738107f $X=8.615 $Y=1.765 $X2=0
+ $Y2=0
cc_614 N_A_1446_368#_c_922_n N_Q_N_c_1141_n 0.00540128f $X=8.625 $Y=1.22 $X2=0
+ $Y2=0
cc_615 N_A_1446_368#_c_924_n N_Q_N_c_1141_n 0.010885f $X=8.525 $Y=1.22 $X2=0
+ $Y2=0
cc_616 N_A_1446_368#_c_927_n N_Q_N_c_1141_n 0.0250802f $X=8.065 $Y=1.385 $X2=0
+ $Y2=0
cc_617 N_A_1446_368#_c_925_n N_VGND_c_1170_n 0.0285932f $X=7.38 $Y=0.515 $X2=0
+ $Y2=0
cc_618 N_A_1446_368#_c_918_n N_VGND_c_1171_n 0.00531218f $X=8.155 $Y=1.22 $X2=0
+ $Y2=0
cc_619 N_A_1446_368#_c_923_n N_VGND_c_1171_n 0.00597676f $X=8.075 $Y=1.385 $X2=0
+ $Y2=0
cc_620 N_A_1446_368#_c_925_n N_VGND_c_1171_n 0.0463564f $X=7.38 $Y=0.515 $X2=0
+ $Y2=0
cc_621 N_A_1446_368#_c_927_n N_VGND_c_1171_n 0.0208454f $X=8.065 $Y=1.385 $X2=0
+ $Y2=0
cc_622 N_A_1446_368#_c_922_n N_VGND_c_1173_n 0.00663052f $X=8.625 $Y=1.22 $X2=0
+ $Y2=0
cc_623 N_A_1446_368#_c_925_n N_VGND_c_1180_n 0.0145639f $X=7.38 $Y=0.515 $X2=0
+ $Y2=0
cc_624 N_A_1446_368#_c_918_n N_VGND_c_1181_n 0.00461464f $X=8.155 $Y=1.22 $X2=0
+ $Y2=0
cc_625 N_A_1446_368#_c_922_n N_VGND_c_1181_n 0.00461464f $X=8.625 $Y=1.22 $X2=0
+ $Y2=0
cc_626 N_A_1446_368#_c_918_n N_VGND_c_1187_n 0.00913494f $X=8.155 $Y=1.22 $X2=0
+ $Y2=0
cc_627 N_A_1446_368#_c_922_n N_VGND_c_1187_n 0.00912153f $X=8.625 $Y=1.22 $X2=0
+ $Y2=0
cc_628 N_A_1446_368#_c_925_n N_VGND_c_1187_n 0.0119984f $X=7.38 $Y=0.515 $X2=0
+ $Y2=0
cc_629 N_VPWR_c_992_n Q_N 0.0781509f $X=7.94 $Y=1.985 $X2=0 $Y2=0
cc_630 N_VPWR_c_994_n Q_N 0.0847451f $X=8.84 $Y=1.985 $X2=0 $Y2=0
cc_631 N_VPWR_c_1001_n Q_N 0.0153846f $X=8.755 $Y=3.33 $X2=0 $Y2=0
cc_632 N_VPWR_c_987_n Q_N 0.0126213f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_633 Q N_VGND_c_1169_n 0.0134502f $X=6.395 $Y=0.84 $X2=0 $Y2=0
cc_634 Q N_VGND_c_1187_n 0.0129173f $X=6.395 $Y=0.84 $X2=0 $Y2=0
cc_635 N_Q_N_c_1141_n N_VGND_c_1173_n 0.00347369f $X=8.4 $Y=1.82 $X2=0 $Y2=0
