* File: sky130_fd_sc_ls__dlxbn_1.spice
* Created: Fri Aug 28 13:19:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dlxbn_1.pex.spice"
.subckt sky130_fd_sc_ls__dlxbn_1  VNB VPB D GATE_N VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_D_M1017_g N_A_27_120#_M1017_s VNB NSHORT L=0.15 W=0.55
+ AD=0.161184 AS=0.15675 PD=1.20233 PS=1.67 NRD=51.936 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1001 N_A_232_82#_M1001_d N_GATE_N_M1001_g N_VGND_M1017_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.216866 PD=2.05 PS=1.61767 NRD=0 NRS=38.604 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_232_82#_M1007_g N_A_343_80#_M1007_s VNB NSHORT L=0.15
+ W=0.74 AD=0.193727 AS=0.3182 PD=1.49072 PS=2.34 NRD=33.528 NRS=1.62 M=1
+ R=4.93333 SA=75000.4 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1013 A_575_79# N_A_27_120#_M1013_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.167548 PD=0.88 PS=1.28928 NRD=12.18 NRS=15.936 M=1 R=4.26667
+ SA=75000.9 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1012 N_A_653_79#_M1012_d N_A_232_82#_M1012_g A_575_79# VNB NSHORT L=0.15
+ W=0.64 AD=0.247487 AS=0.0768 PD=1.79321 PS=0.88 NRD=18.744 NRS=12.18 M=1
+ R=4.26667 SA=75001.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1010 A_852_123# N_A_343_80#_M1010_g N_A_653_79#_M1012_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.162413 PD=0.66 PS=1.17679 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75002.3 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_863_294#_M1004_g A_852_123# VNB NSHORT L=0.15 W=0.42
+ AD=0.101262 AS=0.0504 PD=0.84 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75002.7 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1002 N_A_863_294#_M1002_d N_A_653_79#_M1002_g N_VGND_M1004_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2183 AS=0.178413 PD=2.07 PS=1.48 NRD=1.62 NRS=9.72 M=1 R=4.93333
+ SA=75002 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A_863_294#_M1008_g N_Q_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.140829 AS=0.2109 PD=1.26202 PS=2.05 NRD=7.296 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_A_1347_424#_M1016_d N_A_863_294#_M1016_g N_VGND_M1008_d VNB NSHORT
+ L=0.15 W=0.55 AD=0.15675 AS=0.104671 PD=1.67 PS=0.937984 NRD=0 NRS=7.632 M=1
+ R=3.66667 SA=75000.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1005 N_Q_N_M1005_d N_A_1347_424#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2072 AS=0.2109 PD=2.04 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_VPWR_M1006_d N_D_M1006_g N_A_27_120#_M1006_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.147 AS=0.294 PD=1.19 PS=2.38 NRD=2.3443 NRS=18.7544 M=1 R=5.6 SA=75000.3
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1011 N_A_232_82#_M1011_d N_GATE_N_M1011_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.147 PD=2.27 PS=1.19 NRD=2.3443 NRS=14.0658 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1018 N_VPWR_M1018_d N_A_232_82#_M1018_g N_A_343_80#_M1018_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.173752 AS=0.2478 PD=1.2737 PS=2.27 NRD=23.443 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1003 A_571_392# N_A_27_120#_M1003_g N_VPWR_M1018_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.206848 PD=1.27 PS=1.5163 NRD=15.7403 NRS=3.9203 M=1 R=6.66667
+ SA=75000.7 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1021 N_A_653_79#_M1021_d N_A_343_80#_M1021_g A_571_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.285704 AS=0.135 PD=2.25352 PS=1.27 NRD=22.6353 NRS=15.7403 M=1 R=6.66667
+ SA=75001.1 SB=75001 A=0.15 P=2.3 MULT=1
MM1000 A_805_392# N_A_232_82#_M1000_g N_A_653_79#_M1021_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.07035 AS=0.119996 PD=0.755 PS=0.946479 NRD=52.7566 NRS=96.136 M=1
+ R=2.8 SA=75001.9 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1015 N_VPWR_M1015_d N_A_863_294#_M1015_g A_805_392# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.121364 AS=0.07035 PD=0.924545 PS=0.755 NRD=46.886 NRS=52.7566 M=1 R=2.8
+ SA=75002.4 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1014 N_A_863_294#_M1014_d N_A_653_79#_M1014_g N_VPWR_M1015_d VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.3136 AS=0.323636 PD=2.8 PS=2.46545 NRD=1.7533 NRS=18.0255
+ M=1 R=7.46667 SA=75001.3 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1019 N_VPWR_M1019_d N_A_863_294#_M1019_g N_Q_M1019_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2128 AS=0.3136 PD=1.68571 PS=2.8 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1020 N_A_1347_424#_M1020_d N_A_863_294#_M1020_g N_VPWR_M1019_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2478 AS=0.1596 PD=2.27 PS=1.26429 NRD=3.5066 NRS=14.0658
+ M=1 R=5.6 SA=75000.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_Q_N_M1009_d N_A_1347_424#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.3136 PD=2.83 PS=2.8 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX22_noxref VNB VPB NWDIODE A=15.97 P=20.96
*
.include "sky130_fd_sc_ls__dlxbn_1.pxi.spice"
*
.ends
*
*
