* File: sky130_fd_sc_ls__or3_4.pex.spice
* Created: Fri Aug 28 13:58:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__OR3_4%A 2 3 5 7 8 10 13 16 17 19 21 25 27 37 41 45
c94 45 0 1.22748e-19 $X=0.24 $Y=1.295
c95 21 0 1.25197e-19 $X=2.905 $Y=1.195
c96 8 0 6.43787e-20 $X=2.89 $Y=1.865
c97 3 0 8.22769e-20 $X=0.505 $Y=1.865
r98 43 45 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.27 $Y=1.28
+ $X2=0.27 $Y2=1.295
r99 37 39 40.5227 $w=4.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.35 $Y=1.465
+ $X2=0.35 $Y2=1.63
r100 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r101 30 37 8.73518 $w=4.9e-07 $l=8e-08 $layer=POLY_cond $X=0.35 $Y=1.385
+ $X2=0.35 $Y2=1.465
r102 30 34 28.3893 $w=4.9e-07 $l=2.6e-07 $layer=POLY_cond $X=0.35 $Y=1.385
+ $X2=0.35 $Y2=1.125
r103 27 43 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=1.195
+ $X2=0.27 $Y2=1.28
r104 27 38 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.27 $Y=1.33
+ $X2=0.27 $Y2=1.465
r105 27 45 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.27 $Y=1.33
+ $X2=0.27 $Y2=1.295
r106 27 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.125 $X2=0.27 $Y2=1.125
r107 25 42 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.92 $Y=1.385
+ $X2=2.92 $Y2=1.55
r108 25 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.92 $Y=1.385
+ $X2=2.92 $Y2=1.22
r109 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.92
+ $Y=1.385 $X2=2.92 $Y2=1.385
r110 21 24 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=2.905 $Y=1.195
+ $X2=2.905 $Y2=1.385
r111 20 27 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=1.195
+ $X2=0.27 $Y2=1.195
r112 19 21 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.755 $Y=1.195
+ $X2=2.905 $Y2=1.195
r113 19 20 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=2.755 $Y=1.195
+ $X2=0.435 $Y2=1.195
r114 17 34 74.249 $w=4.9e-07 $l=6.8e-07 $layer=POLY_cond $X=0.35 $Y=0.445
+ $X2=0.35 $Y2=1.125
r115 16 17 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=0.445 $X2=0.27 $Y2=0.445
r116 14 27 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=1.11
+ $X2=0.27 $Y2=1.195
r117 14 16 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=0.27 $Y=1.11
+ $X2=0.27 $Y2=0.445
r118 13 41 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.93 $Y=0.74
+ $X2=2.93 $Y2=1.22
r119 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.89 $Y=1.865
+ $X2=2.89 $Y2=2.44
r120 7 8 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.89 $Y=1.775 $X2=2.89
+ $Y2=1.865
r121 7 42 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=2.89 $Y=1.775
+ $X2=2.89 $Y2=1.55
r122 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.865
+ $X2=0.505 $Y2=2.44
r123 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.775
+ $X2=0.505 $Y2=1.865
r124 2 39 56.3629 $w=1.8e-07 $l=1.45e-07 $layer=POLY_cond $X=0.505 $Y=1.775
+ $X2=0.505 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_LS__OR3_4%B 1 3 4 6 9 11 12 13 14 24
c59 4 0 1.25197e-19 $X=2.39 $Y=1.865
c60 1 0 1.22748e-19 $X=0.955 $Y=1.865
r61 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=1.615 $X2=2.38 $Y2=1.615
r62 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.615 $X2=0.97 $Y2=1.615
r63 14 24 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.16 $Y=1.615
+ $X2=2.38 $Y2=1.615
r64 13 14 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.615
+ $X2=2.16 $Y2=1.615
r65 12 13 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.68 $Y2=1.615
r66 12 21 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=0.97 $Y2=1.615
r67 11 21 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.97 $Y2=1.615
r68 7 23 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.44 $Y=1.45
+ $X2=2.38 $Y2=1.615
r69 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.44 $Y=1.45 $X2=2.44
+ $Y2=0.74
r70 4 23 52.2586 $w=2.99e-07 $l=2.54951e-07 $layer=POLY_cond $X=2.39 $Y=1.865
+ $X2=2.38 $Y2=1.615
r71 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.39 $Y=1.865
+ $X2=2.39 $Y2=2.44
r72 1 20 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=0.955 $Y=1.865
+ $X2=0.97 $Y2=1.615
r73 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.955 $Y=1.865
+ $X2=0.955 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_LS__OR3_4%C 2 3 5 7 8 10 11 13 17 19 22 23
r57 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.215
+ $Y=0.435 $X2=1.215 $Y2=0.435
r58 19 23 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.215 $Y=0.555
+ $X2=1.215 $Y2=0.435
r59 17 18 9.34914 $w=2.32e-07 $l=4.5e-08 $layer=POLY_cond $X=1.885 $Y=1.345
+ $X2=1.93 $Y2=1.345
r60 16 17 93.4914 $w=2.32e-07 $l=4.5e-07 $layer=POLY_cond $X=1.435 $Y=1.345
+ $X2=1.885 $Y2=1.345
r61 15 22 93.7338 $w=4.45e-07 $l=7.5e-07 $layer=POLY_cond $X=1.272 $Y=1.185
+ $X2=1.272 $Y2=0.435
r62 15 16 33.8647 $w=2.32e-07 $l=2.29454e-07 $layer=POLY_cond $X=1.272 $Y=1.185
+ $X2=1.435 $Y2=1.345
r63 11 18 12.995 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.93 $Y=1.185
+ $X2=1.93 $Y2=1.345
r64 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.93 $Y=1.185
+ $X2=1.93 $Y2=0.74
r65 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.885 $Y=1.865
+ $X2=1.885 $Y2=2.44
r66 7 8 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.885 $Y=1.775 $X2=1.885
+ $Y2=1.865
r67 6 17 8.79421 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=1.885 $Y=1.505
+ $X2=1.885 $Y2=1.345
r68 6 7 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=1.885 $Y=1.505
+ $X2=1.885 $Y2=1.775
r69 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.865
+ $X2=1.435 $Y2=2.44
r70 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.435 $Y=1.775 $X2=1.435
+ $Y2=1.865
r71 1 16 8.79421 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=1.435 $Y=1.505
+ $X2=1.435 $Y2=1.345
r72 1 2 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=1.435 $Y=1.505
+ $X2=1.435 $Y2=1.775
.ends

.subckt PM_SKY130_FD_SC_LS__OR3_4%A_302_388# 1 2 3 10 12 15 19 21 23 24 26 29 31
+ 33 36 40 42 44 45 48 50 53 55 61 67 69 70 79
c166 79 0 1.44954e-19 $X=4.775 $Y=1.532
r167 79 80 1.22646 $w=3.93e-07 $l=1e-08 $layer=POLY_cond $X=4.775 $Y=1.532
+ $X2=4.785 $Y2=1.532
r168 76 77 3.67939 $w=3.93e-07 $l=3e-08 $layer=POLY_cond $X=4.325 $Y=1.532
+ $X2=4.355 $Y2=1.532
r169 75 76 55.1908 $w=3.93e-07 $l=4.5e-07 $layer=POLY_cond $X=3.875 $Y=1.532
+ $X2=4.325 $Y2=1.532
r170 74 75 1.22646 $w=3.93e-07 $l=1e-08 $layer=POLY_cond $X=3.865 $Y=1.532
+ $X2=3.875 $Y2=1.532
r171 71 72 0.613232 $w=3.93e-07 $l=5e-09 $layer=POLY_cond $X=3.425 $Y=1.532
+ $X2=3.43 $Y2=1.532
r172 65 67 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.66 $Y=2.075
+ $X2=1.825 $Y2=2.075
r173 62 79 31.2748 $w=3.93e-07 $l=2.55e-07 $layer=POLY_cond $X=4.52 $Y=1.532
+ $X2=4.775 $Y2=1.532
r174 62 77 20.2366 $w=3.93e-07 $l=1.65e-07 $layer=POLY_cond $X=4.52 $Y=1.532
+ $X2=4.355 $Y2=1.532
r175 61 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.52
+ $Y=1.465 $X2=4.52 $Y2=1.465
r176 59 74 44.7659 $w=3.93e-07 $l=3.65e-07 $layer=POLY_cond $X=3.5 $Y=1.532
+ $X2=3.865 $Y2=1.532
r177 59 72 8.58524 $w=3.93e-07 $l=7e-08 $layer=POLY_cond $X=3.5 $Y=1.532
+ $X2=3.43 $Y2=1.532
r178 58 61 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=3.5 $Y=1.465
+ $X2=4.52 $Y2=1.465
r179 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.5
+ $Y=1.465 $X2=3.5 $Y2=1.465
r180 56 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.395 $Y=1.465
+ $X2=3.31 $Y2=1.465
r181 56 58 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.395 $Y=1.465
+ $X2=3.5 $Y2=1.465
r182 54 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.31 $Y=1.63
+ $X2=3.31 $Y2=1.465
r183 54 55 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.31 $Y=1.63
+ $X2=3.31 $Y2=1.95
r184 53 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.31 $Y=1.3
+ $X2=3.31 $Y2=1.465
r185 52 53 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.31 $Y=0.94
+ $X2=3.31 $Y2=1.3
r186 51 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.88 $Y=0.855
+ $X2=2.715 $Y2=0.855
r187 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.225 $Y=0.855
+ $X2=3.31 $Y2=0.94
r188 50 51 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.225 $Y=0.855
+ $X2=2.88 $Y2=0.855
r189 46 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0.77
+ $X2=2.715 $Y2=0.855
r190 46 48 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.715 $Y=0.77
+ $X2=2.715 $Y2=0.515
r191 44 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=0.855
+ $X2=2.715 $Y2=0.855
r192 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.55 $Y=0.855
+ $X2=1.88 $Y2=0.855
r193 42 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.225 $Y=2.035
+ $X2=3.31 $Y2=1.95
r194 42 67 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=3.225 $Y=2.035
+ $X2=1.825 $Y2=2.035
r195 38 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.715 $Y=0.77
+ $X2=1.88 $Y2=0.855
r196 38 40 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.715 $Y=0.77
+ $X2=1.715 $Y2=0.515
r197 34 80 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.785 $Y=1.3
+ $X2=4.785 $Y2=1.532
r198 34 36 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.785 $Y=1.3
+ $X2=4.785 $Y2=0.74
r199 31 79 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.775 $Y=1.765
+ $X2=4.775 $Y2=1.532
r200 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.775 $Y=1.765
+ $X2=4.775 $Y2=2.4
r201 27 77 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.355 $Y=1.3
+ $X2=4.355 $Y2=1.532
r202 27 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.355 $Y=1.3
+ $X2=4.355 $Y2=0.74
r203 24 76 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.325 $Y=1.765
+ $X2=4.325 $Y2=1.532
r204 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.325 $Y=1.765
+ $X2=4.325 $Y2=2.4
r205 21 75 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.875 $Y=1.765
+ $X2=3.875 $Y2=1.532
r206 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.875 $Y=1.765
+ $X2=3.875 $Y2=2.4
r207 17 74 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.865 $Y=1.3
+ $X2=3.865 $Y2=1.532
r208 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.865 $Y=1.3
+ $X2=3.865 $Y2=0.74
r209 13 72 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.43 $Y=1.3
+ $X2=3.43 $Y2=1.532
r210 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.43 $Y=1.3
+ $X2=3.43 $Y2=0.74
r211 10 71 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.425 $Y=1.765
+ $X2=3.425 $Y2=1.532
r212 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.425 $Y=1.765
+ $X2=3.425 $Y2=2.4
r213 3 65 600 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.94 $X2=1.66 $Y2=2.1
r214 2 69 182 $w=1.7e-07 $l=5.7639e-07 $layer=licon1_NDIFF $count=1 $X=2.515
+ $Y=0.37 $X2=2.715 $Y2=0.855
r215 2 48 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=2.515
+ $Y=0.37 $X2=2.715 $Y2=0.515
r216 1 40 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.57
+ $Y=0.37 $X2=1.715 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR3_4%VPWR 1 2 3 4 13 15 21 25 27 29 31 33 41 46 55
+ 58 62
r70 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r71 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r72 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r73 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 50 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r75 50 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r76 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r77 47 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.06 $Y2=3.33
r78 47 49 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.56 $Y2=3.33
r79 46 61 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=4.915 $Y=3.33
+ $X2=5.097 $Y2=3.33
r80 46 49 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.915 $Y=3.33
+ $X2=4.56 $Y2=3.33
r81 45 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r82 45 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r83 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r84 42 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.2 $Y2=3.33
r85 42 44 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.6 $Y2=3.33
r86 41 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.935 $Y=3.33
+ $X2=4.06 $Y2=3.33
r87 41 44 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.935 $Y=3.33
+ $X2=3.6 $Y2=3.33
r88 37 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r89 36 39 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r90 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r91 34 52 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r92 34 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r93 33 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=3.2 $Y2=3.33
r94 33 39 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=2.64 $Y2=3.33
r95 31 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r96 31 37 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=0.72 $Y2=3.33
r97 31 39 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r98 27 61 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.04 $Y=3.245
+ $X2=5.097 $Y2=3.33
r99 27 29 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=5.04 $Y=3.245
+ $X2=5.04 $Y2=2.305
r100 23 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.06 $Y=3.245
+ $X2=4.06 $Y2=3.33
r101 23 25 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=4.06 $Y=3.245
+ $X2=4.06 $Y2=2.305
r102 19 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=3.245 $X2=3.2
+ $Y2=3.33
r103 19 21 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.2 $Y=3.245
+ $X2=3.2 $Y2=2.455
r104 15 18 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.24 $Y=2.085
+ $X2=0.24 $Y2=2.795
r105 13 52 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r106 13 18 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.795
r107 4 29 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=4.85
+ $Y=1.84 $X2=5 $Y2=2.305
r108 3 25 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=3.95
+ $Y=1.84 $X2=4.1 $Y2=2.305
r109 2 21 300 $w=1.7e-07 $l=6.2149e-07 $layer=licon1_PDIFF $count=2 $X=2.965
+ $Y=1.94 $X2=3.2 $Y2=2.455
r110 1 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.94 $X2=0.28 $Y2=2.795
r111 1 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.94 $X2=0.28 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LS__OR3_4%A_116_388# 1 2 9 13 15 17 19 22
r37 17 24 2.94173 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=2.665 $Y=2.54
+ $X2=2.665 $Y2=2.415
r38 17 19 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.665 $Y=2.54
+ $X2=2.665 $Y2=2.795
r39 16 22 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.815 $Y=2.455
+ $X2=0.69 $Y2=2.455
r40 15 24 4.82444 $w=1.7e-07 $l=1.83916e-07 $layer=LI1_cond $X=2.5 $Y=2.455
+ $X2=2.665 $Y2=2.415
r41 15 16 109.93 $w=1.68e-07 $l=1.685e-06 $layer=LI1_cond $X=2.5 $Y=2.455
+ $X2=0.815 $Y2=2.455
r42 11 22 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.54 $X2=0.69
+ $Y2=2.455
r43 11 13 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.69 $Y=2.54
+ $X2=0.69 $Y2=2.795
r44 7 22 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.37 $X2=0.69
+ $Y2=2.455
r45 7 9 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.69 $Y=2.37 $X2=0.69
+ $Y2=2.115
r46 2 24 600 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.94 $X2=2.665 $Y2=2.455
r47 2 19 600 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.94 $X2=2.665 $Y2=2.795
r48 1 22 600 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.94 $X2=0.73 $Y2=2.455
r49 1 13 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.94 $X2=0.73 $Y2=2.795
r50 1 9 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.94 $X2=0.73 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__OR3_4%A_206_388# 1 2 11
c14 11 0 1.46656e-19 $X=2.135 $Y=2.795
r15 8 11 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=1.195 $Y=2.835
+ $X2=2.135 $Y2=2.835
r16 2 11 600 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.94 $X2=2.135 $Y2=2.795
r17 1 8 600 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.94 $X2=1.195 $Y2=2.795
.ends

.subckt PM_SKY130_FD_SC_LS__OR3_4%X 1 2 3 4 15 19 23 24 25 26 29 35 37 39 41 42
+ 45 46
c83 37 0 1.44954e-19 $X=4.925 $Y=1.045
r84 45 46 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.665
r85 44 46 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.04 $Y=1.8
+ $X2=5.04 $Y2=1.665
r86 43 45 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.04 $Y=1.13
+ $X2=5.04 $Y2=1.295
r87 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=1.885
+ $X2=4.55 $Y2=1.885
r88 39 44 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.925 $Y=1.885
+ $X2=5.04 $Y2=1.8
r89 39 40 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.925 $Y=1.885
+ $X2=4.715 $Y2=1.885
r90 38 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.655 $Y=1.045
+ $X2=4.53 $Y2=1.045
r91 37 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.925 $Y=1.045
+ $X2=5.04 $Y2=1.13
r92 37 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.925 $Y=1.045
+ $X2=4.655 $Y2=1.045
r93 33 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=0.96
+ $X2=4.53 $Y2=1.045
r94 33 35 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=4.53 $Y=0.96
+ $X2=4.53 $Y2=0.515
r95 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.55 $Y=1.985
+ $X2=4.55 $Y2=2.815
r96 27 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=1.97 $X2=4.55
+ $Y2=1.885
r97 27 29 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.55 $Y=1.97
+ $X2=4.55 $Y2=1.985
r98 25 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.385 $Y=1.885
+ $X2=4.55 $Y2=1.885
r99 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.385 $Y=1.885
+ $X2=3.735 $Y2=1.885
r100 23 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.405 $Y=1.045
+ $X2=4.53 $Y2=1.045
r101 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.405 $Y=1.045
+ $X2=3.735 $Y2=1.045
r102 19 21 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.65 $Y=1.985
+ $X2=3.65 $Y2=2.815
r103 17 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.65 $Y=1.97
+ $X2=3.735 $Y2=1.885
r104 17 19 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.65 $Y=1.97
+ $X2=3.65 $Y2=1.985
r105 13 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.65 $Y=0.96
+ $X2=3.735 $Y2=1.045
r106 13 15 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.65 $Y=0.96
+ $X2=3.65 $Y2=0.515
r107 4 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.4
+ $Y=1.84 $X2=4.55 $Y2=2.815
r108 4 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.4
+ $Y=1.84 $X2=4.55 $Y2=1.985
r109 3 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.5
+ $Y=1.84 $X2=3.65 $Y2=2.815
r110 3 19 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.5
+ $Y=1.84 $X2=3.65 $Y2=1.985
r111 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.43
+ $Y=0.37 $X2=4.57 $Y2=0.515
r112 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=3.505
+ $Y=0.37 $X2=3.65 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR3_4%VGND 1 2 3 4 15 17 21 25 27 29 31 33 41 46 52
+ 55 58 62
r74 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r75 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r76 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r77 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r78 50 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r79 50 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r80 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r81 47 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.165 $Y=0 $X2=4.04
+ $Y2=0
r82 47 49 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.165 $Y=0 $X2=4.56
+ $Y2=0
r83 46 61 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5.057
+ $Y2=0
r84 46 49 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=4.56
+ $Y2=0
r85 45 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r86 45 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r87 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r88 42 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.38 $Y=0 $X2=3.215
+ $Y2=0
r89 42 44 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.38 $Y=0 $X2=3.6
+ $Y2=0
r90 41 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.915 $Y=0 $X2=4.04
+ $Y2=0
r91 41 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.915 $Y=0 $X2=3.6
+ $Y2=0
r92 40 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r93 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r94 36 40 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r95 35 39 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r96 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r97 33 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.05 $Y=0 $X2=2.215
+ $Y2=0
r98 33 39 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.05 $Y=0 $X2=1.68
+ $Y2=0
r99 31 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r100 31 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r101 27 61 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5 $Y=0.085
+ $X2=5.057 $Y2=0
r102 27 29 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.61
r103 23 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0
r104 23 25 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.57
r105 19 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=0.085
+ $X2=3.215 $Y2=0
r106 19 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.215 $Y=0.085
+ $X2=3.215 $Y2=0.515
r107 18 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.38 $Y=0 $X2=2.215
+ $Y2=0
r108 17 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=0 $X2=3.215
+ $Y2=0
r109 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.05 $Y=0 $X2=2.38
+ $Y2=0
r110 13 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.215 $Y=0.085
+ $X2=2.215 $Y2=0
r111 13 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.215 $Y=0.085
+ $X2=2.215 $Y2=0.515
r112 4 29 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.37 $X2=5 $Y2=0.61
r113 3 25 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=3.94
+ $Y=0.37 $X2=4.08 $Y2=0.57
r114 2 21 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.005
+ $Y=0.37 $X2=3.215 $Y2=0.515
r115 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.37 $X2=2.215 $Y2=0.515
.ends

