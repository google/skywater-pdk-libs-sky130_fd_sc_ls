* File: sky130_fd_sc_ls__a2bb2oi_4.pxi.spice
* Created: Wed Sep  2 10:51:23 2020
* 
x_PM_SKY130_FD_SC_LS__A2BB2OI_4%A2_N N_A2_N_c_147_n N_A2_N_M1026_g
+ N_A2_N_c_148_n N_A2_N_M1027_g N_A2_N_c_142_n N_A2_N_c_143_n N_A2_N_c_144_n
+ N_A2_N_M1022_g A2_N A2_N A2_N N_A2_N_c_146_n
+ PM_SKY130_FD_SC_LS__A2BB2OI_4%A2_N
x_PM_SKY130_FD_SC_LS__A2BB2OI_4%A1_N N_A1_N_c_196_n N_A1_N_M1005_g
+ N_A1_N_M1004_g N_A1_N_c_197_n N_A1_N_M1013_g A1_N A1_N N_A1_N_c_195_n
+ PM_SKY130_FD_SC_LS__A2BB2OI_4%A1_N
x_PM_SKY130_FD_SC_LS__A2BB2OI_4%A_114_392# N_A_114_392#_M1022_d
+ N_A_114_392#_M1026_d N_A_114_392#_c_241_n N_A_114_392#_M1002_g
+ N_A_114_392#_c_242_n N_A_114_392#_c_243_n N_A_114_392#_c_244_n
+ N_A_114_392#_M1003_g N_A_114_392#_c_259_n N_A_114_392#_M1000_g
+ N_A_114_392#_c_245_n N_A_114_392#_M1014_g N_A_114_392#_c_260_n
+ N_A_114_392#_M1006_g N_A_114_392#_c_246_n N_A_114_392#_M1023_g
+ N_A_114_392#_c_247_n N_A_114_392#_c_248_n N_A_114_392#_c_262_n
+ N_A_114_392#_M1019_g N_A_114_392#_c_249_n N_A_114_392#_c_263_n
+ N_A_114_392#_M1024_g N_A_114_392#_c_250_n N_A_114_392#_c_251_n
+ N_A_114_392#_c_266_n N_A_114_392#_c_252_n N_A_114_392#_c_253_n
+ N_A_114_392#_c_254_n N_A_114_392#_c_255_n N_A_114_392#_c_256_n
+ N_A_114_392#_c_257_n N_A_114_392#_c_258_n
+ PM_SKY130_FD_SC_LS__A2BB2OI_4%A_114_392#
x_PM_SKY130_FD_SC_LS__A2BB2OI_4%B2 N_B2_c_397_n N_B2_M1001_g N_B2_M1008_g
+ N_B2_c_398_n N_B2_M1016_g N_B2_M1011_g N_B2_c_399_n N_B2_M1018_g N_B2_M1012_g
+ N_B2_c_400_n N_B2_M1021_g N_B2_M1029_g B2 B2 B2 B2 N_B2_c_396_n
+ PM_SKY130_FD_SC_LS__A2BB2OI_4%B2
x_PM_SKY130_FD_SC_LS__A2BB2OI_4%B1 N_B1_M1010_g N_B1_c_482_n N_B1_M1007_g
+ N_B1_M1020_g N_B1_c_483_n N_B1_M1009_g N_B1_M1025_g N_B1_c_484_n N_B1_M1015_g
+ N_B1_M1028_g N_B1_c_485_n N_B1_M1017_g B1 B1 B1 B1 N_B1_c_481_n
+ PM_SKY130_FD_SC_LS__A2BB2OI_4%B1
x_PM_SKY130_FD_SC_LS__A2BB2OI_4%A_29_392# N_A_29_392#_M1026_s
+ N_A_29_392#_M1027_s N_A_29_392#_M1013_s N_A_29_392#_c_558_n
+ N_A_29_392#_c_559_n N_A_29_392#_c_560_n N_A_29_392#_c_561_n
+ N_A_29_392#_c_589_n N_A_29_392#_c_573_n N_A_29_392#_c_562_n
+ N_A_29_392#_c_563_n PM_SKY130_FD_SC_LS__A2BB2OI_4%A_29_392#
x_PM_SKY130_FD_SC_LS__A2BB2OI_4%VPWR N_VPWR_M1005_d N_VPWR_M1001_s
+ N_VPWR_M1018_s N_VPWR_M1007_d N_VPWR_M1015_d N_VPWR_c_607_n N_VPWR_c_608_n
+ N_VPWR_c_609_n N_VPWR_c_610_n N_VPWR_c_611_n N_VPWR_c_612_n N_VPWR_c_613_n
+ N_VPWR_c_614_n N_VPWR_c_615_n N_VPWR_c_616_n VPWR N_VPWR_c_617_n
+ N_VPWR_c_618_n N_VPWR_c_619_n N_VPWR_c_606_n N_VPWR_c_621_n N_VPWR_c_622_n
+ N_VPWR_c_623_n PM_SKY130_FD_SC_LS__A2BB2OI_4%VPWR
x_PM_SKY130_FD_SC_LS__A2BB2OI_4%A_539_368# N_A_539_368#_M1000_s
+ N_A_539_368#_M1006_s N_A_539_368#_M1024_s N_A_539_368#_M1016_d
+ N_A_539_368#_M1021_d N_A_539_368#_M1009_s N_A_539_368#_M1017_s
+ N_A_539_368#_c_712_n N_A_539_368#_c_713_n N_A_539_368#_c_714_n
+ N_A_539_368#_c_730_n N_A_539_368#_c_715_n N_A_539_368#_c_736_n
+ N_A_539_368#_c_737_n N_A_539_368#_c_746_n N_A_539_368#_c_716_n
+ N_A_539_368#_c_754_n N_A_539_368#_c_717_n N_A_539_368#_c_765_n
+ N_A_539_368#_c_718_n N_A_539_368#_c_773_n N_A_539_368#_c_719_n
+ N_A_539_368#_c_720_n N_A_539_368#_c_721_n N_A_539_368#_c_759_n
+ N_A_539_368#_c_722_n N_A_539_368#_c_782_n
+ PM_SKY130_FD_SC_LS__A2BB2OI_4%A_539_368#
x_PM_SKY130_FD_SC_LS__A2BB2OI_4%Y N_Y_M1002_s N_Y_M1014_s N_Y_M1008_d
+ N_Y_M1012_d N_Y_M1000_d N_Y_M1019_d N_Y_c_847_n N_Y_c_835_n N_Y_c_851_n
+ N_Y_c_855_n N_Y_c_836_n N_Y_c_843_n N_Y_c_844_n N_Y_c_837_n N_Y_c_869_n
+ N_Y_c_838_n N_Y_c_839_n N_Y_c_871_n N_Y_c_845_n N_Y_c_840_n Y Y
+ PM_SKY130_FD_SC_LS__A2BB2OI_4%Y
x_PM_SKY130_FD_SC_LS__A2BB2OI_4%VGND N_VGND_M1022_s N_VGND_M1004_d
+ N_VGND_M1003_d N_VGND_M1023_d N_VGND_M1010_d N_VGND_M1025_d N_VGND_c_934_n
+ N_VGND_c_935_n N_VGND_c_936_n N_VGND_c_937_n N_VGND_c_938_n N_VGND_c_939_n
+ N_VGND_c_940_n N_VGND_c_941_n N_VGND_c_942_n N_VGND_c_943_n N_VGND_c_944_n
+ N_VGND_c_945_n N_VGND_c_946_n N_VGND_c_947_n N_VGND_c_948_n N_VGND_c_949_n
+ N_VGND_c_950_n VGND N_VGND_c_951_n N_VGND_c_952_n N_VGND_c_953_n
+ PM_SKY130_FD_SC_LS__A2BB2OI_4%VGND
x_PM_SKY130_FD_SC_LS__A2BB2OI_4%A_914_74# N_A_914_74#_M1008_s
+ N_A_914_74#_M1011_s N_A_914_74#_M1029_s N_A_914_74#_M1020_s
+ N_A_914_74#_M1028_s N_A_914_74#_c_1045_n N_A_914_74#_c_1046_n
+ N_A_914_74#_c_1047_n N_A_914_74#_c_1048_n N_A_914_74#_c_1049_n
+ N_A_914_74#_c_1050_n N_A_914_74#_c_1051_n N_A_914_74#_c_1052_n
+ PM_SKY130_FD_SC_LS__A2BB2OI_4%A_914_74#
cc_1 VNB N_A2_N_c_142_n 0.0251068f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.26
cc_2 VNB N_A2_N_c_143_n 0.0849064f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.26
cc_3 VNB N_A2_N_c_144_n 0.0173058f $X=-0.19 $Y=-0.245 $X2=1.32 $Y2=1.185
cc_4 VNB A2_N 0.00316394f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_5 VNB N_A2_N_c_146_n 0.122325f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.585
cc_6 VNB N_A1_N_M1004_g 0.033515f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.46
cc_7 VNB A1_N 0.00955002f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_8 VNB N_A1_N_c_195_n 0.0282149f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.29
cc_9 VNB N_A_114_392#_c_241_n 0.0169153f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.26
cc_10 VNB N_A_114_392#_c_242_n 0.0218365f $X=-0.19 $Y=-0.245 $X2=1.32 $Y2=0.74
cc_11 VNB N_A_114_392#_c_243_n 0.00949263f $X=-0.19 $Y=-0.245 $X2=1.32 $Y2=0.74
cc_12 VNB N_A_114_392#_c_244_n 0.0157654f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_13 VNB N_A_114_392#_c_245_n 0.0157622f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.29
cc_14 VNB N_A_114_392#_c_246_n 0.0192435f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.605
cc_15 VNB N_A_114_392#_c_247_n 0.0143567f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.535
cc_16 VNB N_A_114_392#_c_248_n 0.0790595f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.535
cc_17 VNB N_A_114_392#_c_249_n 0.0144441f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.925
cc_18 VNB N_A_114_392#_c_250_n 0.0136869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_114_392#_c_251_n 0.0151935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_114_392#_c_252_n 0.00712702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_114_392#_c_253_n 0.0111501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_114_392#_c_254_n 0.00211602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_114_392#_c_255_n 0.0073757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_114_392#_c_256_n 0.00618867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_114_392#_c_257_n 0.00167115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_114_392#_c_258_n 0.0120196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B2_M1008_g 0.0299032f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.46
cc_28 VNB N_B2_M1011_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_29 VNB N_B2_M1012_g 0.0234234f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.585
cc_30 VNB N_B2_M1029_g 0.0240886f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.535
cc_31 VNB B2 0.00365188f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.925
cc_32 VNB N_B2_c_396_n 0.0712771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_B1_M1010_g 0.0230056f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.46
cc_34 VNB N_B1_M1020_g 0.0230578f $X=-0.19 $Y=-0.245 $X2=1.32 $Y2=0.74
cc_35 VNB N_B1_M1025_g 0.0224931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B1_M1028_g 0.0326336f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.605
cc_37 VNB B1 0.0257216f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.925
cc_38 VNB N_B1_c_481_n 0.0747886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VPWR_c_606_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_835_n 0.00206283f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.585
cc_41 VNB N_Y_c_836_n 0.00178621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_837_n 0.00312482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_838_n 0.00135831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_Y_c_839_n 0.00645039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_Y_c_840_n 0.0149701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB Y 0.0116167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB Y 0.00762606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_934_n 0.0176435f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.585
cc_49 VNB N_VGND_c_935_n 0.00451436f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.605
cc_50 VNB N_VGND_c_936_n 0.0026136f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.555
cc_51 VNB N_VGND_c_937_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_938_n 0.0138193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_939_n 0.00481913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_940_n 0.00497771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_941_n 0.0298226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_942_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_943_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_944_n 0.00538852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_945_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_946_n 0.00601765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_947_n 0.0731998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_948_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_949_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_950_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_951_n 0.0266297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_952_n 0.484031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_953_n 0.00613324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_914_74#_c_1045_n 0.0151254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_914_74#_c_1046_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_914_74#_c_1047_n 0.00472705f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.535
cc_71 VNB N_A_914_74#_c_1048_n 0.0037698f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.535
cc_72 VNB N_A_914_74#_c_1049_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_914_74#_c_1050_n 0.0126873f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.925
cc_74 VNB N_A_914_74#_c_1051_n 0.0281813f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.605
cc_75 VNB N_A_914_74#_c_1052_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VPB N_A2_N_c_147_n 0.0185168f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.885
cc_77 VPB N_A2_N_c_148_n 0.0145865f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.885
cc_78 VPB N_A2_N_c_143_n 0.0536943f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.26
cc_79 VPB A2_N 0.00261477f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_80 VPB N_A1_N_c_196_n 0.0153912f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.885
cc_81 VPB N_A1_N_c_197_n 0.0211544f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.26
cc_82 VPB A1_N 0.00757432f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_83 VPB N_A1_N_c_195_n 0.0357514f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.29
cc_84 VPB N_A_114_392#_c_259_n 0.0180164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_114_392#_c_260_n 0.0141056f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.585
cc_86 VPB N_A_114_392#_c_248_n 0.0144253f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.535
cc_87 VPB N_A_114_392#_c_262_n 0.0141056f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.555
cc_88 VPB N_A_114_392#_c_263_n 0.0148127f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.295
cc_89 VPB N_A_114_392#_c_250_n 0.00580711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_114_392#_c_251_n 0.00632584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_114_392#_c_266_n 0.00175613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_B2_c_397_n 0.0152427f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.885
cc_93 VPB N_B2_c_398_n 0.0155127f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.26
cc_94 VPB N_B2_c_399_n 0.0155119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_B2_c_400_n 0.0154187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB B2 0.0112766f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.925
cc_97 VPB N_B2_c_396_n 0.0461514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_B1_c_482_n 0.0154186f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.46
cc_99 VPB N_B1_c_483_n 0.0155119f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_100 VPB N_B1_c_484_n 0.0155127f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=0.585
cc_101 VPB N_B1_c_485_n 0.0208611f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.535
cc_102 VPB B1 0.0222744f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.925
cc_103 VPB N_B1_c_481_n 0.0477908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_29_392#_c_558_n 0.0399513f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_105 VPB N_A_29_392#_c_559_n 0.00478015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_29_392#_c_560_n 0.00987235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_29_392#_c_561_n 0.0025445f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.29
cc_108 VPB N_A_29_392#_c_562_n 0.00288429f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.605
cc_109 VPB N_A_29_392#_c_563_n 0.015297f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.535
cc_110 VPB N_VPWR_c_607_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.29
cc_111 VPB N_VPWR_c_608_n 0.0810243f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.585
cc_112 VPB N_VPWR_c_609_n 0.00770537f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.605
cc_113 VPB N_VPWR_c_610_n 0.00504372f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.535
cc_114 VPB N_VPWR_c_611_n 0.00504372f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.925
cc_115 VPB N_VPWR_c_612_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.605
cc_116 VPB N_VPWR_c_613_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_614_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_615_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_616_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_617_n 0.0371815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_618_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_619_n 0.0245612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_606_n 0.123084f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_621_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_622_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_623_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_539_368#_c_712_n 0.0221874f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.605
cc_128 VPB N_A_539_368#_c_713_n 0.00213603f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.535
cc_129 VPB N_A_539_368#_c_714_n 0.00784407f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.555
cc_130 VPB N_A_539_368#_c_715_n 0.00431993f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.295
cc_131 VPB N_A_539_368#_c_716_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_539_368#_c_717_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_539_368#_c_718_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_539_368#_c_719_n 0.0075508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_539_368#_c_720_n 0.0360166f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_539_368#_c_721_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_539_368#_c_722_n 0.00324197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_Y_c_843_n 0.00749758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_Y_c_844_n 0.00267017f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.295
cc_140 VPB N_Y_c_845_n 0.00118167f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB Y 3.55613e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 N_A2_N_c_148_n N_A1_N_c_196_n 0.00778285f $X=0.945 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A2_N_c_143_n N_A1_N_M1004_g 0.0036141f $X=1.035 $Y=1.26 $X2=0 $Y2=0
cc_144 N_A2_N_c_144_n N_A1_N_M1004_g 0.0176901f $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_145 N_A2_N_c_143_n A1_N 0.00445968f $X=1.035 $Y=1.26 $X2=0 $Y2=0
cc_146 N_A2_N_c_142_n N_A1_N_c_195_n 0.0040525f $X=1.245 $Y=1.26 $X2=0 $Y2=0
cc_147 N_A2_N_c_143_n N_A1_N_c_195_n 0.0153964f $X=1.035 $Y=1.26 $X2=0 $Y2=0
cc_148 N_A2_N_c_147_n N_A_114_392#_c_266_n 0.00456202f $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_149 N_A2_N_c_148_n N_A_114_392#_c_266_n 0.0106243f $X=0.945 $Y=1.885 $X2=0
+ $Y2=0
cc_150 N_A2_N_c_143_n N_A_114_392#_c_266_n 0.0456725f $X=1.035 $Y=1.26 $X2=0
+ $Y2=0
cc_151 A2_N N_A_114_392#_c_266_n 0.0329548f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_152 N_A2_N_c_142_n N_A_114_392#_c_252_n 0.0153082f $X=1.245 $Y=1.26 $X2=0
+ $Y2=0
cc_153 N_A2_N_c_143_n N_A_114_392#_c_252_n 0.0104158f $X=1.035 $Y=1.26 $X2=0
+ $Y2=0
cc_154 N_A2_N_c_144_n N_A_114_392#_c_252_n 0.00832909f $X=1.32 $Y=1.185 $X2=0
+ $Y2=0
cc_155 N_A2_N_c_143_n N_A_114_392#_c_253_n 0.00589853f $X=1.035 $Y=1.26 $X2=0
+ $Y2=0
cc_156 A2_N N_A_114_392#_c_253_n 0.0136491f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_157 N_A2_N_c_146_n N_A_114_392#_c_253_n 0.00181472f $X=0.29 $Y=0.585 $X2=0
+ $Y2=0
cc_158 N_A2_N_c_144_n N_A_114_392#_c_254_n 8.30306e-19 $X=1.32 $Y=1.185 $X2=0
+ $Y2=0
cc_159 N_A2_N_c_147_n N_A_29_392#_c_558_n 0.0118211f $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_160 N_A2_N_c_148_n N_A_29_392#_c_558_n 7.34739e-19 $X=0.945 $Y=1.885 $X2=0
+ $Y2=0
cc_161 N_A2_N_c_143_n N_A_29_392#_c_558_n 0.00265083f $X=1.035 $Y=1.26 $X2=0
+ $Y2=0
cc_162 A2_N N_A_29_392#_c_558_n 0.0273964f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_163 N_A2_N_c_147_n N_A_29_392#_c_559_n 0.0107904f $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_164 N_A2_N_c_148_n N_A_29_392#_c_559_n 0.012504f $X=0.945 $Y=1.885 $X2=0
+ $Y2=0
cc_165 N_A2_N_c_147_n N_A_29_392#_c_560_n 0.00262934f $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_166 N_A2_N_c_148_n N_A_29_392#_c_561_n 9.27995e-19 $X=0.945 $Y=1.885 $X2=0
+ $Y2=0
cc_167 N_A2_N_c_142_n N_A_29_392#_c_561_n 0.00264727f $X=1.245 $Y=1.26 $X2=0
+ $Y2=0
cc_168 N_A2_N_c_142_n N_A_29_392#_c_573_n 0.00102227f $X=1.245 $Y=1.26 $X2=0
+ $Y2=0
cc_169 N_A2_N_c_147_n N_VPWR_c_617_n 0.00278257f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_170 N_A2_N_c_148_n N_VPWR_c_617_n 0.00278271f $X=0.945 $Y=1.885 $X2=0 $Y2=0
cc_171 N_A2_N_c_147_n N_VPWR_c_606_n 0.00357282f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_172 N_A2_N_c_148_n N_VPWR_c_606_n 0.00353907f $X=0.945 $Y=1.885 $X2=0 $Y2=0
cc_173 N_A2_N_c_143_n N_VGND_c_934_n 0.00192879f $X=1.035 $Y=1.26 $X2=0 $Y2=0
cc_174 N_A2_N_c_144_n N_VGND_c_934_n 0.011643f $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_175 A2_N N_VGND_c_934_n 0.0195009f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_176 N_A2_N_c_146_n N_VGND_c_934_n 0.00569436f $X=0.29 $Y=0.585 $X2=0 $Y2=0
cc_177 N_A2_N_c_144_n N_VGND_c_935_n 4.85748e-19 $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_178 A2_N N_VGND_c_941_n 0.0105202f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_179 N_A2_N_c_146_n N_VGND_c_941_n 0.00476771f $X=0.29 $Y=0.585 $X2=0 $Y2=0
cc_180 N_A2_N_c_144_n N_VGND_c_943_n 0.00383152f $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_181 N_A2_N_c_144_n N_VGND_c_952_n 0.00757637f $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_182 A2_N N_VGND_c_952_n 0.0112802f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_183 N_A2_N_c_146_n N_VGND_c_952_n 0.00333647f $X=0.29 $Y=0.585 $X2=0 $Y2=0
cc_184 N_A1_N_M1004_g N_A_114_392#_c_241_n 0.0280367f $X=1.75 $Y=0.74 $X2=0
+ $Y2=0
cc_185 A1_N N_A_114_392#_c_243_n 0.00377293f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_186 A1_N N_A_114_392#_c_259_n 8.03386e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_187 A1_N N_A_114_392#_c_248_n 0.00571268f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_188 N_A1_N_c_195_n N_A_114_392#_c_248_n 9.7315e-19 $X=1.77 $Y=1.635 $X2=0
+ $Y2=0
cc_189 N_A1_N_c_196_n N_A_114_392#_c_266_n 2.66772e-19 $X=1.395 $Y=1.885 $X2=0
+ $Y2=0
cc_190 N_A1_N_c_195_n N_A_114_392#_c_266_n 0.00122825f $X=1.77 $Y=1.635 $X2=0
+ $Y2=0
cc_191 N_A1_N_c_195_n N_A_114_392#_c_252_n 0.00180648f $X=1.77 $Y=1.635 $X2=0
+ $Y2=0
cc_192 N_A1_N_M1004_g N_A_114_392#_c_254_n 8.30306e-19 $X=1.75 $Y=0.74 $X2=0
+ $Y2=0
cc_193 A1_N N_A_114_392#_c_255_n 0.00455708f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_194 A1_N N_A_114_392#_c_257_n 0.00480329f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_195 N_A1_N_c_195_n N_A_114_392#_c_257_n 0.00314031f $X=1.77 $Y=1.635 $X2=0
+ $Y2=0
cc_196 N_A1_N_M1004_g N_A_114_392#_c_258_n 0.0145425f $X=1.75 $Y=0.74 $X2=0
+ $Y2=0
cc_197 A1_N N_A_114_392#_c_258_n 0.04954f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_198 N_A1_N_c_195_n N_A_114_392#_c_258_n 0.00408777f $X=1.77 $Y=1.635 $X2=0
+ $Y2=0
cc_199 N_A1_N_c_196_n N_A_29_392#_c_559_n 0.00125031f $X=1.395 $Y=1.885 $X2=0
+ $Y2=0
cc_200 N_A1_N_c_196_n N_A_29_392#_c_561_n 6.73255e-19 $X=1.395 $Y=1.885 $X2=0
+ $Y2=0
cc_201 N_A1_N_c_196_n N_A_29_392#_c_573_n 0.0140585f $X=1.395 $Y=1.885 $X2=0
+ $Y2=0
cc_202 N_A1_N_c_197_n N_A_29_392#_c_573_n 0.0119563f $X=1.845 $Y=1.885 $X2=0
+ $Y2=0
cc_203 A1_N N_A_29_392#_c_573_n 0.0226735f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_204 N_A1_N_c_195_n N_A_29_392#_c_573_n 0.00597172f $X=1.77 $Y=1.635 $X2=0
+ $Y2=0
cc_205 N_A1_N_c_197_n N_A_29_392#_c_562_n 4.27055e-19 $X=1.845 $Y=1.885 $X2=0
+ $Y2=0
cc_206 A1_N N_A_29_392#_c_562_n 0.0259138f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_207 N_A1_N_c_196_n N_A_29_392#_c_563_n 6.63228e-19 $X=1.395 $Y=1.885 $X2=0
+ $Y2=0
cc_208 N_A1_N_c_197_n N_A_29_392#_c_563_n 0.0104882f $X=1.845 $Y=1.885 $X2=0
+ $Y2=0
cc_209 N_A1_N_c_196_n N_VPWR_c_607_n 0.00975803f $X=1.395 $Y=1.885 $X2=0 $Y2=0
cc_210 N_A1_N_c_197_n N_VPWR_c_607_n 0.0051932f $X=1.845 $Y=1.885 $X2=0 $Y2=0
cc_211 N_A1_N_c_197_n N_VPWR_c_608_n 0.00445602f $X=1.845 $Y=1.885 $X2=0 $Y2=0
cc_212 N_A1_N_c_196_n N_VPWR_c_617_n 0.00413917f $X=1.395 $Y=1.885 $X2=0 $Y2=0
cc_213 N_A1_N_c_196_n N_VPWR_c_606_n 0.0081781f $X=1.395 $Y=1.885 $X2=0 $Y2=0
cc_214 N_A1_N_c_197_n N_VPWR_c_606_n 0.00862391f $X=1.845 $Y=1.885 $X2=0 $Y2=0
cc_215 N_A1_N_M1004_g N_VGND_c_934_n 5.07446e-19 $X=1.75 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A1_N_M1004_g N_VGND_c_935_n 0.0114017f $X=1.75 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A1_N_M1004_g N_VGND_c_943_n 0.00383152f $X=1.75 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A1_N_M1004_g N_VGND_c_952_n 0.00757637f $X=1.75 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A_114_392#_c_263_n N_B2_c_397_n 0.0120464f $X=4.395 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_220 N_A_114_392#_c_263_n B2 0.00100541f $X=4.395 $Y=1.765 $X2=0 $Y2=0
cc_221 N_A_114_392#_c_251_n B2 0.0105313f $X=4.395 $Y=1.475 $X2=0 $Y2=0
cc_222 N_A_114_392#_c_251_n N_B2_c_396_n 0.0173801f $X=4.395 $Y=1.475 $X2=0
+ $Y2=0
cc_223 N_A_114_392#_c_266_n N_A_29_392#_c_558_n 0.0533352f $X=0.72 $Y=2.105
+ $X2=0 $Y2=0
cc_224 N_A_114_392#_M1026_d N_A_29_392#_c_559_n 0.00222494f $X=0.57 $Y=1.96
+ $X2=0 $Y2=0
cc_225 N_A_114_392#_c_266_n N_A_29_392#_c_559_n 0.0144323f $X=0.72 $Y=2.105
+ $X2=0 $Y2=0
cc_226 N_A_114_392#_c_266_n N_A_29_392#_c_561_n 0.0140969f $X=0.72 $Y=2.105
+ $X2=0 $Y2=0
cc_227 N_A_114_392#_c_252_n N_A_29_392#_c_561_n 0.00503831f $X=1.45 $Y=1.215
+ $X2=0 $Y2=0
cc_228 N_A_114_392#_c_266_n N_A_29_392#_c_589_n 0.0379077f $X=0.72 $Y=2.105
+ $X2=0 $Y2=0
cc_229 N_A_114_392#_c_252_n N_A_29_392#_c_573_n 0.00375932f $X=1.45 $Y=1.215
+ $X2=0 $Y2=0
cc_230 N_A_114_392#_c_257_n N_A_29_392#_c_573_n 0.00273982f $X=1.535 $Y=1.215
+ $X2=0 $Y2=0
cc_231 N_A_114_392#_c_259_n N_VPWR_c_608_n 0.00278257f $X=3.045 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_A_114_392#_c_260_n N_VPWR_c_608_n 0.00278257f $X=3.495 $Y=1.765 $X2=0
+ $Y2=0
cc_233 N_A_114_392#_c_262_n N_VPWR_c_608_n 0.00278257f $X=3.945 $Y=1.765 $X2=0
+ $Y2=0
cc_234 N_A_114_392#_c_263_n N_VPWR_c_608_n 0.00278257f $X=4.395 $Y=1.765 $X2=0
+ $Y2=0
cc_235 N_A_114_392#_c_259_n N_VPWR_c_606_n 0.00358623f $X=3.045 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_A_114_392#_c_260_n N_VPWR_c_606_n 0.00353822f $X=3.495 $Y=1.765 $X2=0
+ $Y2=0
cc_237 N_A_114_392#_c_262_n N_VPWR_c_606_n 0.00353822f $X=3.945 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_A_114_392#_c_263_n N_VPWR_c_606_n 0.00353905f $X=4.395 $Y=1.765 $X2=0
+ $Y2=0
cc_239 N_A_114_392#_c_259_n N_A_539_368#_c_712_n 0.0139063f $X=3.045 $Y=1.765
+ $X2=0 $Y2=0
cc_240 N_A_114_392#_c_260_n N_A_539_368#_c_712_n 7.22826e-19 $X=3.495 $Y=1.765
+ $X2=0 $Y2=0
cc_241 N_A_114_392#_c_248_n N_A_539_368#_c_712_n 0.00779138f $X=3.585 $Y=1.475
+ $X2=0 $Y2=0
cc_242 N_A_114_392#_c_255_n N_A_539_368#_c_712_n 0.0198519f $X=2.995 $Y=1.34
+ $X2=0 $Y2=0
cc_243 N_A_114_392#_c_259_n N_A_539_368#_c_713_n 0.0108414f $X=3.045 $Y=1.765
+ $X2=0 $Y2=0
cc_244 N_A_114_392#_c_260_n N_A_539_368#_c_713_n 0.0108414f $X=3.495 $Y=1.765
+ $X2=0 $Y2=0
cc_245 N_A_114_392#_c_259_n N_A_539_368#_c_714_n 0.00262934f $X=3.045 $Y=1.765
+ $X2=0 $Y2=0
cc_246 N_A_114_392#_c_259_n N_A_539_368#_c_730_n 6.41034e-19 $X=3.045 $Y=1.765
+ $X2=0 $Y2=0
cc_247 N_A_114_392#_c_260_n N_A_539_368#_c_730_n 0.0125495f $X=3.495 $Y=1.765
+ $X2=0 $Y2=0
cc_248 N_A_114_392#_c_262_n N_A_539_368#_c_730_n 0.0125495f $X=3.945 $Y=1.765
+ $X2=0 $Y2=0
cc_249 N_A_114_392#_c_263_n N_A_539_368#_c_730_n 6.41034e-19 $X=4.395 $Y=1.765
+ $X2=0 $Y2=0
cc_250 N_A_114_392#_c_262_n N_A_539_368#_c_715_n 0.0108414f $X=3.945 $Y=1.765
+ $X2=0 $Y2=0
cc_251 N_A_114_392#_c_263_n N_A_539_368#_c_715_n 0.0125587f $X=4.395 $Y=1.765
+ $X2=0 $Y2=0
cc_252 N_A_114_392#_c_263_n N_A_539_368#_c_736_n 0.00193585f $X=4.395 $Y=1.765
+ $X2=0 $Y2=0
cc_253 N_A_114_392#_c_262_n N_A_539_368#_c_737_n 6.22492e-19 $X=3.945 $Y=1.765
+ $X2=0 $Y2=0
cc_254 N_A_114_392#_c_263_n N_A_539_368#_c_737_n 0.00919154f $X=4.395 $Y=1.765
+ $X2=0 $Y2=0
cc_255 N_A_114_392#_c_260_n N_A_539_368#_c_721_n 0.00175197f $X=3.495 $Y=1.765
+ $X2=0 $Y2=0
cc_256 N_A_114_392#_c_262_n N_A_539_368#_c_721_n 0.00175197f $X=3.945 $Y=1.765
+ $X2=0 $Y2=0
cc_257 N_A_114_392#_c_241_n N_Y_c_847_n 0.00273433f $X=2.22 $Y=1.22 $X2=0 $Y2=0
cc_258 N_A_114_392#_c_242_n N_Y_c_847_n 6.28576e-19 $X=2.575 $Y=1.295 $X2=0
+ $Y2=0
cc_259 N_A_114_392#_c_258_n N_Y_c_847_n 0.0176844f $X=2.575 $Y=1.34 $X2=0 $Y2=0
cc_260 N_A_114_392#_c_241_n N_Y_c_835_n 0.004978f $X=2.22 $Y=1.22 $X2=0 $Y2=0
cc_261 N_A_114_392#_c_244_n N_Y_c_851_n 0.00947324f $X=2.65 $Y=1.22 $X2=0 $Y2=0
cc_262 N_A_114_392#_c_245_n N_Y_c_851_n 0.00947324f $X=3.08 $Y=1.22 $X2=0 $Y2=0
cc_263 N_A_114_392#_c_248_n N_Y_c_851_n 5.58069e-19 $X=3.585 $Y=1.475 $X2=0
+ $Y2=0
cc_264 N_A_114_392#_c_258_n N_Y_c_851_n 0.0442631f $X=2.575 $Y=1.34 $X2=0 $Y2=0
cc_265 N_A_114_392#_c_259_n N_Y_c_855_n 0.00351644f $X=3.045 $Y=1.765 $X2=0
+ $Y2=0
cc_266 N_A_114_392#_c_260_n N_Y_c_855_n 0.006269f $X=3.495 $Y=1.765 $X2=0 $Y2=0
cc_267 N_A_114_392#_c_260_n N_Y_c_843_n 0.0101246f $X=3.495 $Y=1.765 $X2=0 $Y2=0
cc_268 N_A_114_392#_c_247_n N_Y_c_843_n 0.0030813f $X=3.855 $Y=1.475 $X2=0 $Y2=0
cc_269 N_A_114_392#_c_248_n N_Y_c_843_n 0.00459688f $X=3.585 $Y=1.475 $X2=0
+ $Y2=0
cc_270 N_A_114_392#_c_262_n N_Y_c_843_n 0.00633772f $X=3.945 $Y=1.765 $X2=0
+ $Y2=0
cc_271 N_A_114_392#_c_250_n N_Y_c_843_n 0.00558883f $X=3.945 $Y=1.475 $X2=0
+ $Y2=0
cc_272 N_A_114_392#_c_256_n N_Y_c_843_n 0.0168996f $X=3.42 $Y=1.385 $X2=0 $Y2=0
cc_273 N_A_114_392#_c_259_n N_Y_c_844_n 0.00212373f $X=3.045 $Y=1.765 $X2=0
+ $Y2=0
cc_274 N_A_114_392#_c_248_n N_Y_c_844_n 0.00361007f $X=3.585 $Y=1.475 $X2=0
+ $Y2=0
cc_275 N_A_114_392#_c_256_n N_Y_c_844_n 0.0145791f $X=3.42 $Y=1.385 $X2=0 $Y2=0
cc_276 N_A_114_392#_c_246_n N_Y_c_837_n 0.0115138f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_277 N_A_114_392#_c_247_n N_Y_c_837_n 0.0105398f $X=3.855 $Y=1.475 $X2=0 $Y2=0
cc_278 N_A_114_392#_c_256_n N_Y_c_837_n 0.0132645f $X=3.42 $Y=1.385 $X2=0 $Y2=0
cc_279 N_A_114_392#_c_262_n N_Y_c_869_n 0.006269f $X=3.945 $Y=1.765 $X2=0 $Y2=0
cc_280 N_A_114_392#_c_263_n N_Y_c_869_n 0.00447496f $X=4.395 $Y=1.765 $X2=0
+ $Y2=0
cc_281 N_A_114_392#_c_248_n N_Y_c_871_n 6.18925e-19 $X=3.585 $Y=1.475 $X2=0
+ $Y2=0
cc_282 N_A_114_392#_c_256_n N_Y_c_871_n 0.0147027f $X=3.42 $Y=1.385 $X2=0 $Y2=0
cc_283 N_A_114_392#_c_262_n N_Y_c_845_n 0.00415118f $X=3.945 $Y=1.765 $X2=0
+ $Y2=0
cc_284 N_A_114_392#_c_263_n N_Y_c_845_n 0.00339411f $X=4.395 $Y=1.765 $X2=0
+ $Y2=0
cc_285 N_A_114_392#_c_250_n N_Y_c_845_n 9.41993e-19 $X=3.945 $Y=1.475 $X2=0
+ $Y2=0
cc_286 N_A_114_392#_c_251_n N_Y_c_845_n 3.87046e-19 $X=4.395 $Y=1.475 $X2=0
+ $Y2=0
cc_287 N_A_114_392#_c_249_n N_Y_c_840_n 0.00751003f $X=4.305 $Y=1.475 $X2=0
+ $Y2=0
cc_288 N_A_114_392#_c_251_n N_Y_c_840_n 2.51445e-19 $X=4.395 $Y=1.475 $X2=0
+ $Y2=0
cc_289 N_A_114_392#_c_246_n Y 0.00559274f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_290 N_A_114_392#_c_246_n Y 0.00168909f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_291 N_A_114_392#_c_248_n Y 8.71054e-19 $X=3.585 $Y=1.475 $X2=0 $Y2=0
cc_292 N_A_114_392#_c_249_n Y 0.0124449f $X=4.305 $Y=1.475 $X2=0 $Y2=0
cc_293 N_A_114_392#_c_250_n Y 0.0110051f $X=3.945 $Y=1.475 $X2=0 $Y2=0
cc_294 N_A_114_392#_c_251_n Y 0.00132091f $X=4.395 $Y=1.475 $X2=0 $Y2=0
cc_295 N_A_114_392#_c_256_n Y 0.0183585f $X=3.42 $Y=1.385 $X2=0 $Y2=0
cc_296 N_A_114_392#_c_252_n N_VGND_c_934_n 0.0244338f $X=1.45 $Y=1.215 $X2=0
+ $Y2=0
cc_297 N_A_114_392#_c_254_n N_VGND_c_934_n 0.0225498f $X=1.535 $Y=0.515 $X2=0
+ $Y2=0
cc_298 N_A_114_392#_c_241_n N_VGND_c_935_n 0.00242169f $X=2.22 $Y=1.22 $X2=0
+ $Y2=0
cc_299 N_A_114_392#_c_254_n N_VGND_c_935_n 0.0194859f $X=1.535 $Y=0.515 $X2=0
+ $Y2=0
cc_300 N_A_114_392#_c_258_n N_VGND_c_935_n 0.0161099f $X=2.575 $Y=1.34 $X2=0
+ $Y2=0
cc_301 N_A_114_392#_c_241_n N_VGND_c_936_n 4.26297e-19 $X=2.22 $Y=1.22 $X2=0
+ $Y2=0
cc_302 N_A_114_392#_c_244_n N_VGND_c_936_n 0.00720343f $X=2.65 $Y=1.22 $X2=0
+ $Y2=0
cc_303 N_A_114_392#_c_245_n N_VGND_c_936_n 0.00706632f $X=3.08 $Y=1.22 $X2=0
+ $Y2=0
cc_304 N_A_114_392#_c_246_n N_VGND_c_936_n 4.05984e-19 $X=3.51 $Y=1.22 $X2=0
+ $Y2=0
cc_305 N_A_114_392#_c_245_n N_VGND_c_937_n 0.00383152f $X=3.08 $Y=1.22 $X2=0
+ $Y2=0
cc_306 N_A_114_392#_c_246_n N_VGND_c_937_n 0.00383152f $X=3.51 $Y=1.22 $X2=0
+ $Y2=0
cc_307 N_A_114_392#_c_245_n N_VGND_c_938_n 4.05984e-19 $X=3.08 $Y=1.22 $X2=0
+ $Y2=0
cc_308 N_A_114_392#_c_246_n N_VGND_c_938_n 0.00812981f $X=3.51 $Y=1.22 $X2=0
+ $Y2=0
cc_309 N_A_114_392#_c_254_n N_VGND_c_943_n 0.00749631f $X=1.535 $Y=0.515 $X2=0
+ $Y2=0
cc_310 N_A_114_392#_c_241_n N_VGND_c_945_n 0.00434272f $X=2.22 $Y=1.22 $X2=0
+ $Y2=0
cc_311 N_A_114_392#_c_244_n N_VGND_c_945_n 0.00383152f $X=2.65 $Y=1.22 $X2=0
+ $Y2=0
cc_312 N_A_114_392#_c_241_n N_VGND_c_952_n 0.00820742f $X=2.22 $Y=1.22 $X2=0
+ $Y2=0
cc_313 N_A_114_392#_c_244_n N_VGND_c_952_n 0.00373475f $X=2.65 $Y=1.22 $X2=0
+ $Y2=0
cc_314 N_A_114_392#_c_245_n N_VGND_c_952_n 0.00373475f $X=3.08 $Y=1.22 $X2=0
+ $Y2=0
cc_315 N_A_114_392#_c_246_n N_VGND_c_952_n 0.00373475f $X=3.51 $Y=1.22 $X2=0
+ $Y2=0
cc_316 N_A_114_392#_c_254_n N_VGND_c_952_n 0.0062048f $X=1.535 $Y=0.515 $X2=0
+ $Y2=0
cc_317 N_B2_M1029_g N_B1_M1010_g 0.019323f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_318 N_B2_c_400_n N_B1_c_482_n 0.00946753f $X=6.195 $Y=1.765 $X2=0 $Y2=0
cc_319 B2 B1 0.0124148f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_320 N_B2_c_396_n B1 0.00140487f $X=6.195 $Y=1.557 $X2=0 $Y2=0
cc_321 B2 N_B1_c_481_n 0.00143194f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_322 N_B2_c_396_n N_B1_c_481_n 0.0218264f $X=6.195 $Y=1.557 $X2=0 $Y2=0
cc_323 N_B2_c_397_n N_VPWR_c_608_n 0.0044313f $X=4.845 $Y=1.765 $X2=0 $Y2=0
cc_324 N_B2_c_397_n N_VPWR_c_609_n 0.00331651f $X=4.845 $Y=1.765 $X2=0 $Y2=0
cc_325 N_B2_c_398_n N_VPWR_c_609_n 0.00486623f $X=5.295 $Y=1.765 $X2=0 $Y2=0
cc_326 N_B2_c_399_n N_VPWR_c_610_n 0.00526215f $X=5.745 $Y=1.765 $X2=0 $Y2=0
cc_327 N_B2_c_400_n N_VPWR_c_610_n 0.0106464f $X=6.195 $Y=1.765 $X2=0 $Y2=0
cc_328 N_B2_c_400_n N_VPWR_c_611_n 5.37805e-19 $X=6.195 $Y=1.765 $X2=0 $Y2=0
cc_329 N_B2_c_400_n N_VPWR_c_613_n 0.00413917f $X=6.195 $Y=1.765 $X2=0 $Y2=0
cc_330 N_B2_c_398_n N_VPWR_c_618_n 0.00445602f $X=5.295 $Y=1.765 $X2=0 $Y2=0
cc_331 N_B2_c_399_n N_VPWR_c_618_n 0.00445602f $X=5.745 $Y=1.765 $X2=0 $Y2=0
cc_332 N_B2_c_397_n N_VPWR_c_606_n 0.00853445f $X=4.845 $Y=1.765 $X2=0 $Y2=0
cc_333 N_B2_c_398_n N_VPWR_c_606_n 0.00857589f $X=5.295 $Y=1.765 $X2=0 $Y2=0
cc_334 N_B2_c_399_n N_VPWR_c_606_n 0.00857589f $X=5.745 $Y=1.765 $X2=0 $Y2=0
cc_335 N_B2_c_400_n N_VPWR_c_606_n 0.0081781f $X=6.195 $Y=1.765 $X2=0 $Y2=0
cc_336 N_B2_c_397_n N_A_539_368#_c_715_n 0.0032261f $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_337 N_B2_c_397_n N_A_539_368#_c_736_n 4.27055e-19 $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_338 B2 N_A_539_368#_c_736_n 0.02376f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_339 N_B2_c_397_n N_A_539_368#_c_737_n 0.00919154f $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_340 N_B2_c_398_n N_A_539_368#_c_737_n 6.22492e-19 $X=5.295 $Y=1.765 $X2=0
+ $Y2=0
cc_341 N_B2_c_397_n N_A_539_368#_c_746_n 0.0120074f $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_342 N_B2_c_398_n N_A_539_368#_c_746_n 0.0120074f $X=5.295 $Y=1.765 $X2=0
+ $Y2=0
cc_343 B2 N_A_539_368#_c_746_n 0.0393875f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_344 N_B2_c_396_n N_A_539_368#_c_746_n 0.00130859f $X=6.195 $Y=1.557 $X2=0
+ $Y2=0
cc_345 N_B2_c_397_n N_A_539_368#_c_716_n 6.45594e-19 $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_346 N_B2_c_398_n N_A_539_368#_c_716_n 0.0103431f $X=5.295 $Y=1.765 $X2=0
+ $Y2=0
cc_347 N_B2_c_399_n N_A_539_368#_c_716_n 0.0105452f $X=5.745 $Y=1.765 $X2=0
+ $Y2=0
cc_348 N_B2_c_400_n N_A_539_368#_c_716_n 6.69308e-19 $X=6.195 $Y=1.765 $X2=0
+ $Y2=0
cc_349 N_B2_c_399_n N_A_539_368#_c_754_n 0.0120074f $X=5.745 $Y=1.765 $X2=0
+ $Y2=0
cc_350 N_B2_c_400_n N_A_539_368#_c_754_n 0.0172359f $X=6.195 $Y=1.765 $X2=0
+ $Y2=0
cc_351 B2 N_A_539_368#_c_754_n 0.0293546f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_352 N_B2_c_396_n N_A_539_368#_c_754_n 0.00130859f $X=6.195 $Y=1.557 $X2=0
+ $Y2=0
cc_353 N_B2_c_400_n N_A_539_368#_c_717_n 0.0039133f $X=6.195 $Y=1.765 $X2=0
+ $Y2=0
cc_354 N_B2_c_398_n N_A_539_368#_c_759_n 4.27055e-19 $X=5.295 $Y=1.765 $X2=0
+ $Y2=0
cc_355 N_B2_c_399_n N_A_539_368#_c_759_n 4.27055e-19 $X=5.745 $Y=1.765 $X2=0
+ $Y2=0
cc_356 B2 N_A_539_368#_c_759_n 0.0237598f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_357 N_B2_c_396_n N_A_539_368#_c_759_n 0.00144162f $X=6.195 $Y=1.557 $X2=0
+ $Y2=0
cc_358 N_B2_c_400_n N_A_539_368#_c_722_n 0.00262483f $X=6.195 $Y=1.765 $X2=0
+ $Y2=0
cc_359 N_B2_M1008_g N_Y_c_838_n 0.00262032f $X=4.91 $Y=0.74 $X2=0 $Y2=0
cc_360 N_B2_c_396_n N_Y_c_838_n 0.00221317f $X=6.195 $Y=1.557 $X2=0 $Y2=0
cc_361 N_B2_M1011_g N_Y_c_839_n 0.0140439f $X=5.34 $Y=0.74 $X2=0 $Y2=0
cc_362 N_B2_M1012_g N_Y_c_839_n 0.0140439f $X=5.77 $Y=0.74 $X2=0 $Y2=0
cc_363 N_B2_M1029_g N_Y_c_839_n 0.0054657f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_364 N_B2_c_396_n N_Y_c_839_n 0.00443233f $X=6.195 $Y=1.557 $X2=0 $Y2=0
cc_365 B2 N_Y_c_845_n 0.00479467f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_366 N_B2_M1008_g N_Y_c_840_n 0.0159385f $X=4.91 $Y=0.74 $X2=0 $Y2=0
cc_367 B2 N_Y_c_840_n 0.111129f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_368 N_B2_c_396_n N_Y_c_840_n 0.00202793f $X=6.195 $Y=1.557 $X2=0 $Y2=0
cc_369 N_B2_M1008_g Y 0.005219f $X=4.91 $Y=0.74 $X2=0 $Y2=0
cc_370 B2 Y 0.0277618f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_371 N_B2_c_396_n Y 2.69051e-19 $X=6.195 $Y=1.557 $X2=0 $Y2=0
cc_372 N_B2_M1029_g N_VGND_c_939_n 6.37019e-19 $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_373 N_B2_M1008_g N_VGND_c_947_n 0.00291649f $X=4.91 $Y=0.74 $X2=0 $Y2=0
cc_374 N_B2_M1011_g N_VGND_c_947_n 0.00291649f $X=5.34 $Y=0.74 $X2=0 $Y2=0
cc_375 N_B2_M1012_g N_VGND_c_947_n 0.00291649f $X=5.77 $Y=0.74 $X2=0 $Y2=0
cc_376 N_B2_M1029_g N_VGND_c_947_n 0.00291649f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_377 N_B2_M1008_g N_VGND_c_952_n 0.0036412f $X=4.91 $Y=0.74 $X2=0 $Y2=0
cc_378 N_B2_M1011_g N_VGND_c_952_n 0.00359121f $X=5.34 $Y=0.74 $X2=0 $Y2=0
cc_379 N_B2_M1012_g N_VGND_c_952_n 0.00359121f $X=5.77 $Y=0.74 $X2=0 $Y2=0
cc_380 N_B2_M1029_g N_VGND_c_952_n 0.00359219f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_381 N_B2_M1008_g N_A_914_74#_c_1045_n 0.0104692f $X=4.91 $Y=0.74 $X2=0 $Y2=0
cc_382 N_B2_M1011_g N_A_914_74#_c_1045_n 0.010218f $X=5.34 $Y=0.74 $X2=0 $Y2=0
cc_383 N_B2_M1012_g N_A_914_74#_c_1045_n 0.0101492f $X=5.77 $Y=0.74 $X2=0 $Y2=0
cc_384 N_B2_M1029_g N_A_914_74#_c_1045_n 0.014175f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_385 N_B2_M1029_g N_A_914_74#_c_1048_n 0.0017668f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_386 N_B1_c_482_n N_VPWR_c_610_n 5.37805e-19 $X=6.645 $Y=1.765 $X2=0 $Y2=0
cc_387 N_B1_c_482_n N_VPWR_c_611_n 0.0106464f $X=6.645 $Y=1.765 $X2=0 $Y2=0
cc_388 N_B1_c_483_n N_VPWR_c_611_n 0.00526215f $X=7.095 $Y=1.765 $X2=0 $Y2=0
cc_389 N_B1_c_484_n N_VPWR_c_612_n 0.00486623f $X=7.545 $Y=1.765 $X2=0 $Y2=0
cc_390 N_B1_c_485_n N_VPWR_c_612_n 0.00486623f $X=7.995 $Y=1.765 $X2=0 $Y2=0
cc_391 N_B1_c_482_n N_VPWR_c_613_n 0.00413917f $X=6.645 $Y=1.765 $X2=0 $Y2=0
cc_392 N_B1_c_483_n N_VPWR_c_615_n 0.00445602f $X=7.095 $Y=1.765 $X2=0 $Y2=0
cc_393 N_B1_c_484_n N_VPWR_c_615_n 0.00445602f $X=7.545 $Y=1.765 $X2=0 $Y2=0
cc_394 N_B1_c_485_n N_VPWR_c_619_n 0.00445602f $X=7.995 $Y=1.765 $X2=0 $Y2=0
cc_395 N_B1_c_482_n N_VPWR_c_606_n 0.0081781f $X=6.645 $Y=1.765 $X2=0 $Y2=0
cc_396 N_B1_c_483_n N_VPWR_c_606_n 0.00857589f $X=7.095 $Y=1.765 $X2=0 $Y2=0
cc_397 N_B1_c_484_n N_VPWR_c_606_n 0.00857589f $X=7.545 $Y=1.765 $X2=0 $Y2=0
cc_398 N_B1_c_485_n N_VPWR_c_606_n 0.00861464f $X=7.995 $Y=1.765 $X2=0 $Y2=0
cc_399 N_B1_c_482_n N_A_539_368#_c_717_n 0.0039133f $X=6.645 $Y=1.765 $X2=0
+ $Y2=0
cc_400 N_B1_c_482_n N_A_539_368#_c_765_n 0.0172359f $X=6.645 $Y=1.765 $X2=0
+ $Y2=0
cc_401 N_B1_c_483_n N_A_539_368#_c_765_n 0.0120074f $X=7.095 $Y=1.765 $X2=0
+ $Y2=0
cc_402 B1 N_A_539_368#_c_765_n 0.0289213f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_403 N_B1_c_481_n N_A_539_368#_c_765_n 0.00130859f $X=7.92 $Y=1.515 $X2=0
+ $Y2=0
cc_404 N_B1_c_482_n N_A_539_368#_c_718_n 6.69308e-19 $X=6.645 $Y=1.765 $X2=0
+ $Y2=0
cc_405 N_B1_c_483_n N_A_539_368#_c_718_n 0.0105452f $X=7.095 $Y=1.765 $X2=0
+ $Y2=0
cc_406 N_B1_c_484_n N_A_539_368#_c_718_n 0.0103431f $X=7.545 $Y=1.765 $X2=0
+ $Y2=0
cc_407 N_B1_c_485_n N_A_539_368#_c_718_n 6.45594e-19 $X=7.995 $Y=1.765 $X2=0
+ $Y2=0
cc_408 N_B1_c_484_n N_A_539_368#_c_773_n 0.0120074f $X=7.545 $Y=1.765 $X2=0
+ $Y2=0
cc_409 N_B1_c_485_n N_A_539_368#_c_773_n 0.0120074f $X=7.995 $Y=1.765 $X2=0
+ $Y2=0
cc_410 B1 N_A_539_368#_c_773_n 0.0393875f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_411 N_B1_c_481_n N_A_539_368#_c_773_n 0.00130859f $X=7.92 $Y=1.515 $X2=0
+ $Y2=0
cc_412 N_B1_c_485_n N_A_539_368#_c_719_n 4.27055e-19 $X=7.995 $Y=1.765 $X2=0
+ $Y2=0
cc_413 B1 N_A_539_368#_c_719_n 0.0265364f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_414 N_B1_c_484_n N_A_539_368#_c_720_n 6.45594e-19 $X=7.545 $Y=1.765 $X2=0
+ $Y2=0
cc_415 N_B1_c_485_n N_A_539_368#_c_720_n 0.0104891f $X=7.995 $Y=1.765 $X2=0
+ $Y2=0
cc_416 N_B1_c_482_n N_A_539_368#_c_722_n 0.00262483f $X=6.645 $Y=1.765 $X2=0
+ $Y2=0
cc_417 N_B1_c_483_n N_A_539_368#_c_782_n 4.27055e-19 $X=7.095 $Y=1.765 $X2=0
+ $Y2=0
cc_418 N_B1_c_484_n N_A_539_368#_c_782_n 4.27055e-19 $X=7.545 $Y=1.765 $X2=0
+ $Y2=0
cc_419 B1 N_A_539_368#_c_782_n 0.0237598f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_420 N_B1_c_481_n N_A_539_368#_c_782_n 0.00144162f $X=7.92 $Y=1.515 $X2=0
+ $Y2=0
cc_421 N_B1_M1010_g N_VGND_c_939_n 0.0100344f $X=6.63 $Y=0.74 $X2=0 $Y2=0
cc_422 N_B1_M1020_g N_VGND_c_939_n 0.00204878f $X=7.06 $Y=0.74 $X2=0 $Y2=0
cc_423 N_B1_M1020_g N_VGND_c_940_n 5.20618e-19 $X=7.06 $Y=0.74 $X2=0 $Y2=0
cc_424 N_B1_M1025_g N_VGND_c_940_n 0.0101191f $X=7.49 $Y=0.74 $X2=0 $Y2=0
cc_425 N_B1_M1028_g N_VGND_c_940_n 0.00341128f $X=7.92 $Y=0.74 $X2=0 $Y2=0
cc_426 N_B1_M1010_g N_VGND_c_947_n 0.00383152f $X=6.63 $Y=0.74 $X2=0 $Y2=0
cc_427 N_B1_M1020_g N_VGND_c_949_n 0.00434272f $X=7.06 $Y=0.74 $X2=0 $Y2=0
cc_428 N_B1_M1025_g N_VGND_c_949_n 0.00383152f $X=7.49 $Y=0.74 $X2=0 $Y2=0
cc_429 N_B1_M1028_g N_VGND_c_951_n 0.00434272f $X=7.92 $Y=0.74 $X2=0 $Y2=0
cc_430 N_B1_M1010_g N_VGND_c_952_n 0.00757637f $X=6.63 $Y=0.74 $X2=0 $Y2=0
cc_431 N_B1_M1020_g N_VGND_c_952_n 0.00820284f $X=7.06 $Y=0.74 $X2=0 $Y2=0
cc_432 N_B1_M1025_g N_VGND_c_952_n 0.0075754f $X=7.49 $Y=0.74 $X2=0 $Y2=0
cc_433 N_B1_M1028_g N_VGND_c_952_n 0.00824501f $X=7.92 $Y=0.74 $X2=0 $Y2=0
cc_434 N_B1_M1010_g N_A_914_74#_c_1047_n 0.0174499f $X=6.63 $Y=0.74 $X2=0 $Y2=0
cc_435 N_B1_M1020_g N_A_914_74#_c_1047_n 0.0111034f $X=7.06 $Y=0.74 $X2=0 $Y2=0
cc_436 B1 N_A_914_74#_c_1047_n 0.0282658f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_437 N_B1_c_481_n N_A_914_74#_c_1047_n 0.00224206f $X=7.92 $Y=1.515 $X2=0
+ $Y2=0
cc_438 N_B1_M1010_g N_A_914_74#_c_1049_n 6.58468e-19 $X=6.63 $Y=0.74 $X2=0 $Y2=0
cc_439 N_B1_M1020_g N_A_914_74#_c_1049_n 0.00918302f $X=7.06 $Y=0.74 $X2=0 $Y2=0
cc_440 N_B1_M1025_g N_A_914_74#_c_1049_n 3.97481e-19 $X=7.49 $Y=0.74 $X2=0 $Y2=0
cc_441 N_B1_M1025_g N_A_914_74#_c_1050_n 0.0130918f $X=7.49 $Y=0.74 $X2=0 $Y2=0
cc_442 N_B1_M1028_g N_A_914_74#_c_1050_n 0.0132972f $X=7.92 $Y=0.74 $X2=0 $Y2=0
cc_443 B1 N_A_914_74#_c_1050_n 0.0748451f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_444 N_B1_c_481_n N_A_914_74#_c_1050_n 0.00465078f $X=7.92 $Y=1.515 $X2=0
+ $Y2=0
cc_445 N_B1_M1025_g N_A_914_74#_c_1051_n 6.56397e-19 $X=7.49 $Y=0.74 $X2=0 $Y2=0
cc_446 N_B1_M1028_g N_A_914_74#_c_1051_n 0.0100626f $X=7.92 $Y=0.74 $X2=0 $Y2=0
cc_447 N_B1_M1020_g N_A_914_74#_c_1052_n 0.00157732f $X=7.06 $Y=0.74 $X2=0 $Y2=0
cc_448 B1 N_A_914_74#_c_1052_n 0.0213626f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_449 N_B1_c_481_n N_A_914_74#_c_1052_n 0.00232957f $X=7.92 $Y=1.515 $X2=0
+ $Y2=0
cc_450 N_A_29_392#_c_573_n N_VPWR_M1005_d 0.00402456f $X=1.905 $Y=2.055
+ $X2=-0.19 $Y2=1.66
cc_451 N_A_29_392#_c_559_n N_VPWR_c_607_n 0.0123543f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_452 N_A_29_392#_c_589_n N_VPWR_c_607_n 0.0379077f $X=1.17 $Y=2.815 $X2=0
+ $Y2=0
cc_453 N_A_29_392#_c_573_n N_VPWR_c_607_n 0.0154248f $X=1.905 $Y=2.055 $X2=0
+ $Y2=0
cc_454 N_A_29_392#_c_563_n N_VPWR_c_607_n 0.0449538f $X=2.07 $Y=2.815 $X2=0
+ $Y2=0
cc_455 N_A_29_392#_c_563_n N_VPWR_c_608_n 0.0145938f $X=2.07 $Y=2.815 $X2=0
+ $Y2=0
cc_456 N_A_29_392#_c_559_n N_VPWR_c_617_n 0.0531736f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_457 N_A_29_392#_c_560_n N_VPWR_c_617_n 0.0236039f $X=0.435 $Y=2.99 $X2=0
+ $Y2=0
cc_458 N_A_29_392#_c_559_n N_VPWR_c_606_n 0.0297434f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_459 N_A_29_392#_c_560_n N_VPWR_c_606_n 0.012761f $X=0.435 $Y=2.99 $X2=0 $Y2=0
cc_460 N_A_29_392#_c_563_n N_VPWR_c_606_n 0.0120466f $X=2.07 $Y=2.815 $X2=0
+ $Y2=0
cc_461 N_A_29_392#_c_562_n N_A_539_368#_c_712_n 0.00803119f $X=2.07 $Y=2.14
+ $X2=0 $Y2=0
cc_462 N_A_29_392#_c_563_n N_A_539_368#_c_712_n 0.0340606f $X=2.07 $Y=2.815
+ $X2=0 $Y2=0
cc_463 N_A_29_392#_c_563_n N_A_539_368#_c_714_n 0.00354317f $X=2.07 $Y=2.815
+ $X2=0 $Y2=0
cc_464 N_VPWR_c_608_n N_A_539_368#_c_713_n 0.03588f $X=4.985 $Y=3.33 $X2=0 $Y2=0
cc_465 N_VPWR_c_606_n N_A_539_368#_c_713_n 0.0201952f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_466 N_VPWR_c_608_n N_A_539_368#_c_714_n 0.0236039f $X=4.985 $Y=3.33 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_606_n N_A_539_368#_c_714_n 0.012761f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_468 N_VPWR_c_608_n N_A_539_368#_c_715_n 0.0594312f $X=4.985 $Y=3.33 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_609_n N_A_539_368#_c_715_n 0.0119328f $X=5.07 $Y=2.455 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_606_n N_A_539_368#_c_715_n 0.0328875f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_471 N_VPWR_c_609_n N_A_539_368#_c_737_n 0.0400262f $X=5.07 $Y=2.455 $X2=0
+ $Y2=0
cc_472 N_VPWR_M1001_s N_A_539_368#_c_746_n 0.00408911f $X=4.92 $Y=1.84 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_609_n N_A_539_368#_c_746_n 0.0136682f $X=5.07 $Y=2.455 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_609_n N_A_539_368#_c_716_n 0.0449718f $X=5.07 $Y=2.455 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_610_n N_A_539_368#_c_716_n 0.0462948f $X=5.97 $Y=2.455 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_618_n N_A_539_368#_c_716_n 0.014552f $X=5.885 $Y=3.33 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_606_n N_A_539_368#_c_716_n 0.0119791f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_478 N_VPWR_M1018_s N_A_539_368#_c_754_n 0.00384138f $X=5.82 $Y=1.84 $X2=0
+ $Y2=0
cc_479 N_VPWR_c_610_n N_A_539_368#_c_754_n 0.0154248f $X=5.97 $Y=2.455 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_610_n N_A_539_368#_c_717_n 0.0440249f $X=5.97 $Y=2.455 $X2=0
+ $Y2=0
cc_481 N_VPWR_c_611_n N_A_539_368#_c_717_n 0.0440249f $X=6.87 $Y=2.455 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_613_n N_A_539_368#_c_717_n 0.00749631f $X=6.705 $Y=3.33 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_606_n N_A_539_368#_c_717_n 0.0062048f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_484 N_VPWR_M1007_d N_A_539_368#_c_765_n 0.00384138f $X=6.72 $Y=1.84 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_611_n N_A_539_368#_c_765_n 0.0154248f $X=6.87 $Y=2.455 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_611_n N_A_539_368#_c_718_n 0.0462948f $X=6.87 $Y=2.455 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_612_n N_A_539_368#_c_718_n 0.0449718f $X=7.77 $Y=2.455 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_615_n N_A_539_368#_c_718_n 0.014552f $X=7.685 $Y=3.33 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_606_n N_A_539_368#_c_718_n 0.0119791f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_490 N_VPWR_M1015_d N_A_539_368#_c_773_n 0.00408911f $X=7.62 $Y=1.84 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_612_n N_A_539_368#_c_773_n 0.0136682f $X=7.77 $Y=2.455 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_612_n N_A_539_368#_c_720_n 0.0449718f $X=7.77 $Y=2.455 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_619_n N_A_539_368#_c_720_n 0.0145938f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_494 N_VPWR_c_606_n N_A_539_368#_c_720_n 0.0120466f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_495 N_VPWR_c_608_n N_A_539_368#_c_721_n 0.0235512f $X=4.985 $Y=3.33 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_606_n N_A_539_368#_c_721_n 0.0126924f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_497 N_A_539_368#_c_713_n N_Y_M1000_d 0.00243452f $X=3.555 $Y=2.99 $X2=0 $Y2=0
cc_498 N_A_539_368#_c_715_n N_Y_M1019_d 0.00243452f $X=4.455 $Y=2.99 $X2=0 $Y2=0
cc_499 N_A_539_368#_c_712_n N_Y_c_855_n 0.0550085f $X=2.82 $Y=1.985 $X2=0 $Y2=0
cc_500 N_A_539_368#_c_713_n N_Y_c_855_n 0.012787f $X=3.555 $Y=2.99 $X2=0 $Y2=0
cc_501 N_A_539_368#_c_730_n N_Y_c_855_n 0.0439674f $X=3.72 $Y=2.225 $X2=0 $Y2=0
cc_502 N_A_539_368#_M1006_s N_Y_c_843_n 0.00197722f $X=3.57 $Y=1.84 $X2=0 $Y2=0
cc_503 N_A_539_368#_c_730_n N_Y_c_843_n 0.0171813f $X=3.72 $Y=2.225 $X2=0 $Y2=0
cc_504 N_A_539_368#_c_712_n N_Y_c_844_n 0.00513432f $X=2.82 $Y=1.985 $X2=0 $Y2=0
cc_505 N_A_539_368#_c_730_n N_Y_c_869_n 0.0439674f $X=3.72 $Y=2.225 $X2=0 $Y2=0
cc_506 N_A_539_368#_c_715_n N_Y_c_869_n 0.012787f $X=4.455 $Y=2.99 $X2=0 $Y2=0
cc_507 N_A_539_368#_c_736_n N_Y_c_869_n 0.0117758f $X=4.62 $Y=2.12 $X2=0 $Y2=0
cc_508 N_A_539_368#_c_737_n N_Y_c_869_n 0.0400262f $X=4.62 $Y=2.815 $X2=0 $Y2=0
cc_509 N_A_539_368#_c_722_n N_A_914_74#_c_1048_n 0.00609927f $X=6.42 $Y=1.985
+ $X2=0 $Y2=0
cc_510 N_Y_c_851_n N_VGND_M1003_d 0.00330219f $X=3.21 $Y=0.875 $X2=0 $Y2=0
cc_511 N_Y_c_837_n N_VGND_M1023_d 0.00668617f $X=3.965 $Y=0.875 $X2=0 $Y2=0
cc_512 N_Y_c_835_n N_VGND_c_935_n 0.0158235f $X=2.435 $Y=0.515 $X2=0 $Y2=0
cc_513 N_Y_c_835_n N_VGND_c_936_n 0.0104051f $X=2.435 $Y=0.515 $X2=0 $Y2=0
cc_514 N_Y_c_851_n N_VGND_c_936_n 0.0166744f $X=3.21 $Y=0.875 $X2=0 $Y2=0
cc_515 N_Y_c_836_n N_VGND_c_936_n 0.0103637f $X=3.295 $Y=0.515 $X2=0 $Y2=0
cc_516 N_Y_c_836_n N_VGND_c_937_n 0.00743725f $X=3.295 $Y=0.515 $X2=0 $Y2=0
cc_517 N_Y_c_836_n N_VGND_c_938_n 0.0103637f $X=3.295 $Y=0.515 $X2=0 $Y2=0
cc_518 N_Y_c_837_n N_VGND_c_938_n 0.0214241f $X=3.965 $Y=0.875 $X2=0 $Y2=0
cc_519 N_Y_c_835_n N_VGND_c_945_n 0.0109081f $X=2.435 $Y=0.515 $X2=0 $Y2=0
cc_520 N_Y_c_835_n N_VGND_c_952_n 0.00901008f $X=2.435 $Y=0.515 $X2=0 $Y2=0
cc_521 N_Y_c_851_n N_VGND_c_952_n 0.0122738f $X=3.21 $Y=0.875 $X2=0 $Y2=0
cc_522 N_Y_c_836_n N_VGND_c_952_n 0.00618197f $X=3.295 $Y=0.515 $X2=0 $Y2=0
cc_523 N_Y_c_837_n N_VGND_c_952_n 0.00943228f $X=3.965 $Y=0.875 $X2=0 $Y2=0
cc_524 N_Y_c_840_n N_VGND_c_952_n 0.0113458f $X=4.96 $Y=0.95 $X2=0 $Y2=0
cc_525 Y N_VGND_c_952_n 0.0119508f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_526 N_Y_c_840_n N_A_914_74#_M1008_s 0.00382948f $X=4.96 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_527 N_Y_c_839_n N_A_914_74#_M1011_s 0.00177442f $X=5.985 $Y=0.95 $X2=0 $Y2=0
cc_528 N_Y_M1008_d N_A_914_74#_c_1045_n 0.00179007f $X=4.985 $Y=0.37 $X2=0 $Y2=0
cc_529 N_Y_M1012_d N_A_914_74#_c_1045_n 0.00179007f $X=5.845 $Y=0.37 $X2=0 $Y2=0
cc_530 N_Y_c_838_n N_A_914_74#_c_1045_n 0.0628697f $X=5.14 $Y=0.95 $X2=0 $Y2=0
cc_531 N_Y_c_840_n N_A_914_74#_c_1045_n 0.0253733f $X=4.96 $Y=0.95 $X2=0 $Y2=0
cc_532 N_Y_c_839_n N_A_914_74#_c_1048_n 0.00561736f $X=5.985 $Y=0.95 $X2=0 $Y2=0
cc_533 N_VGND_c_938_n N_A_914_74#_c_1045_n 0.00868144f $X=3.725 $Y=0.525 $X2=0
+ $Y2=0
cc_534 N_VGND_c_947_n N_A_914_74#_c_1045_n 0.0729484f $X=6.68 $Y=0 $X2=0 $Y2=0
cc_535 N_VGND_c_952_n N_A_914_74#_c_1045_n 0.0614753f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_536 N_VGND_c_939_n N_A_914_74#_c_1046_n 0.00947603f $X=6.845 $Y=0.675 $X2=0
+ $Y2=0
cc_537 N_VGND_c_947_n N_A_914_74#_c_1046_n 0.00758556f $X=6.68 $Y=0 $X2=0 $Y2=0
cc_538 N_VGND_c_952_n N_A_914_74#_c_1046_n 0.00627867f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_539 N_VGND_M1010_d N_A_914_74#_c_1047_n 0.00176461f $X=6.705 $Y=0.37 $X2=0
+ $Y2=0
cc_540 N_VGND_c_939_n N_A_914_74#_c_1047_n 0.0152916f $X=6.845 $Y=0.675 $X2=0
+ $Y2=0
cc_541 N_VGND_c_939_n N_A_914_74#_c_1049_n 0.0175587f $X=6.845 $Y=0.675 $X2=0
+ $Y2=0
cc_542 N_VGND_c_940_n N_A_914_74#_c_1049_n 0.0175587f $X=7.705 $Y=0.675 $X2=0
+ $Y2=0
cc_543 N_VGND_c_949_n N_A_914_74#_c_1049_n 0.0109942f $X=7.54 $Y=0 $X2=0 $Y2=0
cc_544 N_VGND_c_952_n N_A_914_74#_c_1049_n 0.00904371f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_545 N_VGND_M1025_d N_A_914_74#_c_1050_n 0.00176461f $X=7.565 $Y=0.37 $X2=0
+ $Y2=0
cc_546 N_VGND_c_940_n N_A_914_74#_c_1050_n 0.0152916f $X=7.705 $Y=0.675 $X2=0
+ $Y2=0
cc_547 N_VGND_c_940_n N_A_914_74#_c_1051_n 0.0182902f $X=7.705 $Y=0.675 $X2=0
+ $Y2=0
cc_548 N_VGND_c_951_n N_A_914_74#_c_1051_n 0.0145639f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_549 N_VGND_c_952_n N_A_914_74#_c_1051_n 0.0119984f $X=8.4 $Y=0 $X2=0 $Y2=0
