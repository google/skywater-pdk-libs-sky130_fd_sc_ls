* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
M1000 Q a_2580_74# VGND VNB nshort w=740000u l=150000u
+  ad=5.291e+11p pd=4.39e+06u as=2.27325e+12p ps=1.996e+07u
M1001 VPWR SCD a_414_464# VPB phighvt w=640000u l=150000u
+  ad=3.1281e+12p pd=2.706e+07u as=1.728e+11p ps=1.82e+06u
M1002 a_1017_81# a_616_74# a_288_464# VNB nshort w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=3.592e+11p ps=3.44e+06u
M1003 VGND SET_B a_1445_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1004 VPWR a_1201_55# a_1140_495# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.8235e+11p ps=1.93e+06u
M1005 a_1823_524# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=6.171e+11p pd=6.09e+06u as=0p ps=0u
M1006 VPWR SET_B a_1201_55# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1007 a_2227_74# a_2191_180# a_2149_74# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=1.008e+11p ps=1.32e+06u
M1008 VGND a_1823_524# a_2580_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1009 a_2103_508# a_803_74# a_1823_524# VPB phighvt w=420000u l=150000u
+  ad=1.995e+11p pd=1.79e+06u as=0p ps=0u
M1010 a_1823_524# a_803_74# a_1677_74# VNB nshort w=640000u l=150000u
+  ad=3.963e+11p pd=3.85e+06u as=3.584e+11p ps=3.68e+06u
M1011 Q a_2580_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1012 a_414_464# a_27_74# a_288_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=4.311e+11p ps=3.67e+06u
M1013 VPWR a_1823_524# a_2191_180# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.239e+11p ps=1.43e+06u
M1014 VGND a_1017_81# a_1677_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Q a_2580_74# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1620_373# a_616_74# a_1823_524# VPB phighvt w=840000u l=150000u
+  ad=5.04e+11p pd=4.56e+06u as=0p ps=0u
M1017 a_417_74# SCE a_288_464# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1018 VGND SCD a_417_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_1201_55# a_1153_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1020 a_1153_81# a_803_74# a_1017_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_803_74# a_616_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1022 a_2580_74# a_1823_524# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1023 VGND a_2580_74# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1445_74# a_1017_81# a_1201_55# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1025 VGND CLK a_616_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1026 a_2149_74# a_616_74# a_1823_524# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_2580_74# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR CLK a_616_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1029 a_1017_81# a_803_74# a_288_464# VPB phighvt w=420000u l=150000u
+  ad=1.9495e+11p pd=1.99e+06u as=0p ps=0u
M1030 a_1823_524# a_616_74# a_1620_373# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1201_55# a_1017_81# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1140_495# a_616_74# a_1017_81# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_1823_524# a_2580_74# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_288_464# D a_204_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1035 a_1620_373# a_1017_81# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1677_74# a_803_74# a_1823_524# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Q a_2580_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND SET_B a_2227_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_2191_180# a_1823_524# VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1040 a_803_74# a_616_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.256e+11p pd=2.93e+06u as=0p ps=0u
M1041 a_222_74# a_27_74# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1042 a_288_464# D a_222_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VPWR SCE a_27_74# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1044 a_204_464# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VGND SCE a_27_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1046 VPWR a_2191_180# a_2103_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VPWR a_1017_81# a_1620_373# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_1677_74# a_1017_81# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VPWR a_2580_74# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 VPWR a_2580_74# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
