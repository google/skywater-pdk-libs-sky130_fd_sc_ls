* File: sky130_fd_sc_ls__o31ai_2.pxi.spice
* Created: Fri Aug 28 13:53:37 2020
* 
x_PM_SKY130_FD_SC_LS__O31AI_2%A1 N_A1_M1012_g N_A1_c_85_n N_A1_M1005_g
+ N_A1_c_86_n N_A1_M1006_g N_A1_c_82_n N_A1_M1014_g A1 A1 A1 N_A1_c_84_n
+ PM_SKY130_FD_SC_LS__O31AI_2%A1
x_PM_SKY130_FD_SC_LS__O31AI_2%A2 N_A2_c_134_n N_A2_M1010_g N_A2_M1004_g
+ N_A2_c_135_n N_A2_M1015_g N_A2_M1011_g A2 A2 N_A2_c_133_n
+ PM_SKY130_FD_SC_LS__O31AI_2%A2
x_PM_SKY130_FD_SC_LS__O31AI_2%A3 N_A3_M1001_g N_A3_c_186_n N_A3_c_187_n
+ N_A3_c_191_n N_A3_M1009_g N_A3_c_192_n N_A3_M1013_g N_A3_M1002_g A3
+ N_A3_c_189_n N_A3_c_190_n PM_SKY130_FD_SC_LS__O31AI_2%A3
x_PM_SKY130_FD_SC_LS__O31AI_2%B1 N_B1_M1007_g N_B1_c_256_n N_B1_M1000_g
+ N_B1_M1008_g N_B1_c_257_n N_B1_M1003_g N_B1_c_253_n B1 N_B1_c_255_n
+ PM_SKY130_FD_SC_LS__O31AI_2%B1
x_PM_SKY130_FD_SC_LS__O31AI_2%A_28_368# N_A_28_368#_M1005_s N_A_28_368#_M1006_s
+ N_A_28_368#_M1015_s N_A_28_368#_c_307_n N_A_28_368#_c_308_n
+ N_A_28_368#_c_313_n N_A_28_368#_c_309_n N_A_28_368#_c_323_n
+ N_A_28_368#_c_319_n N_A_28_368#_c_310_n PM_SKY130_FD_SC_LS__O31AI_2%A_28_368#
x_PM_SKY130_FD_SC_LS__O31AI_2%VPWR N_VPWR_M1005_d N_VPWR_M1000_d N_VPWR_c_350_n
+ N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_353_n VPWR N_VPWR_c_354_n
+ N_VPWR_c_355_n N_VPWR_c_349_n N_VPWR_c_357_n PM_SKY130_FD_SC_LS__O31AI_2%VPWR
x_PM_SKY130_FD_SC_LS__O31AI_2%A_297_368# N_A_297_368#_M1010_d
+ N_A_297_368#_M1009_d N_A_297_368#_c_408_n N_A_297_368#_c_398_n
+ N_A_297_368#_c_399_n N_A_297_368#_c_404_n
+ PM_SKY130_FD_SC_LS__O31AI_2%A_297_368#
x_PM_SKY130_FD_SC_LS__O31AI_2%Y N_Y_M1007_d N_Y_M1009_s N_Y_M1013_s N_Y_M1003_s
+ N_Y_c_427_n N_Y_c_424_n N_Y_c_425_n N_Y_c_440_n N_Y_c_460_n N_Y_c_444_n
+ N_Y_c_428_n N_Y_c_429_n N_Y_c_430_n N_Y_c_426_n N_Y_c_454_n Y Y
+ PM_SKY130_FD_SC_LS__O31AI_2%Y
x_PM_SKY130_FD_SC_LS__O31AI_2%A_27_74# N_A_27_74#_M1012_s N_A_27_74#_M1014_s
+ N_A_27_74#_M1011_s N_A_27_74#_M1002_s N_A_27_74#_M1008_s N_A_27_74#_c_502_n
+ N_A_27_74#_c_503_n N_A_27_74#_c_504_n N_A_27_74#_c_505_n N_A_27_74#_c_506_n
+ N_A_27_74#_c_530_n N_A_27_74#_c_537_n N_A_27_74#_c_541_n N_A_27_74#_c_507_n
+ N_A_27_74#_c_508_n N_A_27_74#_c_509_n N_A_27_74#_c_510_n N_A_27_74#_c_511_n
+ PM_SKY130_FD_SC_LS__O31AI_2%A_27_74#
x_PM_SKY130_FD_SC_LS__O31AI_2%VGND N_VGND_M1012_d N_VGND_M1004_d N_VGND_M1001_d
+ N_VGND_c_583_n N_VGND_c_584_n N_VGND_c_585_n VGND N_VGND_c_586_n
+ N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n N_VGND_c_590_n N_VGND_c_591_n
+ N_VGND_c_592_n PM_SKY130_FD_SC_LS__O31AI_2%VGND
cc_1 VNB N_A1_M1012_g 0.0339584f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_c_82_n 0.0157773f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.185
cc_3 VNB A1 0.0218337f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_4 VNB N_A1_c_84_n 0.0574047f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.475
cc_5 VNB N_A2_M1004_g 0.0254433f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_6 VNB N_A2_M1011_g 0.0253921f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.74
cc_7 VNB A2 0.00408815f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_8 VNB N_A2_c_133_n 0.0491661f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_9 VNB N_A3_M1001_g 0.0254342f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_10 VNB N_A3_c_186_n 0.0144872f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.765
cc_11 VNB N_A3_c_187_n 0.0119391f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_12 VNB N_A3_M1002_g 0.0262448f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_13 VNB N_A3_c_189_n 0.00217772f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.475
cc_14 VNB N_A3_c_190_n 0.0392491f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_15 VNB N_B1_M1007_g 0.0205226f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_16 VNB N_B1_M1008_g 0.0255449f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_17 VNB N_B1_c_253_n 0.00219487f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_18 VNB B1 0.0102709f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.475
cc_19 VNB N_B1_c_255_n 0.08416f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.185
cc_20 VNB N_VPWR_c_349_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_424_n 0.0147535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_425_n 8.30186e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.475
cc_23 VNB N_Y_c_426_n 0.00570061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_502_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_503_n 0.00263637f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.475
cc_26 VNB N_A_27_74#_c_504_n 0.0104987f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.475
cc_27 VNB N_A_27_74#_c_505_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_28 VNB N_A_27_74#_c_506_n 0.010404f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.185
cc_29 VNB N_A_27_74#_c_507_n 0.0126811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_74#_c_508_n 0.00163372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_74#_c_509_n 0.0222992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_74#_c_510_n 0.00322614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_74#_c_511_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_583_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.74
cc_35 VNB N_VGND_c_584_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_36 VNB N_VGND_c_585_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_586_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_38 VNB N_VGND_c_587_n 0.0387921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_588_n 0.271117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_589_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_590_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_591_n 0.0182584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_592_n 0.0206062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_A1_c_85_n 0.0201401f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_45 VPB N_A1_c_86_n 0.0157885f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_46 VPB A1 0.0147904f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_47 VPB N_A1_c_84_n 0.0205655f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.475
cc_48 VPB N_A2_c_134_n 0.015911f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_49 VPB N_A2_c_135_n 0.0183174f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_50 VPB A2 0.00804723f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_51 VPB N_A2_c_133_n 0.0212651f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_52 VPB N_A3_c_191_n 0.017528f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_53 VPB N_A3_c_192_n 0.0158201f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_54 VPB N_A3_c_189_n 0.00461917f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.475
cc_55 VPB N_A3_c_190_n 0.0212204f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_56 VPB N_B1_c_256_n 0.016278f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_57 VPB N_B1_c_257_n 0.0211552f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.74
cc_58 VPB B1 0.00389529f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.475
cc_59 VPB N_B1_c_255_n 0.0243266f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.185
cc_60 VPB N_A_28_368#_c_307_n 0.00739392f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_61 VPB N_A_28_368#_c_308_n 0.0339313f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.74
cc_62 VPB N_A_28_368#_c_309_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_28_368#_c_310_n 0.00763828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_350_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_65 VPB N_VPWR_c_351_n 0.00799266f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.74
cc_66 VPB N_VPWR_c_352_n 0.0788082f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_67 VPB N_VPWR_c_353_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_354_n 0.0181665f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.475
cc_69 VPB N_VPWR_c_355_n 0.0201062f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_70 VPB N_VPWR_c_349_n 0.080252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_357_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_297_368#_c_398_n 0.020921f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.185
cc_73 VPB N_A_297_368#_c_399_n 0.00262155f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.74
cc_74 VPB N_Y_c_427_n 0.00583784f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_75 VPB N_Y_c_428_n 0.007175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_Y_c_429_n 0.0391931f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_77 VPB N_Y_c_430_n 0.0057129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_Y_c_426_n 0.00290204f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB Y 0.00289633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 N_A1_c_86_n N_A2_c_134_n 0.0123855f $X=0.96 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_81 N_A1_c_82_n N_A2_M1004_g 0.0195161f $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_82 N_A1_c_84_n N_A2_M1004_g 0.00742259f $X=0.96 $Y=1.475 $X2=0 $Y2=0
cc_83 A1 A2 0.0288692f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_84 N_A1_c_84_n A2 2.56292e-19 $X=0.96 $Y=1.475 $X2=0 $Y2=0
cc_85 A1 N_A2_c_133_n 0.00490735f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_86 N_A1_c_84_n N_A2_c_133_n 0.00868664f $X=0.96 $Y=1.475 $X2=0 $Y2=0
cc_87 A1 N_A_28_368#_c_307_n 0.021684f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_88 N_A1_c_85_n N_A_28_368#_c_308_n 0.0043207f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A1_c_85_n N_A_28_368#_c_313_n 0.0126853f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A1_c_86_n N_A_28_368#_c_313_n 0.0120074f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_91 A1 N_A_28_368#_c_313_n 0.0435529f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_92 N_A1_c_84_n N_A_28_368#_c_313_n 0.00132059f $X=0.96 $Y=1.475 $X2=0 $Y2=0
cc_93 N_A1_c_85_n N_A_28_368#_c_309_n 6.69308e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A1_c_86_n N_A_28_368#_c_309_n 0.0105394f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A1_c_86_n N_A_28_368#_c_319_n 4.27055e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_96 A1 N_A_28_368#_c_319_n 0.021711f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_97 N_A1_c_85_n N_VPWR_c_350_n 0.0135832f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A1_c_86_n N_VPWR_c_350_n 0.00526215f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A1_c_86_n N_VPWR_c_352_n 0.00445602f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A1_c_85_n N_VPWR_c_354_n 0.00413917f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_101 N_A1_c_85_n N_VPWR_c_349_n 0.00821237f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A1_c_86_n N_VPWR_c_349_n 0.00857673f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A1_M1012_g N_A_27_74#_c_502_n 0.0104846f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A1_c_82_n N_A_27_74#_c_502_n 6.72835e-19 $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_105 N_A1_M1012_g N_A_27_74#_c_503_n 0.0118691f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A1_c_82_n N_A_27_74#_c_503_n 0.0115835f $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_107 A1 N_A_27_74#_c_503_n 0.0506639f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A1_c_84_n N_A_27_74#_c_503_n 0.0104337f $X=0.96 $Y=1.475 $X2=0 $Y2=0
cc_109 N_A1_M1012_g N_A_27_74#_c_504_n 0.00214722f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_110 A1 N_A_27_74#_c_504_n 0.0286342f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_111 N_A1_M1012_g N_A_27_74#_c_505_n 6.72835e-19 $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A1_c_82_n N_A_27_74#_c_505_n 0.00981147f $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_113 N_A1_c_82_n N_A_27_74#_c_510_n 0.0014252f $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_114 A1 N_A_27_74#_c_510_n 0.0179197f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_115 N_A1_M1012_g N_VGND_c_583_n 0.00613492f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A1_c_82_n N_VGND_c_583_n 0.00475299f $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_117 N_A1_c_82_n N_VGND_c_584_n 0.00434272f $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_118 N_A1_M1012_g N_VGND_c_586_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_119 N_A1_M1012_g N_VGND_c_588_n 0.00824951f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A1_c_82_n N_VGND_c_588_n 0.00821391f $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_121 N_A2_M1011_g N_A3_M1001_g 0.0130706f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_122 A2 N_A3_c_187_n 0.00174805f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A2_c_133_n N_A3_c_187_n 0.0130706f $X=1.86 $Y=1.557 $X2=0 $Y2=0
cc_124 A2 N_A3_c_190_n 0.0014638f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A2_c_134_n N_A_28_368#_c_309_n 0.0103267f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A2_c_135_n N_A_28_368#_c_309_n 6.54425e-19 $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A2_c_134_n N_A_28_368#_c_323_n 0.0158599f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_128 N_A2_c_135_n N_A_28_368#_c_323_n 0.0120074f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_129 A2 N_A_28_368#_c_323_n 0.0252692f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_130 N_A2_c_133_n N_A_28_368#_c_323_n 0.00301034f $X=1.86 $Y=1.557 $X2=0 $Y2=0
cc_131 N_A2_c_134_n N_A_28_368#_c_319_n 8.9215e-19 $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_132 N_A2_c_134_n N_A_28_368#_c_310_n 5.7112e-19 $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A2_c_135_n N_A_28_368#_c_310_n 0.00941736f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_134 A2 N_A_28_368#_c_310_n 0.026501f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_135 N_A2_c_133_n N_A_28_368#_c_310_n 7.32687e-19 $X=1.86 $Y=1.557 $X2=0 $Y2=0
cc_136 N_A2_c_134_n N_VPWR_c_352_n 0.00445602f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A2_c_135_n N_VPWR_c_352_n 0.00278271f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A2_c_134_n N_VPWR_c_349_n 0.00858435f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A2_c_135_n N_VPWR_c_349_n 0.00358624f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A2_c_135_n N_A_297_368#_c_398_n 0.0144245f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A2_c_134_n N_A_297_368#_c_399_n 0.00341066f $X=1.41 $Y=1.765 $X2=0
+ $Y2=0
cc_142 N_A2_c_135_n N_Y_c_430_n 0.00432247f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_143 A2 N_Y_c_426_n 0.0198017f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_144 N_A2_M1004_g N_A_27_74#_c_505_n 0.00981147f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A2_M1011_g N_A_27_74#_c_505_n 6.72835e-19 $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A2_M1004_g N_A_27_74#_c_506_n 0.015337f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A2_M1011_g N_A_27_74#_c_506_n 0.0134273f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_148 A2 N_A_27_74#_c_506_n 0.0558786f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_149 N_A2_c_133_n N_A_27_74#_c_506_n 0.00591614f $X=1.86 $Y=1.557 $X2=0 $Y2=0
cc_150 N_A2_M1011_g N_A_27_74#_c_530_n 0.00342095f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A2_M1004_g N_A_27_74#_c_510_n 0.00249368f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A2_c_133_n N_A_27_74#_c_510_n 0.00373746f $X=1.86 $Y=1.557 $X2=0 $Y2=0
cc_153 N_A2_M1004_g N_A_27_74#_c_511_n 6.72158e-19 $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A2_M1011_g N_A_27_74#_c_511_n 0.00637016f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A2_M1004_g N_VGND_c_584_n 0.00434272f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A2_M1004_g N_VGND_c_585_n 0.00475299f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A2_M1011_g N_VGND_c_585_n 0.00613492f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A2_M1004_g N_VGND_c_588_n 0.00821391f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A2_M1011_g N_VGND_c_588_n 0.00821391f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A2_M1011_g N_VGND_c_591_n 0.00434272f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A3_M1002_g N_B1_M1007_g 0.0307304f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A3_c_192_n N_B1_c_256_n 0.0234262f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A3_c_189_n N_B1_c_256_n 2.96261e-19 $X=3.28 $Y=1.515 $X2=0 $Y2=0
cc_164 N_A3_c_189_n N_B1_c_253_n 0.0203452f $X=3.28 $Y=1.515 $X2=0 $Y2=0
cc_165 N_A3_c_190_n N_B1_c_253_n 4.12636e-19 $X=3.345 $Y=1.557 $X2=0 $Y2=0
cc_166 N_A3_M1002_g N_B1_c_255_n 0.021601f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A3_c_189_n N_B1_c_255_n 0.00225382f $X=3.28 $Y=1.515 $X2=0 $Y2=0
cc_168 N_A3_c_190_n N_B1_c_255_n 0.00301396f $X=3.345 $Y=1.557 $X2=0 $Y2=0
cc_169 N_A3_c_191_n N_VPWR_c_352_n 0.00278257f $X=2.895 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A3_c_192_n N_VPWR_c_352_n 0.0044313f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A3_c_191_n N_VPWR_c_349_n 0.00358623f $X=2.895 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A3_c_192_n N_VPWR_c_349_n 0.00854637f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_173 N_A3_c_191_n N_A_297_368#_c_398_n 0.0145139f $X=2.895 $Y=1.765 $X2=0
+ $Y2=0
cc_174 N_A3_c_192_n N_A_297_368#_c_398_n 0.00416253f $X=3.345 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_A3_c_191_n N_A_297_368#_c_404_n 0.0121561f $X=2.895 $Y=1.765 $X2=0
+ $Y2=0
cc_176 N_A3_c_192_n N_A_297_368#_c_404_n 0.00604065f $X=3.345 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_A3_c_191_n N_Y_c_427_n 0.00881943f $X=2.895 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A3_M1002_g N_Y_c_424_n 0.0123777f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A3_c_189_n N_Y_c_424_n 0.0331911f $X=3.28 $Y=1.515 $X2=0 $Y2=0
cc_180 N_A3_c_190_n N_Y_c_424_n 0.0114012f $X=3.345 $Y=1.557 $X2=0 $Y2=0
cc_181 N_A3_M1001_g N_Y_c_425_n 0.00388066f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A3_c_191_n N_Y_c_440_n 0.0160674f $X=2.895 $Y=1.765 $X2=0 $Y2=0
cc_183 N_A3_c_192_n N_Y_c_440_n 0.0150982f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A3_c_189_n N_Y_c_440_n 0.0302663f $X=3.28 $Y=1.515 $X2=0 $Y2=0
cc_185 N_A3_c_190_n N_Y_c_440_n 0.00124412f $X=3.345 $Y=1.557 $X2=0 $Y2=0
cc_186 N_A3_M1002_g N_Y_c_444_n 9.17327e-19 $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A3_c_187_n N_Y_c_430_n 0.00650414f $X=2.57 $Y=1.425 $X2=0 $Y2=0
cc_188 N_A3_c_191_n N_Y_c_430_n 0.00411369f $X=2.895 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A3_M1001_g N_Y_c_426_n 0.00627755f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A3_c_186_n N_Y_c_426_n 0.0104157f $X=2.805 $Y=1.425 $X2=0 $Y2=0
cc_191 N_A3_c_191_n N_Y_c_426_n 0.00171554f $X=2.895 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A3_c_192_n N_Y_c_426_n 8.24949e-19 $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_193 N_A3_M1002_g N_Y_c_426_n 0.00426386f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A3_c_189_n N_Y_c_426_n 0.0318332f $X=3.28 $Y=1.515 $X2=0 $Y2=0
cc_195 N_A3_c_190_n N_Y_c_426_n 0.0118594f $X=3.345 $Y=1.557 $X2=0 $Y2=0
cc_196 N_A3_c_192_n N_Y_c_454_n 0.00274322f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_197 N_A3_c_192_n Y 0.00464012f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A3_M1001_g N_A_27_74#_c_506_n 0.0040258f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A3_M1001_g N_A_27_74#_c_530_n 0.00728117f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A3_M1001_g N_A_27_74#_c_537_n 0.0147088f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A3_c_186_n N_A_27_74#_c_537_n 7.0816e-19 $X=2.805 $Y=1.425 $X2=0 $Y2=0
cc_202 N_A3_M1002_g N_A_27_74#_c_537_n 0.0117184f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A3_c_190_n N_A_27_74#_c_537_n 4.51931e-19 $X=3.345 $Y=1.557 $X2=0 $Y2=0
cc_204 N_A3_M1002_g N_A_27_74#_c_541_n 0.00793893f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A3_M1002_g N_A_27_74#_c_508_n 0.00368639f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A3_M1001_g N_A_27_74#_c_511_n 0.0111378f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A3_M1002_g N_VGND_c_587_n 0.00321293f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A3_M1001_g N_VGND_c_588_n 0.00414829f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A3_M1002_g N_VGND_c_588_n 0.00414843f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A3_M1001_g N_VGND_c_591_n 0.00324657f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A3_M1001_g N_VGND_c_592_n 0.00790404f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A3_M1002_g N_VGND_c_592_n 0.00576111f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_213 N_B1_c_256_n N_VPWR_c_351_n 0.00548829f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_214 N_B1_c_257_n N_VPWR_c_351_n 0.00548829f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_215 N_B1_c_256_n N_VPWR_c_352_n 0.00445602f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_216 N_B1_c_257_n N_VPWR_c_355_n 0.00445602f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_217 N_B1_c_256_n N_VPWR_c_349_n 0.00858104f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_218 N_B1_c_257_n N_VPWR_c_349_n 0.00861084f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_219 N_B1_c_256_n N_A_297_368#_c_398_n 4.63564e-19 $X=3.845 $Y=1.765 $X2=0
+ $Y2=0
cc_220 N_B1_M1007_g N_Y_c_424_n 0.0116769f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_221 N_B1_M1008_g N_Y_c_424_n 0.00283624f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_222 N_B1_c_253_n N_Y_c_424_n 0.0392202f $X=4.365 $Y=1.515 $X2=0 $Y2=0
cc_223 N_B1_c_255_n N_Y_c_424_n 0.0047701f $X=4.295 $Y=1.532 $X2=0 $Y2=0
cc_224 N_B1_c_256_n N_Y_c_460_n 0.0120074f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_225 N_B1_c_257_n N_Y_c_460_n 0.0119773f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_226 N_B1_c_253_n N_Y_c_460_n 0.0372249f $X=4.365 $Y=1.515 $X2=0 $Y2=0
cc_227 N_B1_c_255_n N_Y_c_460_n 0.00644128f $X=4.295 $Y=1.532 $X2=0 $Y2=0
cc_228 N_B1_M1007_g N_Y_c_444_n 0.00625675f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_229 N_B1_c_257_n N_Y_c_428_n 3.69071e-19 $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_230 N_B1_c_253_n N_Y_c_428_n 7.98247e-19 $X=4.365 $Y=1.515 $X2=0 $Y2=0
cc_231 B1 N_Y_c_428_n 0.0259797f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_232 N_B1_c_255_n N_Y_c_428_n 0.00196164f $X=4.295 $Y=1.532 $X2=0 $Y2=0
cc_233 N_B1_c_256_n N_Y_c_429_n 6.7588e-19 $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_234 N_B1_c_257_n N_Y_c_429_n 0.011911f $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_235 N_B1_c_256_n N_Y_c_454_n 0.00283991f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_236 N_B1_c_257_n N_Y_c_454_n 2.94324e-19 $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_237 N_B1_c_253_n N_Y_c_454_n 0.00565856f $X=4.365 $Y=1.515 $X2=0 $Y2=0
cc_238 N_B1_c_255_n N_Y_c_454_n 0.00164753f $X=4.295 $Y=1.532 $X2=0 $Y2=0
cc_239 N_B1_c_256_n Y 0.00959654f $X=3.845 $Y=1.765 $X2=0 $Y2=0
cc_240 N_B1_c_257_n Y 3.80626e-19 $X=4.295 $Y=1.765 $X2=0 $Y2=0
cc_241 N_B1_M1007_g N_A_27_74#_c_507_n 0.0107757f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_242 N_B1_M1008_g N_A_27_74#_c_507_n 0.0140969f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_243 N_B1_M1007_g N_A_27_74#_c_509_n 8.96536e-19 $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_244 N_B1_M1008_g N_A_27_74#_c_509_n 0.00715938f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_245 N_B1_c_253_n N_A_27_74#_c_509_n 3.7446e-19 $X=4.365 $Y=1.515 $X2=0 $Y2=0
cc_246 B1 N_A_27_74#_c_509_n 0.0260711f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_247 N_B1_c_255_n N_A_27_74#_c_509_n 0.00173045f $X=4.295 $Y=1.532 $X2=0 $Y2=0
cc_248 N_B1_M1007_g N_VGND_c_587_n 0.00278271f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_249 N_B1_M1008_g N_VGND_c_587_n 0.00278266f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_250 N_B1_M1007_g N_VGND_c_588_n 0.00354005f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_251 N_B1_M1008_g N_VGND_c_588_n 0.00357648f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_28_368#_c_313_n N_VPWR_M1005_d 0.00384138f $X=1.02 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_253 N_A_28_368#_c_308_n N_VPWR_c_350_n 0.0453479f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_254 N_A_28_368#_c_313_n N_VPWR_c_350_n 0.0154248f $X=1.02 $Y=2.035 $X2=0
+ $Y2=0
cc_255 N_A_28_368#_c_309_n N_VPWR_c_350_n 0.0462948f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_256 N_A_28_368#_c_309_n N_VPWR_c_352_n 0.014552f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_257 N_A_28_368#_c_308_n N_VPWR_c_354_n 0.011066f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_258 N_A_28_368#_c_308_n N_VPWR_c_349_n 0.00915947f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_259 N_A_28_368#_c_309_n N_VPWR_c_349_n 0.0119791f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_260 N_A_28_368#_c_323_n N_A_297_368#_M1010_d 0.004142f $X=1.92 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_261 N_A_28_368#_c_309_n N_A_297_368#_c_408_n 0.040027f $X=1.185 $Y=2.815
+ $X2=0 $Y2=0
cc_262 N_A_28_368#_c_323_n N_A_297_368#_c_408_n 0.0136682f $X=1.92 $Y=2.035
+ $X2=0 $Y2=0
cc_263 N_A_28_368#_c_310_n N_A_297_368#_c_408_n 0.0289859f $X=2.085 $Y=2.115
+ $X2=0 $Y2=0
cc_264 N_A_28_368#_M1015_s N_A_297_368#_c_398_n 0.00287371f $X=1.935 $Y=1.84
+ $X2=0 $Y2=0
cc_265 N_A_28_368#_c_310_n N_A_297_368#_c_398_n 0.0205764f $X=2.085 $Y=2.115
+ $X2=0 $Y2=0
cc_266 N_A_28_368#_c_309_n N_A_297_368#_c_399_n 0.00549849f $X=1.185 $Y=2.815
+ $X2=0 $Y2=0
cc_267 N_A_28_368#_c_310_n N_Y_c_427_n 0.0377583f $X=2.085 $Y=2.115 $X2=0 $Y2=0
cc_268 N_A_28_368#_c_310_n N_Y_c_430_n 0.0113228f $X=2.085 $Y=2.115 $X2=0 $Y2=0
cc_269 N_VPWR_c_352_n N_A_297_368#_c_398_n 0.102223f $X=3.985 $Y=3.33 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_349_n N_A_297_368#_c_398_n 0.0578213f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_352_n N_A_297_368#_c_399_n 0.0121867f $X=3.985 $Y=3.33 $X2=0
+ $Y2=0
cc_272 N_VPWR_c_349_n N_A_297_368#_c_399_n 0.00660921f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_273 N_VPWR_M1000_d N_Y_c_460_n 0.00402933f $X=3.92 $Y=1.84 $X2=0 $Y2=0
cc_274 N_VPWR_c_351_n N_Y_c_460_n 0.0136682f $X=4.07 $Y=2.355 $X2=0 $Y2=0
cc_275 N_VPWR_c_351_n N_Y_c_429_n 0.0514854f $X=4.07 $Y=2.355 $X2=0 $Y2=0
cc_276 N_VPWR_c_355_n N_Y_c_429_n 0.0145938f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_277 N_VPWR_c_349_n N_Y_c_429_n 0.0120466f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_278 N_VPWR_c_351_n Y 0.0514854f $X=4.07 $Y=2.355 $X2=0 $Y2=0
cc_279 N_VPWR_c_352_n Y 0.0145938f $X=3.985 $Y=3.33 $X2=0 $Y2=0
cc_280 N_VPWR_c_349_n Y 0.0120466f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_281 N_A_297_368#_c_398_n N_Y_M1009_s 0.00312144f $X=2.955 $Y=2.99 $X2=0 $Y2=0
cc_282 N_A_297_368#_c_398_n N_Y_c_427_n 0.018931f $X=2.955 $Y=2.99 $X2=0 $Y2=0
cc_283 N_A_297_368#_c_404_n N_Y_c_427_n 0.0298377f $X=3.12 $Y=2.455 $X2=0 $Y2=0
cc_284 N_A_297_368#_M1009_d N_Y_c_440_n 0.00359365f $X=2.97 $Y=1.84 $X2=0 $Y2=0
cc_285 N_A_297_368#_c_404_n N_Y_c_440_n 0.0171813f $X=3.12 $Y=2.455 $X2=0 $Y2=0
cc_286 N_A_297_368#_c_398_n Y 0.00395311f $X=2.955 $Y=2.99 $X2=0 $Y2=0
cc_287 N_Y_c_424_n N_A_27_74#_M1002_s 0.00176461f $X=3.85 $Y=1.095 $X2=0 $Y2=0
cc_288 N_Y_c_425_n N_A_27_74#_c_506_n 0.012289f $X=2.835 $Y=1.095 $X2=0 $Y2=0
cc_289 N_Y_c_424_n N_A_27_74#_c_537_n 0.0528952f $X=3.85 $Y=1.095 $X2=0 $Y2=0
cc_290 N_Y_c_425_n N_A_27_74#_c_537_n 0.013831f $X=2.835 $Y=1.095 $X2=0 $Y2=0
cc_291 N_Y_M1007_d N_A_27_74#_c_507_n 0.00237956f $X=3.875 $Y=0.37 $X2=0 $Y2=0
cc_292 N_Y_c_424_n N_A_27_74#_c_507_n 0.0030313f $X=3.85 $Y=1.095 $X2=0 $Y2=0
cc_293 N_Y_c_444_n N_A_27_74#_c_507_n 0.0166105f $X=4.015 $Y=0.775 $X2=0 $Y2=0
cc_294 N_Y_c_424_n N_VGND_M1001_d 0.00581259f $X=3.85 $Y=1.095 $X2=0 $Y2=0
cc_295 N_Y_c_425_n N_VGND_M1001_d 0.00372663f $X=2.835 $Y=1.095 $X2=0 $Y2=0
cc_296 N_A_27_74#_c_503_n N_VGND_M1012_d 0.00369983f $X=1.115 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_297 N_A_27_74#_c_506_n N_VGND_M1004_d 0.00369983f $X=2.115 $Y=1.095 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_c_537_n N_VGND_M1001_d 0.0164865f $X=3.42 $Y=0.755 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_502_n N_VGND_c_583_n 0.0186136f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_503_n N_VGND_c_583_n 0.0233713f $X=1.115 $Y=1.095 $X2=0
+ $Y2=0
cc_301 N_A_27_74#_c_505_n N_VGND_c_583_n 0.0186136f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_302 N_A_27_74#_c_505_n N_VGND_c_584_n 0.0144922f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_303 N_A_27_74#_c_505_n N_VGND_c_585_n 0.0186136f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_304 N_A_27_74#_c_506_n N_VGND_c_585_n 0.0233713f $X=2.115 $Y=1.095 $X2=0
+ $Y2=0
cc_305 N_A_27_74#_c_511_n N_VGND_c_585_n 0.0186136f $X=2.28 $Y=0.515 $X2=0 $Y2=0
cc_306 N_A_27_74#_c_502_n N_VGND_c_586_n 0.0145639f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_307 N_A_27_74#_c_537_n N_VGND_c_587_n 0.00236055f $X=3.42 $Y=0.755 $X2=0
+ $Y2=0
cc_308 N_A_27_74#_c_507_n N_VGND_c_587_n 0.0665294f $X=4.35 $Y=0.34 $X2=0 $Y2=0
cc_309 N_A_27_74#_c_508_n N_VGND_c_587_n 0.0176331f $X=3.67 $Y=0.34 $X2=0 $Y2=0
cc_310 N_A_27_74#_c_502_n N_VGND_c_588_n 0.0119984f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_311 N_A_27_74#_c_505_n N_VGND_c_588_n 0.0118826f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_312 N_A_27_74#_c_537_n N_VGND_c_588_n 0.0113479f $X=3.42 $Y=0.755 $X2=0 $Y2=0
cc_313 N_A_27_74#_c_507_n N_VGND_c_588_n 0.0370234f $X=4.35 $Y=0.34 $X2=0 $Y2=0
cc_314 N_A_27_74#_c_508_n N_VGND_c_588_n 0.00956698f $X=3.67 $Y=0.34 $X2=0 $Y2=0
cc_315 N_A_27_74#_c_511_n N_VGND_c_588_n 0.0118826f $X=2.28 $Y=0.515 $X2=0 $Y2=0
cc_316 N_A_27_74#_c_537_n N_VGND_c_591_n 0.0023667f $X=3.42 $Y=0.755 $X2=0 $Y2=0
cc_317 N_A_27_74#_c_511_n N_VGND_c_591_n 0.0144922f $X=2.28 $Y=0.515 $X2=0 $Y2=0
cc_318 N_A_27_74#_c_537_n N_VGND_c_592_n 0.0468302f $X=3.42 $Y=0.755 $X2=0 $Y2=0
cc_319 N_A_27_74#_c_508_n N_VGND_c_592_n 0.0119157f $X=3.67 $Y=0.34 $X2=0 $Y2=0
cc_320 N_A_27_74#_c_511_n N_VGND_c_592_n 0.00620201f $X=2.28 $Y=0.515 $X2=0
+ $Y2=0
