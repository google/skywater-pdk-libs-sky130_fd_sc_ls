* NGSPICE file created from sky130_fd_sc_ls__nand4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
M1000 a_374_74# a_27_114# Y VNB nshort w=740000u l=150000u
+  ad=1.0508e+12p pd=1.024e+07u as=4.921e+11p ps=4.29e+06u
M1001 VPWR B_N a_232_114# VPB phighvt w=840000u l=150000u
+  ad=3.9592e+12p pd=3.104e+07u as=2.52e+11p ps=2.28e+06u
M1002 a_828_74# a_232_114# a_374_74# VNB nshort w=740000u l=150000u
+  ad=9.53e+11p pd=8.52e+06u as=0p ps=0u
M1003 a_1229_74# D VGND VNB nshort w=740000u l=150000u
+  ad=1.0434e+12p pd=1.022e+07u as=9.049e+11p ps=7.36e+06u
M1004 VPWR a_232_114# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=2.744e+12p ps=2.282e+07u
M1005 Y a_27_114# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_27_114# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_374_74# a_27_114# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y D VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_374_74# a_232_114# a_828_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND D a_1229_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y a_27_114# a_374_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND D a_1229_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_27_114# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y C VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_27_114# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR D Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_828_74# a_232_114# a_374_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A_N a_27_114# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1019 VPWR C Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_232_114# B_N VGND VNB nshort w=740000u l=150000u
+  ad=2.368e+11p pd=2.12e+06u as=0p ps=0u
M1021 a_828_74# C a_1229_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y a_232_114# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_828_74# C a_1229_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A_N a_27_114# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.52e+11p ps=2.28e+06u
M1025 Y D VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_114# A_N VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y C VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_374_74# a_232_114# a_828_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y a_27_114# a_374_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_232_114# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR D Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1229_74# D VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_232_114# B_N VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Y a_232_114# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1229_74# C a_828_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1229_74# C a_828_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR C Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

