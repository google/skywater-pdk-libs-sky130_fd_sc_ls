* File: sky130_fd_sc_ls__edfxbp_1.spice
* Created: Fri Aug 28 13:22:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__edfxbp_1.pex.spice"
.subckt sky130_fd_sc_ls__edfxbp_1  VNB VPB D DE CLK VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* CLK	CLK
* DE	DE
* D	D
* VPB	VPB
* VNB	VNB
MM1031 A_145_74# N_D_M1031_g N_A_27_74#_M1031_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1848 PD=0.66 PS=1.72 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_DE_M1017_g A_145_74# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.8 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_DE_M1026_g N_A_161_446#_M1026_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.1281 PD=0.78 PS=1.45 NRD=19.992 NRS=2.856 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1034 A_527_74# N_A_161_446#_M1034_g N_VGND_M1026_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=2.856 M=1 R=2.8 SA=75000.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1035 N_A_27_74#_M1035_d N_A_575_48#_M1035_g A_527_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1027 N_A_818_74#_M1027_d N_CLK_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.2109 PD=2.01 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1028 N_A_1008_74#_M1028_d N_A_818_74#_M1028_g N_VGND_M1028_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1961 AS=0.1961 PD=2.01 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1033 N_A_1198_97#_M1033_d N_A_818_74#_M1033_g N_A_27_74#_M1033_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=0.95 PS=1.37 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1012 A_1334_97# N_A_1008_74#_M1012_g N_A_1198_97#_M1033_d VNB NSHORT L=0.15
+ W=0.42 AD=0.08925 AS=0.1113 PD=0.845 PS=0.95 NRD=45 NRS=0 M=1 R=2.8 SA=75000.9
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_1419_71#_M1019_g A_1334_97# VNB NSHORT L=0.15 W=0.42
+ AD=0.109992 AS=0.08925 PD=0.92717 PS=0.845 NRD=0 NRS=45 M=1 R=2.8 SA=75001.4
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1013 N_A_1419_71#_M1013_d N_A_1198_97#_M1013_g N_VGND_M1019_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.167608 PD=1.85 PS=1.41283 NRD=0 NRS=46.872 M=1
+ R=4.26667 SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 A_1807_74# N_A_1419_71#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.0777 AS=0.2109 PD=0.95 PS=2.05 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1006 N_A_1879_74#_M1006_d N_A_1008_74#_M1006_g A_1807_74# VNB NSHORT L=0.15
+ W=0.74 AD=0.477045 AS=0.0777 PD=2.97276 PS=0.95 NRD=14.592 NRS=8.1 M=1
+ R=4.93333 SA=75000.6 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1025 A_2227_118# N_A_818_74#_M1025_g N_A_1879_74#_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.270755 PD=0.66 PS=1.68724 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75002.3 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_575_48#_M1009_g A_2227_118# VNB NSHORT L=0.15 W=0.42
+ AD=0.114985 AS=0.0504 PD=0.907358 PS=0.66 NRD=45 NRS=18.564 M=1 R=2.8
+ SA=75002.7 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1014 N_A_575_48#_M1014_d N_A_1879_74#_M1014_g N_VGND_M1009_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1824 AS=0.175215 PD=1.85 PS=1.38264 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75002.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1015 N_VGND_M1015_d N_A_1879_74#_M1015_g N_Q_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2257 AS=0.2109 PD=1.35 PS=2.05 NRD=53.508 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001 A=0.111 P=1.78 MULT=1
MM1020 N_Q_N_M1020_d N_A_575_48#_M1020_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.2257 PD=2.05 PS=1.35 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1024 A_116_508# N_D_M1024_g N_A_27_74#_M1024_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1239 PD=0.66 PS=1.43 NRD=30.4759 NRS=4.6886 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1029 N_VPWR_M1029_d N_A_161_446#_M1029_g A_116_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1239 AS=0.0504 PD=1.43 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1032 N_VPWR_M1032_d N_DE_M1032_g N_A_161_446#_M1032_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1888 PD=1.41283 PS=1.87 NRD=73.8553 NRS=3.0732 M=1
+ R=4.26667 SA=75000.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1030 A_556_504# N_DE_M1030_g N_VPWR_M1032_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1113 PD=0.66 PS=0.92717 NRD=30.4759 NRS=4.6886 M=1 R=2.8
+ SA=75000.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_27_74#_M1007_d N_A_575_48#_M1007_g A_556_504# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1239 AS=0.0504 PD=1.43 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.8
+ SA=75001.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_A_818_74#_M1008_d N_CLK_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1003 N_A_1008_74#_M1003_d N_A_818_74#_M1003_g N_VPWR_M1003_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1010 N_A_1198_97#_M1010_d N_A_1008_74#_M1010_g N_A_27_74#_M1010_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.063 AS=0.206 PD=0.72 PS=1.92 NRD=4.6886 NRS=46.886 M=1
+ R=2.8 SA=75000.3 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1001 A_1423_508# N_A_818_74#_M1001_g N_A_1198_97#_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0756 AS=0.063 PD=0.78 PS=0.72 NRD=58.6272 NRS=4.6886 M=1 R=2.8
+ SA=75000.8 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_1419_71#_M1004_g A_1423_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.125617 AS=0.0756 PD=1.03 PS=0.78 NRD=114.477 NRS=58.6272 M=1 R=2.8
+ SA=75001.3 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1016 N_A_1419_71#_M1016_d N_A_1198_97#_M1016_g N_VPWR_M1004_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2478 AS=0.251233 PD=2.27 PS=2.06 NRD=2.3443 NRS=57.2285 M=1
+ R=5.6 SA=75001 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 A_2008_392# N_A_1419_71#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1021 N_A_1879_74#_M1021_d N_A_818_74#_M1021_g A_2008_392# VPB PHIGHVT L=0.15
+ W=1 AD=0.244718 AS=0.135 PD=2 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75000.6 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1018 A_2206_443# N_A_1008_74#_M1018_g N_A_1879_74#_M1021_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0693 AS=0.102782 PD=0.75 PS=0.84 NRD=51.5943 NRS=60.9715 M=1 R=2.8
+ SA=75001.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_575_48#_M1000_g A_2206_443# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.145462 AS=0.0693 PD=1.06775 PS=0.75 NRD=4.6886 NRS=51.5943 M=1 R=2.8
+ SA=75001.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1023 N_A_575_48#_M1023_d N_A_1879_74#_M1023_g N_VPWR_M1000_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.346338 PD=2.59 PS=2.54225 NRD=1.9503 NRS=11.8003 M=1
+ R=6.66667 SA=75001.2 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_A_1879_74#_M1011_g N_Q_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1022 N_Q_N_M1022_d N_A_575_48#_M1022_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX36_noxref VNB VPB NWDIODE A=27.5178 P=33.33
*
.include "sky130_fd_sc_ls__edfxbp_1.pxi.spice"
*
.ends
*
*
