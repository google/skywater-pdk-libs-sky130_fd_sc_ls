* File: sky130_fd_sc_ls__sdfrbp_1.spice
* Created: Wed Sep  2 11:26:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sdfrbp_1.pex.spice"
.subckt sky130_fd_sc_ls__sdfrbp_1  VNB VPB SCE D SCD CLK RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1032 N_VGND_M1032_d N_SCE_M1032_g N_A_27_74#_M1032_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 noxref_26 N_A_27_74#_M1008_g N_noxref_25_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.1197 PD=0.755 PS=1.41 NRD=32.136 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1012 N_A_409_81#_M1012_d N_D_M1012_g noxref_26 VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.07035 PD=0.95 PS=0.755 NRD=71.424 NRS=32.136 M=1 R=2.8
+ SA=75000.7 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1022 noxref_27 N_SCE_M1022_g N_A_409_81#_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1113 PD=0.66 PS=0.95 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1016 N_noxref_25_M1016_d N_SCD_M1016_g noxref_27 VNB NSHORT L=0.15 W=0.42
+ AD=0.0651 AS=0.0504 PD=0.73 PS=0.66 NRD=2.856 NRS=18.564 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_RESET_B_M1036_g N_noxref_25_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0651 PD=1.41 PS=0.73 NRD=0 NRS=5.712 M=1 R=2.8
+ SA=75002.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_CLK_M1025_g N_A_835_98#_M1025_s VNB NSHORT L=0.15 W=0.74
+ AD=0.167375 AS=0.2619 PD=1.295 PS=2.38 NRD=10.536 NRS=10.536 M=1 R=4.93333
+ SA=75000.2 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1033 N_A_1034_392#_M1033_d N_A_835_98#_M1033_g N_VGND_M1025_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.1961 AS=0.167375 PD=2.01 PS=1.295 NRD=0 NRS=10.536 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1035 N_A_1234_119#_M1035_d N_A_835_98#_M1035_g N_A_409_81#_M1035_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1000 A_1320_119# N_A_1034_392#_M1000_g N_A_1234_119#_M1035_d VNB NSHORT L=0.15
+ W=0.42 AD=0.04935 AS=0.0588 PD=0.655 PS=0.7 NRD=17.856 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1021 A_1397_119# N_A_1367_93#_M1021_g A_1320_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.04935 PD=0.66 PS=0.655 NRD=18.564 NRS=17.856 M=1 R=2.8 SA=75001
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_RESET_B_M1011_g A_1397_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.211199 AS=0.0504 PD=1.27189 PS=0.66 NRD=127.956 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1030 N_A_1367_93#_M1030_d N_A_1234_119#_M1030_g N_VGND_M1011_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0928 AS=0.321826 PD=0.93 PS=1.93811 NRD=0 NRS=83.964 M=1
+ R=4.26667 SA=75001.7 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1020 N_A_1747_74#_M1020_d N_A_1034_392#_M1020_g N_A_1367_93#_M1030_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.272845 AS=0.0928 PD=1.91396 PS=0.93 NRD=92.808 NRS=0
+ M=1 R=4.26667 SA=75002.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1009 A_1966_74# N_A_835_98#_M1009_g N_A_1747_74#_M1020_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.179055 PD=0.63 PS=1.25604 NRD=14.28 NRS=48.564 M=1 R=2.8
+ SA=75002.9 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_2008_48#_M1003_g A_1966_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1005 A_2124_74# N_RESET_B_M1005_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_2008_48#_M1007_d N_A_1747_74#_M1007_g A_2124_74# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_Q_N_M1006_d N_A_1747_74#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2072 AS=0.3159 PD=2.04 PS=2.57 NRD=0 NRS=60.3 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A_1747_74#_M1001_g N_A_2513_424#_M1001_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.101196 AS=0.14575 PD=0.92093 PS=1.63 NRD=13.632 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1031 N_Q_M1031_d N_A_2513_424#_M1031_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.136154 PD=2.05 PS=1.23907 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1026 N_VPWR_M1026_d N_SCE_M1026_g N_A_27_74#_M1026_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.112 AS=0.5792 PD=0.99 PS=3.09 NRD=18.4589 NRS=3.0732 M=1 R=4.26667
+ SA=75000.8 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1037 A_338_464# N_SCE_M1037_g N_VPWR_M1026_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.112 PD=0.91 PS=0.99 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75001.3 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1014 N_A_409_81#_M1014_d N_D_M1014_g A_338_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.096 AS=0.0864 PD=0.94 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75001.8 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1019 A_512_464# N_A_27_74#_M1019_g N_A_409_81#_M1014_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.128 AS=0.096 PD=1.04 PS=0.94 NRD=44.6205 NRS=3.0732 M=1 R=4.26667
+ SA=75002.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1023 N_VPWR_M1023_d N_SCD_M1023_g A_512_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1344 AS=0.128 PD=1.06 PS=1.04 NRD=3.0732 NRS=44.6205 M=1 R=4.26667
+ SA=75002.8 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1038 N_A_409_81#_M1038_d N_RESET_B_M1038_g N_VPWR_M1023_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1888 AS=0.1344 PD=1.87 PS=1.06 NRD=3.0732 NRS=40.0107 M=1
+ R=4.26667 SA=75003.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1024 N_VPWR_M1024_d N_CLK_M1024_g N_A_835_98#_M1024_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1028 N_A_1034_392#_M1028_d N_A_835_98#_M1028_g N_VPWR_M1024_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1039 N_A_1234_119#_M1039_d N_A_1034_392#_M1039_g N_A_409_81#_M1039_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.063 AS=0.1239 PD=0.72 PS=1.43 NRD=4.6886 NRS=4.6886
+ M=1 R=2.8 SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1010 A_1332_457# N_A_835_98#_M1010_g N_A_1234_119#_M1039_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.063 PD=0.63 PS=0.72 NRD=23.443 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001 A=0.063 P=1.14 MULT=1
MM1034 N_VPWR_M1034_d N_A_1367_93#_M1034_g A_1332_457# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.063 AS=0.0441 PD=0.72 PS=0.63 NRD=4.6886 NRS=23.443 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1004 N_A_1234_119#_M1004_d N_RESET_B_M1004_g N_VPWR_M1034_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1239 AS=0.063 PD=1.43 PS=0.72 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75001.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1040 N_A_1367_93#_M1040_d N_A_1234_119#_M1040_g N_VPWR_M1040_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.285 PD=1.3 PS=2.57 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1013 N_A_1747_74#_M1013_d N_A_835_98#_M1013_g N_A_1367_93#_M1040_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.292148 AS=0.15 PD=2.47183 PS=1.3 NRD=23.3051 NRS=1.9503 M=1
+ R=6.66667 SA=75000.7 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1015 A_1969_489# N_A_1034_392#_M1015_g N_A_1747_74#_M1013_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.122702 PD=0.66 PS=1.03817 NRD=30.4759 NRS=4.6886 M=1
+ R=2.8 SA=75001.1 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1017 N_VPWR_M1017_d N_A_2008_48#_M1017_g A_1969_489# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.117862 AS=0.0504 PD=1.01 PS=0.66 NRD=49.2303 NRS=30.4759 M=1 R=2.8
+ SA=75001.4 SB=75002 A=0.063 P=1.14 MULT=1
MM1027 N_A_2008_48#_M1027_d N_RESET_B_M1027_g N_VPWR_M1017_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.063 AS=0.117862 PD=0.72 PS=1.01 NRD=4.6886 NRS=51.5943 M=1 R=2.8
+ SA=75002.1 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1041 N_VPWR_M1041_d N_A_1747_74#_M1041_g N_A_2008_48#_M1027_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.121609 AS=0.063 PD=0.9 PS=0.72 NRD=75.0373 NRS=4.6886 M=1
+ R=2.8 SA=75002.5 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1002 N_Q_N_M1002_d N_A_1747_74#_M1002_g N_VPWR_M1041_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.324291 PD=2.83 PS=2.4 NRD=1.7533 NRS=12.017 M=1
+ R=7.46667 SA=75001.4 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1029 N_VPWR_M1029_d N_A_1747_74#_M1029_g N_A_2513_424#_M1029_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1662 AS=0.231 PD=1.27714 PS=2.23 NRD=10.5395 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1018 N_Q_M1018_d N_A_2513_424#_M1018_g N_VPWR_M1029_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.308 AS=0.2216 PD=2.79 PS=1.70286 NRD=1.7533 NRS=5.8509 M=1
+ R=7.46667 SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX42_noxref VNB VPB NWDIODE A=26.7346 P=32.56
c_154 VNB 0 1.61901e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__sdfrbp_1.pxi.spice"
*
.ends
*
*
