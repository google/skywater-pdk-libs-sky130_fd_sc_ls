* NGSPICE file created from sky130_fd_sc_ls__dlxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
M1000 a_664_392# a_231_74# a_586_392# VPB phighvt w=1e+06u l=150000u
+  ad=3.278e+11p pd=2.76e+06u as=2.4e+11p ps=2.48e+06u
M1001 a_231_74# GATE VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.4685e+12p ps=1.184e+07u
M1002 a_815_124# a_231_74# a_664_392# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.028e+11p ps=2.46e+06u
M1003 VGND D a_27_413# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1004 Q_N a_1347_424# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.248e+11p pd=2.82e+06u as=2.07525e+12p ps=1.551e+07u
M1005 a_770_508# a_373_82# a_664_392# VPB phighvt w=420000u l=150000u
+  ad=2.121e+11p pd=1.85e+06u as=0p ps=0u
M1006 a_863_98# a_664_392# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1007 VPWR a_863_98# a_770_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Q_N a_1347_424# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1009 a_664_392# a_373_82# a_589_80# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1010 a_589_80# a_27_413# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_863_98# a_664_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1012 a_586_392# a_27_413# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_863_98# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1014 VPWR a_231_74# a_373_82# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1015 a_1347_424# a_863_98# VGND VNB nshort w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1016 VGND a_231_74# a_373_82# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1017 VPWR D a_27_413# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.436e+11p ps=2.26e+06u
M1018 VGND a_863_98# a_815_124# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_863_98# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1020 a_1347_424# a_863_98# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.436e+11p pd=2.26e+06u as=0p ps=0u
M1021 a_231_74# GATE VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
.ends

