* NGSPICE file created from sky130_fd_sc_ls__o21a_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_376_387# VPB phighvt w=1e+06u l=150000u
+  ad=9.6465e+11p pd=6.12e+06u as=4.2e+11p ps=2.84e+06u
M1001 a_320_74# A1 VGND VNB nshort w=640000u l=150000u
+  ad=3.616e+11p pd=3.69e+06u as=3.901e+11p ps=3.89e+06u
M1002 a_320_74# B1 a_83_244# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1003 a_83_244# B1 VPWR VPB phighvt w=840000u l=150000u
+  ad=3.406e+11p pd=2.71e+06u as=0p ps=0u
M1004 a_376_387# A2 a_83_244# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_83_244# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1006 VGND a_83_244# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1007 VGND A2 a_320_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

