* File: sky130_fd_sc_ls__sdfstp_2.spice
* Created: Fri Aug 28 14:04:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__sdfstp_2.pex.spice"
.subckt sky130_fd_sc_ls__sdfstp_2  VNB VPB SCE D SCD CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1039 N_VGND_M1039_d N_SCE_M1039_g N_A_27_74#_M1039_s VNB NSHORT L=0.15 W=0.42
+ AD=0.09975 AS=0.1197 PD=0.895 PS=1.41 NRD=37.14 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1031 A_239_74# N_A_27_74#_M1031_g N_VGND_M1039_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.09975 PD=0.66 PS=0.895 NRD=18.564 NRS=18.564 M=1 R=2.8
+ SA=75000.8 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1013 N_A_290_464#_M1013_d N_D_M1013_g A_239_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1032 A_403_74# N_SCE_M1032_g N_A_290_464#_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_SCD_M1026_g A_403_74# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0672 PD=1.41 PS=0.74 NRD=0 NRS=30 M=1 R=2.8 SA=75002.1 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_CLK_M1002_g N_A_608_74#_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1000 N_A_795_74#_M1000_d N_A_608_74#_M1000_g N_VGND_M1002_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2072 AS=0.1295 PD=2.04 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_991_81#_M1008_d N_A_608_74#_M1008_g N_A_290_464#_M1008_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1281 AS=0.1176 PD=1.03 PS=1.4 NRD=94.284 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1020 A_1143_81# N_A_795_74#_M1020_g N_A_991_81#_M1008_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1281 PD=0.63 PS=1.03 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_1185_55#_M1006_g A_1143_81# VNB NSHORT L=0.15 W=0.42
+ AD=0.2316 AS=0.0441 PD=2.11 PS=0.63 NRD=141.828 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1011 A_1429_74# N_A_991_81#_M1011_g N_A_1185_55#_M1011_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_SET_B_M1012_g A_1429_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.108328 AS=0.0504 PD=0.919245 PS=0.66 NRD=24.276 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1014 N_A_1641_74#_M1014_d N_A_991_81#_M1014_g N_VGND_M1012_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.165072 PD=0.92 PS=1.40075 NRD=0 NRS=29.052 M=1 R=4.26667
+ SA=75000.9 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1025 N_A_1641_74#_M1014_d N_A_991_81#_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.2336 PD=0.92 PS=2.01 NRD=0 NRS=14.988 M=1 R=4.26667
+ SA=75001.3 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1028 N_A_1641_74#_M1028_d N_A_795_74#_M1028_g N_A_1804_424#_M1028_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.2272 PD=0.92 PS=1.99 NRD=0 NRS=13.116 M=1
+ R=4.26667 SA=75000.3 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1042 N_A_1641_74#_M1028_d N_A_795_74#_M1042_g N_A_1804_424#_M1042_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.121962 PD=0.92 PS=1.19547 NRD=0 NRS=13.116 M=1
+ R=4.26667 SA=75000.7 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1040 A_2141_74# N_A_608_74#_M1040_g N_A_1804_424#_M1042_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0800377 PD=0.66 PS=0.784528 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75001.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1038 A_2219_74# N_A_2186_367#_M1038_g A_2141_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0504 PD=0.84 PS=0.66 NRD=44.28 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_SET_B_M1009_g A_2219_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.14385 AS=0.0882 PD=1.105 PS=0.84 NRD=0 NRS=44.28 M=1 R=2.8 SA=75002.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1015 N_A_2186_367#_M1015_d N_A_1804_424#_M1015_g N_VGND_M1009_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.14385 PD=1.41 PS=1.105 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75003 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_1804_424#_M1007_g N_A_2611_98#_M1007_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.124754 AS=0.1824 PD=1.0342 PS=1.85 NRD=17.34 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1003 N_Q_M1003_d N_A_2611_98#_M1003_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.144246 PD=1.02 PS=1.1958 NRD=0 NRS=0.804 M=1 R=4.93333
+ SA=75000.7 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1029 N_Q_M1003_d N_A_2611_98#_M1029_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.222 PD=1.02 PS=2.08 NRD=0 NRS=2.424 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1021 N_VPWR_M1021_d N_SCE_M1021_g N_A_27_74#_M1021_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.096 AS=0.1888 PD=0.94 PS=1.87 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1022 A_206_464# N_SCE_M1022_g N_VPWR_M1021_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.096 PD=0.91 PS=0.94 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1010 N_A_290_464#_M1010_d N_D_M1010_g A_206_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1536 AS=0.0864 PD=1.12 PS=0.91 NRD=30.7714 NRS=24.625 M=1 R=4.26667
+ SA=75001.1 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1044 A_416_464# N_A_27_74#_M1044_g N_A_290_464#_M1010_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0864 AS=0.1536 PD=0.91 PS=1.12 NRD=24.625 NRS=30.7714 M=1
+ R=4.26667 SA=75001.7 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1034 N_VPWR_M1034_d N_SCD_M1034_g A_416_464# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.2749 AS=0.0864 PD=2.35 PS=0.91 NRD=27.6982 NRS=24.625 M=1 R=4.26667
+ SA=75002.1 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1045 N_VPWR_M1045_d N_CLK_M1045_g N_A_608_74#_M1045_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1004 N_A_795_74#_M1004_d N_A_608_74#_M1004_g N_VPWR_M1045_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3076 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1019 N_A_991_81#_M1019_d N_A_795_74#_M1019_g N_A_290_464#_M1019_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.092225 AS=0.1239 PD=0.935 PS=1.43 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1017 A_1117_483# N_A_608_74#_M1017_g N_A_991_81#_M1019_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0857 AS=0.092225 PD=0.89 PS=0.935 NRD=69.8956 NRS=46.886 M=1 R=2.8
+ SA=75000.6 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1030 N_VPWR_M1030_d N_A_1185_55#_M1030_g A_1117_483# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.11235 AS=0.0857 PD=0.955 PS=0.89 NRD=7.0329 NRS=69.8956 M=1 R=2.8
+ SA=75001 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1023 N_A_1185_55#_M1023_d N_A_991_81#_M1023_g N_VPWR_M1030_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.07245 AS=0.11235 PD=0.765 PS=0.955 NRD=4.6886 NRS=112.566
+ M=1 R=2.8 SA=75001.7 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1041 N_VPWR_M1041_d N_SET_B_M1041_g N_A_1185_55#_M1023_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.07245 PD=0.883333 PS=0.765 NRD=91.4474 NRS=25.7873 M=1
+ R=2.8 SA=75002.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1018 N_A_1584_379#_M1018_d N_A_991_81#_M1018_g N_VPWR_M1041_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.126 AS=0.2184 PD=1.14 PS=1.76667 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75001.5 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1027 N_A_1584_379#_M1018_d N_A_991_81#_M1027_g N_VPWR_M1027_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.126 AS=0.2352 PD=1.14 PS=2.24 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75002 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_A_1584_379#_M1005_d N_A_608_74#_M1005_g N_A_1804_424#_M1005_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.126 AS=0.2898 PD=1.14 PS=2.37 NRD=2.3443
+ NRS=14.0658 M=1 R=5.6 SA=75000.3 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1016 N_A_1584_379#_M1005_d N_A_608_74#_M1016_g N_A_1804_424#_M1016_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.126 AS=0.2394 PD=1.14 PS=1.90667 NRD=2.3443
+ NRS=38.6908 M=1 R=5.6 SA=75000.7 SB=75001 A=0.126 P=1.98 MULT=1
MM1024 A_2141_508# N_A_795_74#_M1024_g N_A_1804_424#_M1016_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=0.953333 NRD=30.4759 NRS=68.0044 M=1
+ R=2.8 SA=75001.5 SB=75001 A=0.063 P=1.14 MULT=1
MM1035 N_VPWR_M1035_d N_A_2186_367#_M1035_g A_2141_508# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.063 AS=0.0504 PD=0.72 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.8
+ SA=75001.8 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_1804_424#_M1001_d N_SET_B_M1001_g N_VPWR_M1035_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1176 AS=0.063 PD=1.4 PS=0.72 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75002.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1036 N_VPWR_M1036_d N_A_1804_424#_M1036_g N_A_2186_367#_M1036_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1037 N_VPWR_M1037_d N_A_1804_424#_M1037_g N_A_2611_98#_M1037_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.182453 AS=0.28 PD=1.39151 PS=2.56 NRD=11.8003 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1033 N_Q_M1033_d N_A_2611_98#_M1033_g N_VPWR_M1037_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.204347 PD=1.42 PS=1.55849 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75000.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1043 N_Q_M1033_d N_A_2611_98#_M1043_g N_VPWR_M1043_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX46_noxref VNB VPB NWDIODE A=28.3836 P=34.24
c_163 VNB 0 7.29682e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__sdfstp_2.pxi.spice"
*
.ends
*
*
