* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 a_114_74# A3 VGND VNB nshort w=740000u l=150000u
+  ad=4.292e+11p pd=4.12e+06u as=9.093e+11p ps=5.45e+06u
M1001 a_119_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.024e+11p pd=2.78e+06u as=6.608e+11p ps=5.66e+06u
M1002 VPWR B1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=7.728e+11p ps=3.62e+06u
M1003 Y B1 a_114_74# VNB nshort w=740000u l=150000u
+  ad=2.479e+11p pd=2.15e+06u as=0p ps=0u
M1004 Y A3 a_203_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=3.08e+06u
M1005 a_114_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_114_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_203_368# A2 a_119_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
