* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__clkbuf_16 A VGND VNB VPB VPWR X
M1000 X a_114_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=2.688e+12p pd=2.272e+07u as=3.7184e+12p ps=3.128e+07u
M1001 VPWR a_114_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 X a_114_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_114_74# VGND VNB nshort w=420000u l=150000u
+  ad=9.408e+11p pd=1.12e+07u as=1.4826e+12p ps=1.63e+07u
M1004 X a_114_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_114_74# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_114_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_114_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_114_74# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_114_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_114_74# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_114_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_114_74# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_114_74# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_114_74# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_114_74# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_114_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_114_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_114_74# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_114_74# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_114_74# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1021 VPWR A a_114_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A a_114_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1023 VPWR a_114_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_114_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_114_74# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_114_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_114_74# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 X a_114_74# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_114_74# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND A a_114_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND a_114_74# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 X a_114_74# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 X a_114_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR a_114_74# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 X a_114_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_114_74# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_114_74# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR A a_114_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND a_114_74# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
