# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__and4b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.190000 0.595000 1.860000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.550000 2.275000 1.960000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 0.255000 2.810000 0.670000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 1.550000 3.315000 1.880000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.875000 0.480000 4.230000 1.180000 ;
        RECT 3.875000 1.850000 4.230000 2.980000 ;
        RECT 4.060000 1.180000 4.230000 1.850000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.350000 0.405000 0.850000 ;
      RECT 0.115000  0.850000 0.945000 1.020000 ;
      RECT 0.115000  2.030000 0.945000 2.200000 ;
      RECT 0.115000  2.200000 0.445000 2.980000 ;
      RECT 0.575000  0.085000 0.875000 0.680000 ;
      RECT 0.615000  2.370000 0.945000 3.245000 ;
      RECT 0.775000  1.020000 0.945000 1.550000 ;
      RECT 0.775000  1.550000 1.255000 1.880000 ;
      RECT 0.775000  1.880000 0.945000 2.030000 ;
      RECT 1.115000  2.130000 3.095000 2.350000 ;
      RECT 1.115000  2.350000 1.460000 2.460000 ;
      RECT 1.310000  0.600000 1.640000 1.210000 ;
      RECT 1.310000  1.210000 3.705000 1.350000 ;
      RECT 1.310000  1.350000 3.890000 1.380000 ;
      RECT 1.645000  2.535000 2.595000 3.245000 ;
      RECT 2.595000  1.380000 2.765000 2.100000 ;
      RECT 2.595000  2.100000 3.095000 2.130000 ;
      RECT 2.765000  2.350000 3.095000 2.980000 ;
      RECT 3.335000  2.100000 3.665000 3.245000 ;
      RECT 3.375000  0.085000 3.705000 1.040000 ;
      RECT 3.535000  1.380000 3.890000 1.680000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_ls__and4b_1
END LIBRARY
