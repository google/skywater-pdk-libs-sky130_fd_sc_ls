# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__sdfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__sdfxtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.48000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.455000 1.655000 1.785000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.149300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685000 1.800000 12.355000 1.970000 ;
        RECT 10.685000 1.970000 11.015000 2.980000 ;
        RECT 10.745000 0.350000 10.995000 0.880000 ;
        RECT 10.745000 0.880000 12.355000 1.130000 ;
        RECT 11.665000 1.970000 12.355000 2.015000 ;
        RECT 11.665000 2.015000 11.855000 2.980000 ;
        RECT 11.675000 0.350000 11.865000 0.880000 ;
        RECT 11.760000 1.130000 12.355000 1.800000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.435000 1.550000 2.765000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.955000 2.195000 1.285000 ;
        RECT 1.565000 0.810000 2.195000 0.955000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.275000 1.180000 3.685000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.480000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.480000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.480000 0.085000 ;
      RECT  0.000000  3.245000 12.480000 3.415000 ;
      RECT  0.085000  0.350000  0.490000 0.785000 ;
      RECT  0.085000  0.785000  0.255000 1.525000 ;
      RECT  0.085000  1.525000  0.915000 1.955000 ;
      RECT  0.085000  1.955000  2.195000 2.125000 ;
      RECT  0.085000  2.125000  0.555000 2.980000 ;
      RECT  0.660000  0.085000  0.990000 0.785000 ;
      RECT  0.725000  2.300000  1.055000 3.245000 ;
      RECT  1.480000  0.390000  2.535000 0.640000 ;
      RECT  1.595000  2.310000  1.925000 2.390000 ;
      RECT  1.595000  2.390000  4.815000 2.540000 ;
      RECT  1.595000  2.540000  5.405000 2.560000 ;
      RECT  1.595000  2.560000  1.925000 2.980000 ;
      RECT  1.865000  1.470000  2.195000 1.955000 ;
      RECT  1.865000  2.125000  2.195000 2.140000 ;
      RECT  2.365000  0.640000  2.535000 1.180000 ;
      RECT  2.365000  1.180000  3.105000 1.350000 ;
      RECT  2.585000  2.730000  3.205000 3.245000 ;
      RECT  2.705000  0.085000  2.955000 0.810000 ;
      RECT  2.935000  1.350000  3.105000 2.390000 ;
      RECT  3.125000  0.350000  3.455000 0.840000 ;
      RECT  3.125000  0.840000  4.025000 1.010000 ;
      RECT  3.325000  1.820000  4.165000 1.990000 ;
      RECT  3.325000  1.990000  3.655000 2.220000 ;
      RECT  3.685000  0.085000  4.015000 0.670000 ;
      RECT  3.855000  1.010000  4.025000 1.300000 ;
      RECT  3.855000  1.300000  4.165000 1.820000 ;
      RECT  3.885000  2.730000  4.475000 3.245000 ;
      RECT  4.195000  0.255000  5.945000 0.425000 ;
      RECT  4.195000  0.425000  4.445000 1.130000 ;
      RECT  4.335000  1.480000  4.925000 1.650000 ;
      RECT  4.335000  1.650000  4.505000 2.390000 ;
      RECT  4.645000  2.560000  5.405000 2.710000 ;
      RECT  4.675000  0.595000  4.925000 1.480000 ;
      RECT  4.675000  1.820000  4.925000 2.040000 ;
      RECT  4.675000  2.040000  5.405000 2.220000 ;
      RECT  5.075000  2.220000  5.405000 2.370000 ;
      RECT  5.095000  0.425000  5.265000 2.040000 ;
      RECT  5.155000  2.710000  5.405000 2.970000 ;
      RECT  5.435000  0.595000  5.605000 1.610000 ;
      RECT  5.435000  1.610000  7.160000 1.780000 ;
      RECT  5.575000  1.780000  5.745000 2.510000 ;
      RECT  5.575000  2.510000  5.935000 2.970000 ;
      RECT  5.775000  0.425000  5.945000 0.770000 ;
      RECT  5.775000  0.770000  7.160000 0.940000 ;
      RECT  5.775000  0.940000  6.075000 1.360000 ;
      RECT  5.915000  1.950000  6.275000 2.280000 ;
      RECT  6.105000  2.280000  6.275000 2.515000 ;
      RECT  6.105000  2.515000  8.100000 2.685000 ;
      RECT  6.295000  1.110000  7.500000 1.440000 ;
      RECT  6.490000  0.085000  6.820000 0.600000 ;
      RECT  6.680000  2.855000  7.010000 3.245000 ;
      RECT  6.835000  1.780000  7.160000 1.940000 ;
      RECT  6.990000  0.295000  8.125000 0.465000 ;
      RECT  6.990000  0.465000  7.160000 0.770000 ;
      RECT  7.215000  2.175000  7.760000 2.345000 ;
      RECT  7.330000  0.635000  7.785000 0.885000 ;
      RECT  7.330000  0.885000  7.500000 1.110000 ;
      RECT  7.330000  1.440000  7.500000 2.175000 ;
      RECT  7.670000  1.055000  8.125000 1.240000 ;
      RECT  7.670000  1.240000  8.845000 1.410000 ;
      RECT  7.770000  1.625000  8.100000 1.955000 ;
      RECT  7.930000  1.955000  8.100000 2.515000 ;
      RECT  7.955000  0.465000  8.125000 1.055000 ;
      RECT  8.270000  2.020000  9.185000 2.190000 ;
      RECT  8.270000  2.190000  8.600000 2.820000 ;
      RECT  8.295000  0.350000  8.625000 0.900000 ;
      RECT  8.295000  0.900000  9.185000 1.070000 ;
      RECT  8.535000  1.410000  8.845000 1.715000 ;
      RECT  9.015000  1.070000  9.185000 1.470000 ;
      RECT  9.015000  1.470000  9.795000 1.800000 ;
      RECT  9.015000  1.800000  9.185000 2.020000 ;
      RECT  9.195000  0.085000  9.525000 0.730000 ;
      RECT  9.225000  2.360000  9.555000 3.245000 ;
      RECT  9.355000  0.900000  9.665000 1.130000 ;
      RECT  9.355000  1.130000 10.135000 1.300000 ;
      RECT  9.730000  1.970000 10.135000 2.820000 ;
      RECT  9.835000  0.350000 10.005000 1.130000 ;
      RECT  9.965000  1.300000 11.545000 1.630000 ;
      RECT  9.965000  1.630000 10.135000 1.970000 ;
      RECT 10.185000  0.085000 10.515000 0.960000 ;
      RECT 10.305000  1.940000 10.475000 3.245000 ;
      RECT 11.175000  0.085000 11.505000 0.710000 ;
      RECT 11.215000  2.140000 11.465000 3.245000 ;
      RECT 12.035000  0.085000 12.365000 0.710000 ;
      RECT 12.035000  2.185000 12.365000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
  END
END sky130_fd_sc_ls__sdfxtp_4
END LIBRARY
