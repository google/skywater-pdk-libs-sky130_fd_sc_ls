* File: sky130_fd_sc_ls__xor2_4.pex.spice
* Created: Wed Sep  2 11:31:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__XOR2_4%A 1 3 6 8 10 13 15 17 20 22 24 27 31 33 35 36
+ 37 38 40 43 46 50 52 53 55 58 61 62 63 65 66 67 68 69 70 71 76 83 91
c228 63 0 1.24044e-19 $X=3.04 $Y=1.105
c229 55 0 4.48662e-20 $X=0.945 $Y=1.585
c230 36 0 1.17531e-19 $X=6.255 $Y=1.485
c231 22 0 3.52062e-20 $X=5.315 $Y=1.765
c232 15 0 9.55446e-20 $X=4.725 $Y=1.765
c233 6 0 1.34713e-19 $X=0.725 $Y=0.86
r234 88 90 40.1667 $w=3.78e-07 $l=3.15e-07 $layer=POLY_cond $X=5.45 $Y=1.557
+ $X2=5.765 $Y2=1.557
r235 88 89 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.45
+ $Y=1.515 $X2=5.45 $Y2=1.515
r236 86 88 14.664 $w=3.78e-07 $l=1.15e-07 $layer=POLY_cond $X=5.335 $Y=1.557
+ $X2=5.45 $Y2=1.557
r237 85 86 2.55026 $w=3.78e-07 $l=2e-08 $layer=POLY_cond $X=5.315 $Y=1.557
+ $X2=5.335 $Y2=1.557
r238 80 81 22.7358 $w=3.71e-07 $l=1.75e-07 $layer=POLY_cond $X=0.55 $Y=1.652
+ $X2=0.725 $Y2=1.652
r239 79 89 9.21954 $w=4.23e-07 $l=3.4e-07 $layer=LI1_cond $X=5.11 $Y=1.562
+ $X2=5.45 $Y2=1.562
r240 78 79 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.11
+ $Y=1.515 $X2=5.11 $Y2=1.515
r241 76 85 12.3802 $w=3.78e-07 $l=1.08995e-07 $layer=POLY_cond $X=5.225 $Y=1.515
+ $X2=5.315 $Y2=1.557
r242 76 78 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=5.225 $Y=1.515
+ $X2=5.11 $Y2=1.515
r243 71 89 1.89814 $w=4.23e-07 $l=7e-08 $layer=LI1_cond $X=5.52 $Y=1.562
+ $X2=5.45 $Y2=1.562
r244 70 79 1.89814 $w=4.23e-07 $l=7e-08 $layer=LI1_cond $X=5.04 $Y=1.562
+ $X2=5.11 $Y2=1.562
r245 69 70 13.0158 $w=4.23e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.562
+ $X2=5.04 $Y2=1.562
r246 69 91 4.60977 $w=4.23e-07 $l=1.7e-07 $layer=LI1_cond $X=4.56 $Y=1.562
+ $X2=4.39 $Y2=1.562
r247 68 91 9.38859 $w=4.25e-07 $l=3.1e-07 $layer=LI1_cond $X=4.08 $Y=1.562
+ $X2=4.39 $Y2=1.562
r248 66 67 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=1.275 $Y=0.675
+ $X2=1.445 $Y2=0.675
r249 65 68 8.18076 $w=3.43e-07 $l=3.18842e-07 $layer=LI1_cond $X=3.85 $Y=1.35
+ $X2=4.08 $Y2=1.562
r250 64 65 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.85 $Y=1.19
+ $X2=3.85 $Y2=1.35
r251 62 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=1.105
+ $X2=3.85 $Y2=1.19
r252 62 63 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.765 $Y=1.105
+ $X2=3.04 $Y2=1.105
r253 61 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.955 $Y=1.02
+ $X2=3.04 $Y2=1.105
r254 60 61 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.955 $Y=0.77
+ $X2=2.955 $Y2=1.02
r255 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.87 $Y=0.685
+ $X2=2.955 $Y2=0.77
r256 58 67 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=2.87 $Y=0.685
+ $X2=1.445 $Y2=0.685
r257 56 83 13.6415 $w=3.71e-07 $l=1.05e-07 $layer=POLY_cond $X=0.945 $Y=1.652
+ $X2=1.05 $Y2=1.652
r258 56 81 28.5822 $w=3.71e-07 $l=2.2e-07 $layer=POLY_cond $X=0.945 $Y=1.652
+ $X2=0.725 $Y2=1.652
r259 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.945
+ $Y=1.585 $X2=0.945 $Y2=1.585
r260 53 55 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=0.685 $Y=1.585
+ $X2=0.945 $Y2=1.585
r261 52 66 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.685 $Y=0.665
+ $X2=1.275 $Y2=0.665
r262 50 53 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.6 $Y=1.42
+ $X2=0.685 $Y2=1.585
r263 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.6 $Y=0.75
+ $X2=0.685 $Y2=0.665
r264 49 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.6 $Y=0.75 $X2=0.6
+ $Y2=1.42
r265 45 78 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=4.82 $Y=1.515
+ $X2=5.11 $Y2=1.515
r266 45 46 5.03009 $w=3.3e-07 $l=2.85832e-07 $layer=POLY_cond $X=4.82 $Y=1.515
+ $X2=4.605 $Y2=1.35
r267 43 48 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.355 $Y=0.74
+ $X2=6.355 $Y2=1.35
r268 38 40 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.345 $Y=1.765
+ $X2=6.345 $Y2=2.4
r269 37 90 15.4823 $w=3.78e-07 $l=1.20748e-07 $layer=POLY_cond $X=5.855 $Y=1.485
+ $X2=5.765 $Y2=1.557
r270 36 38 110.989 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=6.345 $Y=1.485
+ $X2=6.345 $Y2=1.765
r271 36 48 54.6256 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=6.345 $Y=1.485
+ $X2=6.345 $Y2=1.35
r272 36 37 88.8695 $w=2.7e-07 $l=4e-07 $layer=POLY_cond $X=6.255 $Y=1.485
+ $X2=5.855 $Y2=1.485
r273 33 90 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.765 $Y=1.765
+ $X2=5.765 $Y2=1.557
r274 33 35 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.765 $Y=1.765
+ $X2=5.765 $Y2=2.4
r275 29 90 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.765 $Y=1.35
+ $X2=5.765 $Y2=1.557
r276 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.765 $Y=1.35
+ $X2=5.765 $Y2=0.74
r277 25 86 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.335 $Y=1.35
+ $X2=5.335 $Y2=1.557
r278 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.335 $Y=1.35
+ $X2=5.335 $Y2=0.74
r279 22 85 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.315 $Y=1.765
+ $X2=5.315 $Y2=1.557
r280 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.315 $Y=1.765
+ $X2=5.315 $Y2=2.4
r281 18 46 37.0704 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=4.745 $Y=1.35
+ $X2=4.605 $Y2=1.35
r282 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.745 $Y=1.35
+ $X2=4.745 $Y2=0.74
r283 15 46 37.0704 $w=1.5e-07 $l=4.71195e-07 $layer=POLY_cond $X=4.725 $Y=1.765
+ $X2=4.605 $Y2=1.35
r284 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.725 $Y=1.765
+ $X2=4.725 $Y2=2.4
r285 11 83 13.6415 $w=3.71e-07 $l=2.79614e-07 $layer=POLY_cond $X=1.155 $Y=1.42
+ $X2=1.05 $Y2=1.652
r286 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.155 $Y=1.42
+ $X2=1.155 $Y2=0.86
r287 8 83 24.032 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.05 $Y=1.885
+ $X2=1.05 $Y2=1.652
r288 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.05 $Y=1.885
+ $X2=1.05 $Y2=2.46
r289 4 81 24.032 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.725 $Y=1.42
+ $X2=0.725 $Y2=1.652
r290 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.725 $Y=1.42
+ $X2=0.725 $Y2=0.86
r291 1 80 24.032 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.55 $Y=1.885
+ $X2=0.55 $Y2=1.652
r292 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.55 $Y=1.885
+ $X2=0.55 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_4%B 1 3 6 8 10 13 15 16 20 21 23 24 25 29 30 32
+ 33 35 38 40 42 44 46 50 51 53 54 55 57 58 59 63 64 65 66 67 88 92
c205 57 0 3.52062e-20 $X=5.89 $Y=1.78
c206 15 0 1.53262e-19 $X=6.795 $Y=1.275
c207 13 0 1.24044e-19 $X=2.285 $Y=0.86
c208 6 0 1.87977e-19 $X=1.745 $Y=0.86
r209 90 92 0.670025 $w=4.28e-07 $l=2.5e-08 $layer=LI1_cond $X=5.975 $Y=1.565
+ $X2=6 $Y2=1.565
r210 87 88 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8
+ $Y=1.515 $X2=8 $Y2=1.515
r211 82 84 46.1097 $w=3.92e-07 $l=3.75e-07 $layer=POLY_cond $X=7.32 $Y=1.475
+ $X2=7.695 $Y2=1.475
r212 82 83 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.32
+ $Y=1.515 $X2=7.32 $Y2=1.515
r213 80 82 9.22194 $w=3.92e-07 $l=7.5e-08 $layer=POLY_cond $X=7.245 $Y=1.475
+ $X2=7.32 $Y2=1.475
r214 79 80 3.68878 $w=3.92e-07 $l=3e-08 $layer=POLY_cond $X=7.215 $Y=1.475
+ $X2=7.245 $Y2=1.475
r215 75 76 26.8505 $w=3.68e-07 $l=2.05e-07 $layer=POLY_cond $X=1.745 $Y=1.677
+ $X2=1.95 $Y2=1.677
r216 74 75 32.0897 $w=3.68e-07 $l=2.45e-07 $layer=POLY_cond $X=1.5 $Y=1.677
+ $X2=1.745 $Y2=1.677
r217 67 88 2.14408 $w=4.28e-07 $l=8e-08 $layer=LI1_cond $X=7.92 $Y=1.565 $X2=8
+ $Y2=1.565
r218 66 67 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.92 $Y2=1.565
r219 66 83 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.32 $Y2=1.565
r220 65 83 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.32 $Y2=1.565
r221 64 65 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.96 $Y2=1.565
r222 63 90 2.44569 $w=4.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.89 $Y=1.565
+ $X2=5.975 $Y2=1.565
r223 63 64 12.0604 $w=4.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.03 $Y=1.565
+ $X2=6.48 $Y2=1.565
r224 63 92 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=6.03 $Y=1.565 $X2=6
+ $Y2=1.565
r225 59 61 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.57 $Y=1.935
+ $X2=3.57 $Y2=2.03
r226 57 63 6.18617 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=5.89 $Y=1.78
+ $X2=5.89 $Y2=1.565
r227 57 58 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.89 $Y=1.78
+ $X2=5.89 $Y2=1.945
r228 56 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=2.03
+ $X2=3.57 $Y2=2.03
r229 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.805 $Y=2.03
+ $X2=5.89 $Y2=1.945
r230 55 56 140.267 $w=1.68e-07 $l=2.15e-06 $layer=LI1_cond $X=5.805 $Y=2.03
+ $X2=3.655 $Y2=2.03
r231 53 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.485 $Y=1.935
+ $X2=3.57 $Y2=1.935
r232 53 54 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=3.485 $Y=1.935
+ $X2=2.36 $Y2=1.935
r233 51 78 11.788 $w=3.68e-07 $l=9e-08 $layer=POLY_cond $X=2.195 $Y=1.677
+ $X2=2.285 $Y2=1.677
r234 51 76 32.0897 $w=3.68e-07 $l=2.45e-07 $layer=POLY_cond $X=2.195 $Y=1.677
+ $X2=1.95 $Y2=1.677
r235 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.195
+ $Y=1.635 $X2=2.195 $Y2=1.635
r236 48 54 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.195 $Y=1.85
+ $X2=2.36 $Y2=1.935
r237 48 50 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.195 $Y=1.85
+ $X2=2.195 $Y2=1.635
r238 44 46 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.145 $Y=1.765
+ $X2=8.145 $Y2=2.4
r239 40 44 25.3688 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.145 $Y=1.475
+ $X2=8.145 $Y2=1.765
r240 40 87 17.8291 $w=3.92e-07 $l=1.45e-07 $layer=POLY_cond $X=8.145 $Y=1.475
+ $X2=8 $Y2=1.475
r241 40 42 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.145 $Y=1.35
+ $X2=8.145 $Y2=0.74
r242 36 87 35.0434 $w=3.92e-07 $l=2.85e-07 $layer=POLY_cond $X=7.715 $Y=1.475
+ $X2=8 $Y2=1.475
r243 36 84 2.45918 $w=3.92e-07 $l=2e-08 $layer=POLY_cond $X=7.715 $Y=1.475
+ $X2=7.695 $Y2=1.475
r244 36 38 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.715 $Y=1.35
+ $X2=7.715 $Y2=0.74
r245 33 84 25.3688 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.695 $Y=1.765
+ $X2=7.695 $Y2=1.475
r246 33 35 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.695 $Y=1.765
+ $X2=7.695 $Y2=2.4
r247 30 80 25.3688 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.245 $Y=1.765
+ $X2=7.245 $Y2=1.475
r248 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.245 $Y=1.765
+ $X2=7.245 $Y2=2.4
r249 27 79 25.3688 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.215 $Y=1.185
+ $X2=7.215 $Y2=1.475
r250 27 29 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.215 $Y=1.185
+ $X2=7.215 $Y2=0.74
r251 26 29 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.215 $Y=0.295
+ $X2=7.215 $Y2=0.74
r252 24 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.14 $Y=0.22
+ $X2=7.215 $Y2=0.295
r253 24 25 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=7.14 $Y=0.22
+ $X2=6.86 $Y2=0.22
r254 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.795 $Y=1.765
+ $X2=6.795 $Y2=2.4
r255 20 47 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.785 $Y=0.74
+ $X2=6.785 $Y2=1.185
r256 17 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.785 $Y=0.295
+ $X2=6.86 $Y2=0.22
r257 17 20 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.785 $Y=0.295
+ $X2=6.785 $Y2=0.74
r258 16 21 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.795 $Y=1.675
+ $X2=6.795 $Y2=1.765
r259 15 47 36.5962 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.795 $Y=1.275
+ $X2=6.795 $Y2=1.185
r260 15 16 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=6.795 $Y=1.275
+ $X2=6.795 $Y2=1.675
r261 11 78 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.285 $Y=1.47
+ $X2=2.285 $Y2=1.677
r262 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.285 $Y=1.47
+ $X2=2.285 $Y2=0.86
r263 8 76 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.95 $Y=1.885
+ $X2=1.95 $Y2=1.677
r264 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.95 $Y=1.885
+ $X2=1.95 $Y2=2.46
r265 4 75 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.745 $Y=1.47
+ $X2=1.745 $Y2=1.677
r266 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.745 $Y=1.47
+ $X2=1.745 $Y2=0.86
r267 1 74 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.5 $Y=1.885
+ $X2=1.5 $Y2=1.677
r268 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.5 $Y=1.885 $X2=1.5
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_4%A_160_98# 1 2 3 10 12 13 15 16 18 19 21 22 24
+ 25 26 27 29 30 32 36 38 43 44 49 55 56
c140 55 0 2.77823e-19 $X=1.105 $Y=1.085
r141 62 63 34.3242 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=3.59 $Y=1.557
+ $X2=3.825 $Y2=1.557
r142 59 60 65.7273 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=2.925 $Y=1.557
+ $X2=3.375 $Y2=1.557
r143 58 59 7.30303 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=2.875 $Y=1.557
+ $X2=2.925 $Y2=1.557
r144 53 55 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.94 $Y=1.085
+ $X2=1.105 $Y2=1.085
r145 50 62 23.3697 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.43 $Y=1.557
+ $X2=3.59 $Y2=1.557
r146 50 60 8.03333 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.43 $Y=1.557
+ $X2=3.375 $Y2=1.557
r147 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.515 $X2=3.43 $Y2=1.515
r148 47 58 18.2576 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.75 $Y=1.557
+ $X2=2.875 $Y2=1.557
r149 46 49 24.4894 $w=3.18e-07 $l=6.8e-07 $layer=LI1_cond $X=2.75 $Y=1.52
+ $X2=3.43 $Y2=1.52
r150 46 47 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.75
+ $Y=1.515 $X2=2.75 $Y2=1.515
r151 44 46 1.80069 $w=3.18e-07 $l=5e-08 $layer=LI1_cond $X=2.7 $Y=1.52 $X2=2.75
+ $Y2=1.52
r152 43 44 7.68211 $w=3.2e-07 $l=1.9799e-07 $layer=LI1_cond $X=2.615 $Y=1.36
+ $X2=2.7 $Y2=1.52
r153 42 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.615 $Y=1.19
+ $X2=2.615 $Y2=1.36
r154 39 56 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.81 $Y=1.065
+ $X2=1.685 $Y2=1.065
r155 39 41 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=1.81 $Y=1.065
+ $X2=2.015 $Y2=1.065
r156 38 42 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.53 $Y=1.065
+ $X2=2.615 $Y2=1.19
r157 38 41 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=2.53 $Y=1.065
+ $X2=2.015 $Y2=1.065
r158 34 56 1.34256 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.685 $Y=1.19
+ $X2=1.685 $Y2=1.065
r159 34 36 42.1794 $w=2.48e-07 $l=9.15e-07 $layer=LI1_cond $X=1.685 $Y=1.19
+ $X2=1.685 $Y2=2.105
r160 32 56 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.56 $Y=1.065
+ $X2=1.685 $Y2=1.065
r161 32 55 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=1.56 $Y=1.065
+ $X2=1.105 $Y2=1.065
r162 27 30 64.3434 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=4.275 $Y=1.765
+ $X2=4.275 $Y2=1.605
r163 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.275 $Y=1.765
+ $X2=4.275 $Y2=2.4
r164 26 63 27.6456 $w=3.3e-07 $l=1.11445e-07 $layer=POLY_cond $X=3.915 $Y=1.605
+ $X2=3.825 $Y2=1.557
r165 25 30 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.185 $Y=1.605
+ $X2=4.275 $Y2=1.605
r166 25 26 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.185 $Y=1.605
+ $X2=3.915 $Y2=1.605
r167 22 63 21.2229 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.825 $Y=1.765
+ $X2=3.825 $Y2=1.557
r168 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.825 $Y=1.765
+ $X2=3.825 $Y2=2.4
r169 19 62 21.2229 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.59 $Y=1.35
+ $X2=3.59 $Y2=1.557
r170 19 21 157.453 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.59 $Y=1.35
+ $X2=3.59 $Y2=0.86
r171 16 60 21.2229 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.375 $Y=1.765
+ $X2=3.375 $Y2=1.557
r172 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.375 $Y=1.765
+ $X2=3.375 $Y2=2.4
r173 13 59 21.2229 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.925 $Y=1.765
+ $X2=2.925 $Y2=1.557
r174 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.925 $Y=1.765
+ $X2=2.925 $Y2=2.4
r175 10 58 21.2229 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.875 $Y=1.35
+ $X2=2.875 $Y2=1.557
r176 10 12 157.453 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=2.875 $Y=1.35
+ $X2=2.875 $Y2=0.86
r177 3 36 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.575
+ $Y=1.96 $X2=1.725 $Y2=2.105
r178 2 41 182 $w=1.7e-07 $l=6.2494e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.49 $X2=2.015 $Y2=1.025
r179 1 53 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=0.8
+ $Y=0.49 $X2=0.94 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_4%A_36_392# 1 2 3 12 16 17 21 24 25 28
r46 26 28 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=2.175 $Y=2.905
+ $X2=2.175 $Y2=2.355
r47 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.01 $Y=2.99
+ $X2=2.175 $Y2=2.905
r48 24 25 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.01 $Y=2.99
+ $X2=1.36 $Y2=2.99
r49 21 23 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=1.235 $Y=2.105
+ $X2=1.235 $Y2=2.815
r50 19 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.235 $Y=2.905
+ $X2=1.36 $Y2=2.99
r51 19 23 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.235 $Y=2.905
+ $X2=1.235 $Y2=2.815
r52 18 21 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=1.235 $Y=2.09
+ $X2=1.235 $Y2=2.105
r53 16 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.11 $Y=2.005
+ $X2=1.235 $Y2=2.09
r54 16 17 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.11 $Y=2.005
+ $X2=0.49 $Y2=2.005
r55 12 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.325 $Y=2.105
+ $X2=0.325 $Y2=2.815
r56 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.325 $Y=2.09
+ $X2=0.49 $Y2=2.005
r57 10 12 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.325 $Y=2.09
+ $X2=0.325 $Y2=2.105
r58 3 28 300 $w=1.7e-07 $l=4.63977e-07 $layer=licon1_PDIFF $count=2 $X=2.025
+ $Y=1.96 $X2=2.175 $Y2=2.355
r59 2 23 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.96 $X2=1.275 $Y2=2.815
r60 2 21 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.96 $X2=1.275 $Y2=2.105
r61 1 14 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=1.96 $X2=0.325 $Y2=2.815
r62 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=1.96 $X2=0.325 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_4%VPWR 1 2 3 4 5 20 24 28 30 32 40 45 50 57 58
+ 61 64 71 78 81
r117 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r118 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r119 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r120 71 74 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.055 $Y=3.05
+ $X2=6.055 $Y2=3.33
r121 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r122 64 67 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=5.02 $Y=3.05
+ $X2=5.02 $Y2=3.33
r123 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r124 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r125 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r126 55 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.005 $Y=3.33
+ $X2=7.92 $Y2=3.33
r127 55 57 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.005 $Y=3.33
+ $X2=8.4 $Y2=3.33
r128 54 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r129 54 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r130 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r131 51 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.105 $Y=3.33
+ $X2=6.98 $Y2=3.33
r132 51 53 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.105 $Y=3.33
+ $X2=7.44 $Y2=3.33
r133 50 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.92 $Y2=3.33
r134 50 53 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.44 $Y2=3.33
r135 49 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r136 49 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r137 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r138 46 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.22 $Y=3.33
+ $X2=6.055 $Y2=3.33
r139 46 48 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.22 $Y=3.33
+ $X2=6.48 $Y2=3.33
r140 45 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.855 $Y=3.33
+ $X2=6.98 $Y2=3.33
r141 45 48 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.855 $Y=3.33
+ $X2=6.48 $Y2=3.33
r142 44 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r143 44 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r144 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r145 41 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.185 $Y=3.33
+ $X2=5.02 $Y2=3.33
r146 41 43 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.185 $Y=3.33
+ $X2=5.52 $Y2=3.33
r147 40 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.89 $Y=3.33
+ $X2=6.055 $Y2=3.33
r148 40 43 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.89 $Y=3.33
+ $X2=5.52 $Y2=3.33
r149 39 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r150 38 39 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r151 36 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r152 35 38 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r153 35 36 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r154 33 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.94 $Y=3.33
+ $X2=0.815 $Y2=3.33
r155 33 35 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.94 $Y=3.33
+ $X2=1.2 $Y2=3.33
r156 32 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=5.02 $Y2=3.33
r157 32 38 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=4.56 $Y2=3.33
r158 30 39 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r159 30 36 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=1.2 $Y2=3.33
r160 26 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=3.33
r161 26 28 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=2.805
r162 22 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.98 $Y=3.245
+ $X2=6.98 $Y2=3.33
r163 22 24 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=6.98 $Y=3.245
+ $X2=6.98 $Y2=2.805
r164 18 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r165 18 20 37.8001 $w=2.48e-07 $l=8.2e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.425
r166 5 28 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=7.77
+ $Y=1.84 $X2=7.92 $Y2=2.805
r167 4 24 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=6.87
+ $Y=1.84 $X2=7.02 $Y2=2.805
r168 3 71 600 $w=1.7e-07 $l=1.31311e-06 $layer=licon1_PDIFF $count=1 $X=5.84
+ $Y=1.84 $X2=6.055 $Y2=3.05
r169 2 64 600 $w=1.7e-07 $l=1.31541e-06 $layer=licon1_PDIFF $count=1 $X=4.8
+ $Y=1.84 $X2=5.02 $Y2=3.05
r170 1 20 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=0.625
+ $Y=1.96 $X2=0.775 $Y2=2.425
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_4%A_514_368# 1 2 3 4 5 6 7 24 26 27 30 32 36 38
+ 39 40 44 48 49 57 58 64 66
c117 32 0 9.55446e-20 $X=4.415 $Y=2.99
r118 56 58 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=5.54 $Y=2.802
+ $X2=5.705 $Y2=2.802
r119 56 57 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=5.54 $Y=2.802
+ $X2=5.375 $Y2=2.802
r120 52 53 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=4.54 $Y=2.8
+ $X2=4.54 $Y2=2.99
r121 49 52 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.54 $Y=2.71 $X2=4.54
+ $Y2=2.8
r122 45 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.635 $Y=2.375
+ $X2=7.47 $Y2=2.375
r123 44 66 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.205 $Y=2.375
+ $X2=8.37 $Y2=2.375
r124 44 45 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.205 $Y=2.375
+ $X2=7.635 $Y2=2.375
r125 41 60 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.655 $Y=2.375
+ $X2=6.57 $Y2=2.375
r126 40 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=2.375
+ $X2=7.47 $Y2=2.375
r127 40 41 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=7.305 $Y=2.375
+ $X2=6.655 $Y2=2.375
r128 39 62 3.40825 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=6.57 $Y=2.625
+ $X2=6.57 $Y2=2.802
r129 38 60 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.57 $Y=2.46
+ $X2=6.57 $Y2=2.375
r130 38 39 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.57 $Y=2.46
+ $X2=6.57 $Y2=2.625
r131 36 62 3.40825 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=6.485 $Y=2.71
+ $X2=6.57 $Y2=2.802
r132 36 58 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.485 $Y=2.71
+ $X2=5.705 $Y2=2.71
r133 35 49 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.665 $Y=2.71
+ $X2=4.54 $Y2=2.71
r134 35 57 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.665 $Y=2.71
+ $X2=5.375 $Y2=2.71
r135 33 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=2.99
+ $X2=3.6 $Y2=2.99
r136 32 53 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.415 $Y=2.99
+ $X2=4.54 $Y2=2.99
r137 32 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.415 $Y=2.99
+ $X2=3.685 $Y2=2.99
r138 28 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=2.905 $X2=3.6
+ $Y2=2.99
r139 28 30 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.6 $Y=2.905
+ $X2=3.6 $Y2=2.8
r140 26 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=2.99
+ $X2=3.6 $Y2=2.99
r141 26 27 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.515 $Y=2.99
+ $X2=2.785 $Y2=2.99
r142 22 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.66 $Y=2.905
+ $X2=2.785 $Y2=2.99
r143 22 24 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=2.66 $Y=2.905
+ $X2=2.66 $Y2=2.355
r144 7 66 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=8.22
+ $Y=1.84 $X2=8.37 $Y2=2.455
r145 6 64 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=7.32
+ $Y=1.84 $X2=7.47 $Y2=2.455
r146 5 62 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.42
+ $Y=1.84 $X2=6.57 $Y2=2.815
r147 5 60 600 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=1 $X=6.42
+ $Y=1.84 $X2=6.57 $Y2=2.455
r148 4 56 600 $w=1.7e-07 $l=1.03228e-06 $layer=licon1_PDIFF $count=1 $X=5.39
+ $Y=1.84 $X2=5.54 $Y2=2.8
r149 3 52 600 $w=1.7e-07 $l=1.03228e-06 $layer=licon1_PDIFF $count=1 $X=4.35
+ $Y=1.84 $X2=4.5 $Y2=2.8
r150 2 30 600 $w=1.7e-07 $l=1.03228e-06 $layer=licon1_PDIFF $count=1 $X=3.45
+ $Y=1.84 $X2=3.6 $Y2=2.8
r151 1 24 300 $w=1.7e-07 $l=5.76346e-07 $layer=licon1_PDIFF $count=2 $X=2.57
+ $Y=1.84 $X2=2.7 $Y2=2.355
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_4%X 1 2 3 4 5 18 21 22 24 25 27 28 29 32 34 38
+ 40 43 45 50 54 55 56 60 63
c172 24 0 2.70793e-19 $X=6.835 $Y=1.095
r173 59 60 9.22412 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=2.51
+ $X2=3.885 $Y2=2.51
r174 56 63 8.42674 $w=4.48e-07 $l=1.35e-07 $layer=LI1_cond $X=4.08 $Y=2.51
+ $X2=4.215 $Y2=2.51
r175 56 59 0.797386 $w=4.48e-07 $l=3e-08 $layer=LI1_cond $X=4.08 $Y=2.51
+ $X2=4.05 $Y2=2.51
r176 50 52 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.375 $Y=0.66
+ $X2=3.375 $Y2=0.765
r177 45 47 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.15 $Y=2.275
+ $X2=3.15 $Y2=2.37
r178 42 43 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=8.42 $Y=1.18
+ $X2=8.42 $Y2=1.95
r179 41 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.015 $Y=1.095
+ $X2=7.93 $Y2=1.095
r180 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.335 $Y=1.095
+ $X2=8.42 $Y2=1.18
r181 40 41 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.335 $Y=1.095
+ $X2=8.015 $Y2=1.095
r182 36 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=1.01
+ $X2=7.93 $Y2=1.095
r183 36 38 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.93 $Y=1.01
+ $X2=7.93 $Y2=0.805
r184 35 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.165 $Y=1.095
+ $X2=7 $Y2=1.095
r185 34 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.845 $Y=1.095
+ $X2=7.93 $Y2=1.095
r186 34 35 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.845 $Y=1.095
+ $X2=7.165 $Y2=1.095
r187 30 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=1.01 $X2=7
+ $Y2=1.095
r188 30 32 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=7 $Y=1.01 $X2=7
+ $Y2=0.76
r189 28 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.335 $Y=2.035
+ $X2=8.42 $Y2=1.95
r190 28 29 131.786 $w=1.68e-07 $l=2.02e-06 $layer=LI1_cond $X=8.335 $Y=2.035
+ $X2=6.315 $Y2=2.035
r191 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.23 $Y=2.12
+ $X2=6.315 $Y2=2.035
r192 26 27 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.23 $Y=2.12
+ $X2=6.23 $Y2=2.285
r193 24 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.835 $Y=1.095
+ $X2=7 $Y2=1.095
r194 24 25 167.016 $w=1.68e-07 $l=2.56e-06 $layer=LI1_cond $X=6.835 $Y=1.095
+ $X2=4.275 $Y2=1.095
r195 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.145 $Y=2.37
+ $X2=6.23 $Y2=2.285
r196 22 63 125.914 $w=1.68e-07 $l=1.93e-06 $layer=LI1_cond $X=6.145 $Y=2.37
+ $X2=4.215 $Y2=2.37
r197 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.19 $Y=1.01
+ $X2=4.275 $Y2=1.095
r198 20 21 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.19 $Y=0.85
+ $X2=4.19 $Y2=1.01
r199 19 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.54 $Y=0.765
+ $X2=3.375 $Y2=0.765
r200 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.105 $Y=0.765
+ $X2=4.19 $Y2=0.85
r201 18 19 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.105 $Y=0.765
+ $X2=3.54 $Y2=0.765
r202 17 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.315 $Y=2.37
+ $X2=3.15 $Y2=2.37
r203 17 60 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.315 $Y=2.37
+ $X2=3.885 $Y2=2.37
r204 5 59 600 $w=1.7e-07 $l=7.41215e-07 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=1.84 $X2=4.05 $Y2=2.51
r205 4 45 300 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_PDIFF $count=2 $X=3
+ $Y=1.84 $X2=3.15 $Y2=2.275
r206 3 38 182 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_NDIFF $count=1 $X=7.79
+ $Y=0.37 $X2=7.93 $Y2=0.805
r207 2 32 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=6.86
+ $Y=0.37 $X2=7 $Y2=0.76
r208 1 50 182 $w=1.7e-07 $l=5.02867e-07 $layer=licon1_NDIFF $count=1 $X=2.95
+ $Y=0.49 $X2=3.375 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_4%VGND 1 2 3 4 5 6 19 21 25 29 33 37 39 40 47
+ 48 49 55 63 67 77 78 84 87 90
r122 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r123 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r124 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r125 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r126 77 78 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r127 75 78 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r128 75 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r129 74 77 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r130 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r131 72 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.225 $Y=0 $X2=6.06
+ $Y2=0
r132 72 74 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.225 $Y=0
+ $X2=6.48 $Y2=0
r133 71 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r134 71 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r135 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r136 68 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.205 $Y=0 $X2=5.04
+ $Y2=0
r137 68 70 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.205 $Y=0
+ $X2=5.52 $Y2=0
r138 67 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.895 $Y=0 $X2=6.06
+ $Y2=0
r139 67 70 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.895 $Y=0
+ $X2=5.52 $Y2=0
r140 66 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r141 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r142 63 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=0 $X2=5.04
+ $Y2=0
r143 63 65 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.875 $Y=0
+ $X2=4.56 $Y2=0
r144 62 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r145 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r146 59 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.58
+ $Y2=0
r147 59 61 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=3.6
+ $Y2=0
r148 58 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r149 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r150 55 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.58
+ $Y2=0
r151 55 57 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.415 $Y=0
+ $X2=2.16 $Y2=0
r152 54 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r153 54 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r154 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r155 51 81 4.03846 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r156 51 53 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=1.2
+ $Y2=0
r157 49 66 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r158 49 62 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=0 $X2=3.6
+ $Y2=0
r159 47 61 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.6
+ $Y2=0
r160 47 48 10.0494 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.927
+ $Y2=0
r161 46 65 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=4.135 $Y=0
+ $X2=4.56 $Y2=0
r162 46 48 10.0494 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=4.135 $Y=0
+ $X2=3.927 $Y2=0
r163 42 57 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=1.615 $Y=0
+ $X2=2.16 $Y2=0
r164 40 53 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.2
+ $Y2=0
r165 39 44 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.45
+ $Y2=0.325
r166 39 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.615
+ $Y2=0
r167 39 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.285
+ $Y2=0
r168 35 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.06 $Y=0.085
+ $X2=6.06 $Y2=0
r169 35 37 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6.06 $Y=0.085
+ $X2=6.06 $Y2=0.335
r170 31 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=0.085
+ $X2=5.04 $Y2=0
r171 31 33 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=5.04 $Y=0.085
+ $X2=5.04 $Y2=0.335
r172 27 48 1.57254 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.927 $Y=0.085
+ $X2=3.927 $Y2=0
r173 27 29 7.22012 $w=4.13e-07 $l=2.6e-07 $layer=LI1_cond $X=3.927 $Y=0.085
+ $X2=3.927 $Y2=0.345
r174 23 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=0.085
+ $X2=2.58 $Y2=0
r175 23 25 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.58 $Y=0.085
+ $X2=2.58 $Y2=0.335
r176 19 81 3.10471 $w=2.5e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.22 $Y=0.085
+ $X2=0.172 $Y2=0
r177 19 21 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=0.22 $Y=0.085
+ $X2=0.22 $Y2=0.635
r178 6 37 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=5.84
+ $Y=0.37 $X2=6.06 $Y2=0.335
r179 5 33 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=4.82
+ $Y=0.37 $X2=5.04 $Y2=0.335
r180 4 29 182 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=1 $X=3.665
+ $Y=0.49 $X2=3.925 $Y2=0.345
r181 3 25 182 $w=1.7e-07 $l=2.87228e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.49 $X2=2.58 $Y2=0.335
r182 2 44 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=1.23
+ $Y=0.49 $X2=1.45 $Y2=0.325
r183 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.49 $X2=0.26 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_4%A_877_74# 1 2 3 4 5 20 23 24 25 28 30 34 37
+ 40 41 44
r77 39 41 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.55 $Y=0.595
+ $X2=5.715 $Y2=0.595
r78 39 40 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.55 $Y=0.595
+ $X2=5.385 $Y2=0.595
r79 32 34 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=8.36 $Y=0.425
+ $X2=8.36 $Y2=0.675
r80 31 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.665 $Y=0.34
+ $X2=7.5 $Y2=0.34
r81 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.195 $Y=0.34
+ $X2=8.36 $Y2=0.425
r82 30 31 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.195 $Y=0.34
+ $X2=7.665 $Y2=0.34
r83 26 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=0.425 $X2=7.5
+ $Y2=0.34
r84 26 28 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=7.5 $Y=0.425 $X2=7.5
+ $Y2=0.675
r85 24 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.335 $Y=0.34
+ $X2=7.5 $Y2=0.34
r86 24 25 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.335 $Y=0.34
+ $X2=6.655 $Y2=0.34
r87 23 43 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.53 $Y=0.67 $X2=6.53
+ $Y2=0.755
r88 22 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.53 $Y=0.425
+ $X2=6.655 $Y2=0.34
r89 22 23 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=6.53 $Y=0.425
+ $X2=6.53 $Y2=0.67
r90 20 43 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.405 $Y=0.755
+ $X2=6.53 $Y2=0.755
r91 20 41 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.405 $Y=0.755
+ $X2=5.715 $Y2=0.755
r92 19 37 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.695 $Y=0.755
+ $X2=4.57 $Y2=0.755
r93 19 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.695 $Y=0.755
+ $X2=5.385 $Y2=0.755
r94 5 34 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.37 $X2=8.36 $Y2=0.675
r95 4 28 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=7.29
+ $Y=0.37 $X2=7.5 $Y2=0.675
r96 3 43 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=6.43
+ $Y=0.37 $X2=6.57 $Y2=0.675
r97 2 39 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=5.41
+ $Y=0.37 $X2=5.55 $Y2=0.675
r98 1 37 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.37 $X2=4.53 $Y2=0.675
.ends

