* File: sky130_fd_sc_ls__dfrbp_1.pxi.spice
* Created: Wed Sep  2 11:00:45 2020
* 
x_PM_SKY130_FD_SC_LS__DFRBP_1%D N_D_c_247_n N_D_M1021_g N_D_M1007_g N_D_c_248_n
+ D D D N_D_c_244_n N_D_c_245_n N_D_c_246_n PM_SKY130_FD_SC_LS__DFRBP_1%D
x_PM_SKY130_FD_SC_LS__DFRBP_1%CLK N_CLK_M1000_g N_CLK_M1001_g CLK N_CLK_c_278_n
+ N_CLK_c_279_n PM_SKY130_FD_SC_LS__DFRBP_1%CLK
x_PM_SKY130_FD_SC_LS__DFRBP_1%A_500_392# N_A_500_392#_M1029_d
+ N_A_500_392#_M1030_d N_A_500_392#_c_325_n N_A_500_392#_c_345_n
+ N_A_500_392#_M1023_g N_A_500_392#_c_326_n N_A_500_392#_c_327_n
+ N_A_500_392#_M1010_g N_A_500_392#_c_328_n N_A_500_392#_M1004_g
+ N_A_500_392#_c_329_n N_A_500_392#_c_330_n N_A_500_392#_c_347_n
+ N_A_500_392#_M1018_g N_A_500_392#_c_348_n N_A_500_392#_c_331_n
+ N_A_500_392#_c_332_n N_A_500_392#_c_349_n N_A_500_392#_c_333_n
+ N_A_500_392#_c_334_n N_A_500_392#_c_335_n N_A_500_392#_c_336_n
+ N_A_500_392#_c_359_p N_A_500_392#_c_400_p N_A_500_392#_c_337_n
+ N_A_500_392#_c_371_p N_A_500_392#_c_338_n N_A_500_392#_c_339_n
+ N_A_500_392#_c_382_p N_A_500_392#_c_351_n N_A_500_392#_c_340_n
+ N_A_500_392#_c_341_n N_A_500_392#_c_342_n N_A_500_392#_c_343_n
+ PM_SKY130_FD_SC_LS__DFRBP_1%A_500_392#
x_PM_SKY130_FD_SC_LS__DFRBP_1%A_841_401# N_A_841_401#_M1002_d
+ N_A_841_401#_M1017_d N_A_841_401#_c_539_n N_A_841_401#_M1006_g
+ N_A_841_401#_M1033_g N_A_841_401#_c_540_n N_A_841_401#_c_531_n
+ N_A_841_401#_c_532_n N_A_841_401#_c_533_n N_A_841_401#_c_534_n
+ N_A_841_401#_c_535_n N_A_841_401#_c_536_n N_A_841_401#_c_537_n
+ N_A_841_401#_c_538_n N_A_841_401#_c_544_n
+ PM_SKY130_FD_SC_LS__DFRBP_1%A_841_401#
x_PM_SKY130_FD_SC_LS__DFRBP_1%RESET_B N_RESET_B_M1028_g N_RESET_B_c_642_n
+ N_RESET_B_c_652_n N_RESET_B_c_653_n N_RESET_B_M1022_g N_RESET_B_c_643_n
+ N_RESET_B_c_644_n N_RESET_B_M1015_g N_RESET_B_c_646_n N_RESET_B_c_655_n
+ N_RESET_B_M1019_g N_RESET_B_M1026_g N_RESET_B_c_657_n N_RESET_B_M1014_g
+ N_RESET_B_c_648_n N_RESET_B_c_658_n N_RESET_B_c_659_n N_RESET_B_c_660_n
+ N_RESET_B_c_661_n N_RESET_B_c_662_n N_RESET_B_c_663_n RESET_B
+ N_RESET_B_c_664_n N_RESET_B_c_665_n N_RESET_B_c_649_n N_RESET_B_c_650_n
+ N_RESET_B_c_667_n N_RESET_B_c_668_n PM_SKY130_FD_SC_LS__DFRBP_1%RESET_B
x_PM_SKY130_FD_SC_LS__DFRBP_1%A_705_463# N_A_705_463#_M1013_d
+ N_A_705_463#_M1023_d N_A_705_463#_M1019_d N_A_705_463#_M1002_g
+ N_A_705_463#_c_854_n N_A_705_463#_c_860_n N_A_705_463#_M1017_g
+ N_A_705_463#_c_870_n N_A_705_463#_c_887_n N_A_705_463#_c_861_n
+ N_A_705_463#_c_855_n N_A_705_463#_c_894_n N_A_705_463#_c_856_n
+ N_A_705_463#_c_857_n N_A_705_463#_c_858_n N_A_705_463#_c_864_n
+ PM_SKY130_FD_SC_LS__DFRBP_1%A_705_463#
x_PM_SKY130_FD_SC_LS__DFRBP_1%A_319_392# N_A_319_392#_M1001_s
+ N_A_319_392#_M1000_s N_A_319_392#_M1030_g N_A_319_392#_c_981_n
+ N_A_319_392#_M1029_g N_A_319_392#_c_992_n N_A_319_392#_c_993_n
+ N_A_319_392#_c_994_n N_A_319_392#_c_982_n N_A_319_392#_c_983_n
+ N_A_319_392#_M1013_g N_A_319_392#_c_996_n N_A_319_392#_c_997_n
+ N_A_319_392#_c_998_n N_A_319_392#_M1025_g N_A_319_392#_c_999_n
+ N_A_319_392#_c_1000_n N_A_319_392#_c_1001_n N_A_319_392#_M1012_g
+ N_A_319_392#_c_985_n N_A_319_392#_c_986_n N_A_319_392#_M1032_g
+ N_A_319_392#_c_1005_n N_A_319_392#_c_988_n N_A_319_392#_c_1018_n
+ N_A_319_392#_c_989_n N_A_319_392#_c_990_n N_A_319_392#_c_1007_n
+ PM_SKY130_FD_SC_LS__DFRBP_1%A_319_392#
x_PM_SKY130_FD_SC_LS__DFRBP_1%A_1482_48# N_A_1482_48#_M1027_d
+ N_A_1482_48#_M1014_d N_A_1482_48#_c_1173_n N_A_1482_48#_M1024_g
+ N_A_1482_48#_c_1174_n N_A_1482_48#_c_1182_n N_A_1482_48#_M1016_g
+ N_A_1482_48#_c_1175_n N_A_1482_48#_c_1183_n N_A_1482_48#_c_1176_n
+ N_A_1482_48#_c_1177_n N_A_1482_48#_c_1178_n N_A_1482_48#_c_1185_n
+ N_A_1482_48#_c_1179_n N_A_1482_48#_c_1180_n
+ PM_SKY130_FD_SC_LS__DFRBP_1%A_1482_48#
x_PM_SKY130_FD_SC_LS__DFRBP_1%A_1224_74# N_A_1224_74#_M1004_d
+ N_A_1224_74#_M1012_d N_A_1224_74#_M1027_g N_A_1224_74#_c_1269_n
+ N_A_1224_74#_c_1286_n N_A_1224_74#_M1020_g N_A_1224_74#_c_1270_n
+ N_A_1224_74#_c_1271_n N_A_1224_74#_c_1272_n N_A_1224_74#_M1011_g
+ N_A_1224_74#_M1009_g N_A_1224_74#_c_1274_n N_A_1224_74#_c_1275_n
+ N_A_1224_74#_c_1289_n N_A_1224_74#_M1003_g N_A_1224_74#_M1008_g
+ N_A_1224_74#_c_1277_n N_A_1224_74#_c_1297_n N_A_1224_74#_c_1301_n
+ N_A_1224_74#_c_1278_n N_A_1224_74#_c_1279_n N_A_1224_74#_c_1280_n
+ N_A_1224_74#_c_1281_n N_A_1224_74#_c_1282_n N_A_1224_74#_c_1283_n
+ N_A_1224_74#_c_1284_n PM_SKY130_FD_SC_LS__DFRBP_1%A_1224_74#
x_PM_SKY130_FD_SC_LS__DFRBP_1%A_2026_424# N_A_2026_424#_M1008_s
+ N_A_2026_424#_M1003_s N_A_2026_424#_M1005_g N_A_2026_424#_c_1433_n
+ N_A_2026_424#_M1031_g N_A_2026_424#_c_1434_n N_A_2026_424#_c_1435_n
+ N_A_2026_424#_c_1436_n N_A_2026_424#_c_1437_n
+ PM_SKY130_FD_SC_LS__DFRBP_1%A_2026_424#
x_PM_SKY130_FD_SC_LS__DFRBP_1%VPWR N_VPWR_M1021_s N_VPWR_M1022_d N_VPWR_M1000_d
+ N_VPWR_M1006_d N_VPWR_M1017_s N_VPWR_M1016_d N_VPWR_M1020_d N_VPWR_M1003_d
+ N_VPWR_c_1483_n N_VPWR_c_1484_n N_VPWR_c_1485_n N_VPWR_c_1486_n
+ N_VPWR_c_1487_n N_VPWR_c_1488_n N_VPWR_c_1489_n N_VPWR_c_1490_n
+ N_VPWR_c_1491_n N_VPWR_c_1492_n VPWR N_VPWR_c_1493_n N_VPWR_c_1494_n
+ N_VPWR_c_1495_n N_VPWR_c_1496_n N_VPWR_c_1497_n N_VPWR_c_1498_n
+ N_VPWR_c_1499_n N_VPWR_c_1482_n N_VPWR_c_1501_n N_VPWR_c_1502_n
+ N_VPWR_c_1503_n N_VPWR_c_1504_n N_VPWR_c_1505_n N_VPWR_c_1506_n
+ N_VPWR_c_1507_n PM_SKY130_FD_SC_LS__DFRBP_1%VPWR
x_PM_SKY130_FD_SC_LS__DFRBP_1%A_38_78# N_A_38_78#_M1007_s N_A_38_78#_M1013_s
+ N_A_38_78#_M1021_d N_A_38_78#_M1023_s N_A_38_78#_c_1637_n N_A_38_78#_c_1645_n
+ N_A_38_78#_c_1638_n N_A_38_78#_c_1647_n N_A_38_78#_c_1648_n
+ N_A_38_78#_c_1639_n N_A_38_78#_c_1640_n N_A_38_78#_c_1649_n
+ N_A_38_78#_c_1641_n N_A_38_78#_c_1642_n N_A_38_78#_c_1651_n
+ N_A_38_78#_c_1652_n N_A_38_78#_c_1669_n N_A_38_78#_c_1653_n
+ N_A_38_78#_c_1643_n N_A_38_78#_c_1644_n PM_SKY130_FD_SC_LS__DFRBP_1%A_38_78#
x_PM_SKY130_FD_SC_LS__DFRBP_1%Q_N N_Q_N_M1009_d N_Q_N_M1011_d N_Q_N_c_1770_n Q_N
+ Q_N Q_N N_Q_N_c_1773_n PM_SKY130_FD_SC_LS__DFRBP_1%Q_N
x_PM_SKY130_FD_SC_LS__DFRBP_1%Q N_Q_M1005_d N_Q_M1031_d Q Q Q Q Q N_Q_c_1796_n
+ PM_SKY130_FD_SC_LS__DFRBP_1%Q
x_PM_SKY130_FD_SC_LS__DFRBP_1%VGND N_VGND_M1028_d N_VGND_M1001_d N_VGND_M1015_d
+ N_VGND_M1024_d N_VGND_M1009_s N_VGND_M1008_d N_VGND_c_1817_n N_VGND_c_1818_n
+ N_VGND_c_1819_n N_VGND_c_1820_n N_VGND_c_1821_n N_VGND_c_1822_n VGND
+ N_VGND_c_1823_n N_VGND_c_1824_n N_VGND_c_1825_n N_VGND_c_1826_n
+ N_VGND_c_1827_n N_VGND_c_1828_n N_VGND_c_1829_n N_VGND_c_1830_n
+ N_VGND_c_1831_n N_VGND_c_1832_n N_VGND_c_1833_n N_VGND_c_1834_n
+ N_VGND_c_1835_n PM_SKY130_FD_SC_LS__DFRBP_1%VGND
cc_1 VNB N_D_M1007_g 0.0286427f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.6
cc_2 VNB N_D_c_244_n 0.0408539f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_3 VNB N_D_c_245_n 0.0253354f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_4 VNB N_D_c_246_n 0.0298264f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_5 VNB CLK 0.00260448f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=2.148
cc_6 VNB N_CLK_c_278_n 0.0251051f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_7 VNB N_CLK_c_279_n 0.015704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_500_392#_c_325_n 0.00651136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_500_392#_c_326_n 0.0137458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_500_392#_c_327_n 0.0159053f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.202
cc_11 VNB N_A_500_392#_c_328_n 0.0205313f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.165
cc_12 VNB N_A_500_392#_c_329_n 0.0187502f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1
cc_13 VNB N_A_500_392#_c_330_n 0.00880336f $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.165
cc_14 VNB N_A_500_392#_c_331_n 0.0131415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_500_392#_c_332_n 0.0118314f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.845
cc_16 VNB N_A_500_392#_c_333_n 0.00260346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_500_392#_c_334_n 0.0348735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_500_392#_c_335_n 0.00285435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_500_392#_c_336_n 0.0030846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_500_392#_c_337_n 0.00621215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_500_392#_c_338_n 0.0316981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_500_392#_c_339_n 0.00782104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_500_392#_c_340_n 0.0133198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_500_392#_c_341_n 0.00183605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_500_392#_c_342_n 0.00740079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_500_392#_c_343_n 0.00185238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_841_401#_M1033_g 0.0269879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_841_401#_c_531_n 0.00629371f $X=-0.19 $Y=-0.245 $X2=0.422
+ $Y2=1.165
cc_29 VNB N_A_841_401#_c_532_n 0.0156794f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_30 VNB N_A_841_401#_c_533_n 0.0106545f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1
cc_31 VNB N_A_841_401#_c_534_n 4.52231e-19 $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.165
cc_32 VNB N_A_841_401#_c_535_n 4.96212e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_841_401#_c_536_n 0.00934369f $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.295
cc_34 VNB N_A_841_401#_c_537_n 0.00496873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_841_401#_c_538_n 4.11682e-19 $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.665
cc_36 VNB N_RESET_B_M1028_g 0.0222763f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1
cc_37 VNB N_RESET_B_c_642_n 0.0275892f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.6
cc_38 VNB N_RESET_B_c_643_n 0.286034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_RESET_B_c_644_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_RESET_B_M1015_g 0.0240189f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_41 VNB N_RESET_B_c_646_n 0.01872f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.165
cc_42 VNB N_RESET_B_M1026_g 0.0515393f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.295
cc_43 VNB N_RESET_B_c_648_n 0.0133121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_RESET_B_c_649_n 0.0323124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_RESET_B_c_650_n 0.00371377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_705_463#_M1002_g 0.0297973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_705_463#_c_854_n 0.0206988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_705_463#_c_855_n 0.00342048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_705_463#_c_856_n 0.00364311f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_705_463#_c_857_n 0.0106366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_705_463#_c_858_n 0.0286964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_319_392#_c_981_n 0.0149901f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_53 VNB N_A_319_392#_c_982_n 0.0301015f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_54 VNB N_A_319_392#_c_983_n 0.0627365f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.165
cc_55 VNB N_A_319_392#_M1013_g 0.0225997f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1
cc_56 VNB N_A_319_392#_c_985_n 0.021569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_319_392#_c_986_n 0.00563426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_319_392#_M1032_g 0.0529012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_319_392#_c_988_n 0.00845639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_319_392#_c_989_n 9.79491e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_319_392#_c_990_n 0.010025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1482_48#_c_1173_n 0.0177983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1482_48#_c_1174_n 0.0233363f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_64 VNB N_A_1482_48#_c_1175_n 0.0157083f $X=-0.19 $Y=-0.245 $X2=0.422
+ $Y2=1.202
cc_65 VNB N_A_1482_48#_c_1176_n 0.0117659f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_66 VNB N_A_1482_48#_c_1177_n 0.00518085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1482_48#_c_1178_n 0.00346875f $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.295
cc_68 VNB N_A_1482_48#_c_1179_n 0.00600532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1482_48#_c_1180_n 0.0330587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1224_74#_M1027_g 0.0408739f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_71 VNB N_A_1224_74#_c_1269_n 0.00400132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1224_74#_c_1270_n 0.0327014f $X=-0.19 $Y=-0.245 $X2=0.422
+ $Y2=1.845
cc_73 VNB N_A_1224_74#_c_1271_n 0.0281282f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.845
cc_74 VNB N_A_1224_74#_c_1272_n 0.0364438f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.845
cc_75 VNB N_A_1224_74#_M1009_g 0.0260029f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.165
cc_76 VNB N_A_1224_74#_c_1274_n 0.0888375f $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.295
cc_77 VNB N_A_1224_74#_c_1275_n 0.00400127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1224_74#_M1008_g 0.0355065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1224_74#_c_1277_n 0.0100839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1224_74#_c_1278_n 0.00749917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1224_74#_c_1279_n 0.0120508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1224_74#_c_1280_n 4.69525e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1224_74#_c_1281_n 9.056e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1224_74#_c_1282_n 0.00965329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1224_74#_c_1283_n 5.50055e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1224_74#_c_1284_n 0.00638783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2026_424#_M1005_g 0.0282052f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_88 VNB N_A_2026_424#_c_1433_n 0.0344608f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_89 VNB N_A_2026_424#_c_1434_n 0.00968545f $X=-0.19 $Y=-0.245 $X2=0.422
+ $Y2=1.845
cc_90 VNB N_A_2026_424#_c_1435_n 3.04122e-19 $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_91 VNB N_A_2026_424#_c_1436_n 0.00611923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2026_424#_c_1437_n 3.73161e-19 $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.665
cc_93 VNB N_VPWR_c_1482_n 0.48212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_38_78#_c_1637_n 0.00234225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_38_78#_c_1638_n 0.0151383f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_96 VNB N_A_38_78#_c_1639_n 9.8117e-19 $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.845
cc_97 VNB N_A_38_78#_c_1640_n 0.00164254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_38_78#_c_1641_n 0.00370394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_38_78#_c_1642_n 0.0222631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_38_78#_c_1643_n 5.71893e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_38_78#_c_1644_n 0.00608917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_Q_N_c_1770_n 0.0157896f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_103 VNB Q 0.0267746f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_104 VNB Q 0.0133985f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_105 VNB N_Q_c_1796_n 0.0249767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1817_n 0.00940183f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_107 VNB N_VGND_c_1818_n 0.021454f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.165
cc_108 VNB N_VGND_c_1819_n 0.0132166f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.665
cc_109 VNB N_VGND_c_1820_n 0.00450041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1821_n 0.00944343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1822_n 0.0125104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1823_n 0.0298733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1824_n 0.0605658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1825_n 0.0603291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1826_n 0.0324414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1827_n 0.0347338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1828_n 0.0191572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1829_n 0.609762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1830_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1831_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1832_n 0.0146905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1833_n 0.00846888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1834_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1835_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VPB N_D_c_247_n 0.017902f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.465
cc_126 VPB N_D_c_248_n 0.0399063f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.148
cc_127 VPB N_D_c_244_n 0.0435358f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_128 VPB N_D_c_246_n 0.0215212f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_129 VPB N_CLK_M1000_g 0.0242864f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_130 VPB CLK 0.00380331f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.148
cc_131 VPB N_CLK_c_278_n 0.0133323f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_132 VPB N_A_500_392#_c_325_n 0.0290243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_500_392#_c_345_n 0.00848422f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.148
cc_134 VPB N_A_500_392#_c_326_n 0.0211535f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_500_392#_c_347_n 0.0569971f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_500_392#_c_348_n 0.0211542f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.665
cc_137 VPB N_A_500_392#_c_349_n 0.00500505f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=2.035
cc_138 VPB N_A_500_392#_c_339_n 0.0024834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_500_392#_c_351_n 0.00306084f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_500_392#_c_341_n 0.0021357f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_841_401#_c_539_n 0.0145107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_841_401#_c_540_n 0.0553568f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_841_401#_c_531_n 0.00229128f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.165
cc_144 VPB N_A_841_401#_c_532_n 0.00204604f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_145 VPB N_A_841_401#_c_537_n 6.92353e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_841_401#_c_544_n 0.00398554f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=2.035
cc_147 VPB N_RESET_B_c_642_n 0.0231877f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=0.6
cc_148 VPB N_RESET_B_c_652_n 0.0161426f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.148
cc_149 VPB N_RESET_B_c_653_n 0.0239078f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_150 VPB N_RESET_B_c_646_n 0.0124021f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.165
cc_151 VPB N_RESET_B_c_655_n 0.0191525f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_152 VPB N_RESET_B_M1026_g 0.00974243f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.295
cc_153 VPB N_RESET_B_c_657_n 0.052471f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.665
cc_154 VPB N_RESET_B_c_658_n 0.0189061f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_RESET_B_c_659_n 0.0277252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_RESET_B_c_660_n 0.00333626f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_RESET_B_c_661_n 0.00537181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_RESET_B_c_662_n 0.00350644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_RESET_B_c_663_n 0.00338092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_RESET_B_c_664_n 0.0553546f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_RESET_B_c_665_n 0.00383188f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_RESET_B_c_650_n 9.2757e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_RESET_B_c_667_n 0.0291728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_RESET_B_c_668_n 0.00608672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_705_463#_c_854_n 0.0214001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_705_463#_c_860_n 0.0168657f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.845
cc_167 VPB N_A_705_463#_c_861_n 0.0113023f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_705_463#_c_856_n 0.00939076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_705_463#_c_858_n 3.30851e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_705_463#_c_864_n 0.00604136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_319_392#_M1030_g 0.0214513f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_172 VPB N_A_319_392#_c_992_n 0.0745734f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.202
cc_173 VPB N_A_319_392#_c_993_n 0.0553482f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.845
cc_174 VPB N_A_319_392#_c_994_n 0.012371f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_175 VPB N_A_319_392#_c_983_n 0.0140094f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.165
cc_176 VPB N_A_319_392#_c_996_n 0.00710611f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_319_392#_c_997_n 0.0163876f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.295
cc_178 VPB N_A_319_392#_c_998_n 0.0140534f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_319_392#_c_999_n 0.200724f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.845
cc_180 VPB N_A_319_392#_c_1000_n 0.00738389f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_319_392#_c_1001_n 0.0161081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_319_392#_M1012_g 0.00837835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_319_392#_c_985_n 0.0142262f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_319_392#_c_986_n 0.00505238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_319_392#_c_1005_n 0.0089864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_319_392#_c_988_n 0.0038387f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_319_392#_c_1007_n 0.0126952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_1482_48#_c_1174_n 0.0272407f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_189 VPB N_A_1482_48#_c_1182_n 0.0213103f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1482_48#_c_1183_n 0.0103983f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_191 VPB N_A_1482_48#_c_1177_n 0.00239847f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_1482_48#_c_1185_n 0.00655902f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_1224_74#_c_1269_n 0.0278194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1224_74#_c_1286_n 0.021316f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_1224_74#_c_1272_n 0.0280594f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_196 VPB N_A_1224_74#_c_1275_n 0.0203227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1224_74#_c_1289_n 0.0278562f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.845
cc_198 VPB N_A_1224_74#_c_1281_n 0.00656652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_2026_424#_c_1433_n 0.0290451f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_200 VPB N_A_2026_424#_c_1435_n 0.00753336f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.165
cc_201 VPB N_VPWR_c_1483_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.295
cc_202 VPB N_VPWR_c_1484_n 0.0307191f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.665
cc_203 VPB N_VPWR_c_1485_n 0.010025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1486_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1487_n 0.0139231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1488_n 0.0156795f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1489_n 0.0249508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1490_n 0.021993f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1491_n 0.0118234f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1492_n 0.0143642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1493_n 0.0176642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1494_n 0.0189818f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1495_n 0.0579816f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1496_n 0.0280581f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1497_n 0.0507873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1498_n 0.0430282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1499_n 0.0189171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1482_n 0.120841f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1501_n 0.00614052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1502_n 0.00601569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1503_n 0.00456844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1504_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1505_n 0.00430193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1506_n 0.00410958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1507_n 0.00564836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_38_78#_c_1645_n 0.00241568f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_227 VPB N_A_38_78#_c_1638_n 0.0107846f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_228 VPB N_A_38_78#_c_1647_n 0.0105441f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_229 VPB N_A_38_78#_c_1648_n 0.00305134f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.295
cc_230 VPB N_A_38_78#_c_1649_n 5.84114e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_38_78#_c_1641_n 0.00678795f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_38_78#_c_1651_n 0.00547968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_38_78#_c_1652_n 0.00193012f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_38_78#_c_1653_n 0.00388249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_Q_N_c_1770_n 0.00323856f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_236 VPB Q_N 0.0168178f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_Q_N_c_1773_n 0.00844312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB Q 0.0131162f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_239 VPB Q 0.041687f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.665
cc_240 VPB N_Q_c_1796_n 0.00776073f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 N_D_M1007_g N_RESET_B_M1028_g 0.0261166f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_242 N_D_c_244_n N_RESET_B_c_642_n 0.0261166f $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_243 N_D_c_248_n N_RESET_B_c_652_n 0.00488452f $X=0.422 $Y=2.148 $X2=0 $Y2=0
cc_244 N_D_c_247_n N_RESET_B_c_653_n 0.00893417f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_245 N_D_c_245_n N_RESET_B_c_649_n 0.0261166f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_246 N_D_c_248_n N_RESET_B_c_667_n 0.0261166f $X=0.422 $Y=2.148 $X2=0 $Y2=0
cc_247 N_D_c_247_n N_VPWR_c_1484_n 0.00598914f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_248 N_D_c_248_n N_VPWR_c_1484_n 0.0042702f $X=0.422 $Y=2.148 $X2=0 $Y2=0
cc_249 N_D_c_246_n N_VPWR_c_1484_n 0.013492f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_250 N_D_c_247_n N_VPWR_c_1485_n 4.12155e-19 $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_251 N_D_c_247_n N_VPWR_c_1493_n 0.00445602f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_252 N_D_c_247_n N_VPWR_c_1482_n 0.00861168f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_253 N_D_c_248_n N_VPWR_c_1482_n 3.7828e-19 $X=0.422 $Y=2.148 $X2=0 $Y2=0
cc_254 N_D_M1007_g N_A_38_78#_c_1637_n 0.0116103f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_255 N_D_c_246_n N_A_38_78#_c_1637_n 0.00144733f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_256 N_D_c_247_n N_A_38_78#_c_1645_n 0.00424962f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_257 N_D_M1007_g N_A_38_78#_c_1638_n 0.0152564f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_258 N_D_c_246_n N_A_38_78#_c_1638_n 0.0904243f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_259 N_D_M1007_g N_A_38_78#_c_1642_n 0.0078958f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_260 N_D_c_245_n N_A_38_78#_c_1642_n 0.00191909f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_261 N_D_c_246_n N_A_38_78#_c_1642_n 0.028486f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_262 N_D_c_247_n N_A_38_78#_c_1651_n 0.00395363f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_263 N_D_c_248_n N_A_38_78#_c_1651_n 0.00689915f $X=0.422 $Y=2.148 $X2=0 $Y2=0
cc_264 N_D_M1007_g N_VGND_c_1817_n 0.00200808f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_265 N_D_M1007_g N_VGND_c_1823_n 0.00429844f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_266 N_D_M1007_g N_VGND_c_1829_n 0.00539454f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_267 N_CLK_M1000_g N_A_500_392#_c_349_n 0.00122372f $X=1.965 $Y=2.46 $X2=0
+ $Y2=0
cc_268 N_CLK_M1000_g N_RESET_B_c_642_n 0.00463279f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_269 N_CLK_c_278_n N_RESET_B_c_642_n 0.00731548f $X=1.975 $Y=1.61 $X2=0 $Y2=0
cc_270 N_CLK_c_279_n N_RESET_B_c_643_n 0.0103009f $X=1.962 $Y=1.41 $X2=0 $Y2=0
cc_271 N_CLK_M1000_g N_RESET_B_c_659_n 0.00470044f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_272 CLK N_RESET_B_c_659_n 0.0160477f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_273 N_CLK_c_278_n N_RESET_B_c_659_n 0.00170548f $X=1.975 $Y=1.61 $X2=0 $Y2=0
cc_274 N_CLK_c_279_n N_RESET_B_c_649_n 0.00394671f $X=1.962 $Y=1.41 $X2=0 $Y2=0
cc_275 CLK N_A_319_392#_M1001_s 5.47303e-19 $X=2.075 $Y=1.58 $X2=-0.19
+ $Y2=-0.245
cc_276 N_CLK_M1000_g N_A_319_392#_M1030_g 0.0413937f $X=1.965 $Y=2.46 $X2=0
+ $Y2=0
cc_277 CLK N_A_319_392#_c_981_n 3.85296e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_278 N_CLK_c_279_n N_A_319_392#_c_981_n 0.0217488f $X=1.962 $Y=1.41 $X2=0
+ $Y2=0
cc_279 CLK N_A_319_392#_c_983_n 0.0044164f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_280 N_CLK_c_278_n N_A_319_392#_c_983_n 0.0238169f $X=1.975 $Y=1.61 $X2=0
+ $Y2=0
cc_281 N_CLK_M1000_g N_A_319_392#_c_988_n 0.00181991f $X=1.965 $Y=2.46 $X2=0
+ $Y2=0
cc_282 CLK N_A_319_392#_c_988_n 0.0334879f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_283 N_CLK_c_278_n N_A_319_392#_c_988_n 0.00341993f $X=1.975 $Y=1.61 $X2=0
+ $Y2=0
cc_284 N_CLK_c_279_n N_A_319_392#_c_988_n 0.00388687f $X=1.962 $Y=1.41 $X2=0
+ $Y2=0
cc_285 N_CLK_c_278_n N_A_319_392#_c_1018_n 4.13834e-19 $X=1.975 $Y=1.61 $X2=0
+ $Y2=0
cc_286 N_CLK_c_279_n N_A_319_392#_c_1018_n 0.0115337f $X=1.962 $Y=1.41 $X2=0
+ $Y2=0
cc_287 CLK N_A_319_392#_c_989_n 0.0294479f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_288 N_CLK_c_278_n N_A_319_392#_c_989_n 2.33973e-19 $X=1.975 $Y=1.61 $X2=0
+ $Y2=0
cc_289 CLK N_A_319_392#_c_990_n 0.0270662f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_290 N_CLK_c_278_n N_A_319_392#_c_990_n 0.00134844f $X=1.975 $Y=1.61 $X2=0
+ $Y2=0
cc_291 N_CLK_c_279_n N_A_319_392#_c_990_n 0.0101268f $X=1.962 $Y=1.41 $X2=0
+ $Y2=0
cc_292 N_CLK_M1000_g N_A_319_392#_c_1007_n 0.00429385f $X=1.965 $Y=2.46 $X2=0
+ $Y2=0
cc_293 CLK N_A_319_392#_c_1007_n 0.00114171f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_294 N_CLK_c_278_n N_A_319_392#_c_1007_n 0.00152253f $X=1.975 $Y=1.61 $X2=0
+ $Y2=0
cc_295 N_CLK_M1000_g N_VPWR_c_1485_n 0.00847466f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_296 N_CLK_M1000_g N_VPWR_c_1486_n 0.0164741f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_297 N_CLK_M1000_g N_VPWR_c_1494_n 0.00303184f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_298 N_CLK_M1000_g N_VPWR_c_1482_n 0.00397656f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_299 N_CLK_M1000_g N_A_38_78#_c_1647_n 0.00307891f $X=1.965 $Y=2.46 $X2=0
+ $Y2=0
cc_300 N_CLK_M1000_g N_A_38_78#_c_1648_n 0.00630143f $X=1.965 $Y=2.46 $X2=0
+ $Y2=0
cc_301 CLK N_A_38_78#_c_1648_n 0.00252085f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_302 N_CLK_c_278_n N_A_38_78#_c_1648_n 3.06088e-19 $X=1.975 $Y=1.61 $X2=0
+ $Y2=0
cc_303 N_CLK_c_278_n N_A_38_78#_c_1652_n 9.45729e-19 $X=1.975 $Y=1.61 $X2=0
+ $Y2=0
cc_304 N_CLK_M1000_g N_A_38_78#_c_1669_n 0.00870954f $X=1.965 $Y=2.46 $X2=0
+ $Y2=0
cc_305 CLK N_VGND_M1001_d 0.00211522f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_306 N_CLK_c_279_n N_VGND_c_1817_n 0.00347693f $X=1.962 $Y=1.41 $X2=0 $Y2=0
cc_307 N_CLK_c_279_n N_VGND_c_1819_n 0.00506085f $X=1.962 $Y=1.41 $X2=0 $Y2=0
cc_308 N_CLK_c_279_n N_VGND_c_1829_n 9.39239e-19 $X=1.962 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A_500_392#_c_336_n N_A_841_401#_M1002_d 0.0095109f $X=6.085 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_310 N_A_500_392#_c_327_n N_A_841_401#_M1033_g 0.00963625f $X=4.015 $Y=1.56
+ $X2=0 $Y2=0
cc_311 N_A_500_392#_c_331_n N_A_841_401#_M1033_g 0.0408829f $X=4.05 $Y=1.09
+ $X2=0 $Y2=0
cc_312 N_A_500_392#_c_335_n N_A_841_401#_M1033_g 0.00423512f $X=4.435 $Y=0.58
+ $X2=0 $Y2=0
cc_313 N_A_500_392#_c_336_n N_A_841_401#_M1033_g 0.00295293f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_314 N_A_500_392#_c_359_p N_A_841_401#_M1033_g 0.00422261f $X=4.52 $Y=0.665
+ $X2=0 $Y2=0
cc_315 N_A_500_392#_c_345_n N_A_841_401#_c_540_n 0.0024818f $X=3.462 $Y=2.123
+ $X2=0 $Y2=0
cc_316 N_A_500_392#_c_326_n N_A_841_401#_c_540_n 0.00696445f $X=3.94 $Y=1.635
+ $X2=0 $Y2=0
cc_317 N_A_500_392#_c_327_n N_A_841_401#_c_531_n 9.08379e-19 $X=4.015 $Y=1.56
+ $X2=0 $Y2=0
cc_318 N_A_500_392#_c_332_n N_A_841_401#_c_531_n 4.69143e-19 $X=4.05 $Y=1.24
+ $X2=0 $Y2=0
cc_319 N_A_500_392#_c_327_n N_A_841_401#_c_532_n 0.00696445f $X=4.015 $Y=1.56
+ $X2=0 $Y2=0
cc_320 N_A_500_392#_c_336_n N_A_841_401#_c_533_n 0.0628972f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_321 N_A_500_392#_c_331_n N_A_841_401#_c_534_n 3.46091e-19 $X=4.05 $Y=1.09
+ $X2=0 $Y2=0
cc_322 N_A_500_392#_c_336_n N_A_841_401#_c_534_n 0.00412245f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_323 N_A_500_392#_c_359_p N_A_841_401#_c_534_n 0.00983586f $X=4.52 $Y=0.665
+ $X2=0 $Y2=0
cc_324 N_A_500_392#_c_328_n N_A_841_401#_c_535_n 0.00136384f $X=6.045 $Y=1.085
+ $X2=0 $Y2=0
cc_325 N_A_500_392#_c_336_n N_A_841_401#_c_535_n 0.0136179f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_326 N_A_500_392#_c_371_p N_A_841_401#_c_535_n 0.0108515f $X=6.255 $Y=1.065
+ $X2=0 $Y2=0
cc_327 N_A_500_392#_c_330_n N_A_841_401#_c_536_n 0.00176493f $X=6.12 $Y=1.16
+ $X2=0 $Y2=0
cc_328 N_A_500_392#_c_371_p N_A_841_401#_c_536_n 0.011149f $X=6.255 $Y=1.065
+ $X2=0 $Y2=0
cc_329 N_A_500_392#_c_329_n N_A_841_401#_c_537_n 0.00507154f $X=6.48 $Y=1.16
+ $X2=0 $Y2=0
cc_330 N_A_500_392#_c_330_n N_A_841_401#_c_537_n 0.00303743f $X=6.12 $Y=1.16
+ $X2=0 $Y2=0
cc_331 N_A_500_392#_c_336_n N_A_841_401#_c_537_n 0.00373373f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_332 N_A_500_392#_c_337_n N_A_841_401#_c_537_n 0.0188995f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_333 N_A_500_392#_c_371_p N_A_841_401#_c_537_n 0.0136879f $X=6.255 $Y=1.065
+ $X2=0 $Y2=0
cc_334 N_A_500_392#_c_339_n N_A_841_401#_c_537_n 0.0135711f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_335 N_A_500_392#_c_347_n N_A_841_401#_c_544_n 0.00141721f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_336 N_A_500_392#_c_339_n N_A_841_401#_c_544_n 0.016501f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_337 N_A_500_392#_c_382_p N_A_841_401#_c_544_n 0.0140459f $X=6.82 $Y=2.03
+ $X2=0 $Y2=0
cc_338 N_A_500_392#_c_331_n N_RESET_B_c_643_n 0.00882199f $X=4.05 $Y=1.09 $X2=0
+ $Y2=0
cc_339 N_A_500_392#_c_334_n N_RESET_B_c_643_n 0.0261266f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_340 N_A_500_392#_c_336_n N_RESET_B_c_643_n 0.00286781f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_341 N_A_500_392#_c_340_n N_RESET_B_c_643_n 0.0121156f $X=2.862 $Y=0.34 $X2=0
+ $Y2=0
cc_342 N_A_500_392#_c_334_n N_RESET_B_M1015_g 0.00386847f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_343 N_A_500_392#_c_335_n N_RESET_B_M1015_g 0.00191339f $X=4.435 $Y=0.58 $X2=0
+ $Y2=0
cc_344 N_A_500_392#_c_336_n N_RESET_B_M1015_g 0.012028f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_345 N_A_500_392#_c_325_n N_RESET_B_c_659_n 9.88559e-19 $X=3.462 $Y=1.985
+ $X2=0 $Y2=0
cc_346 N_A_500_392#_c_345_n N_RESET_B_c_659_n 0.0035746f $X=3.462 $Y=2.123 $X2=0
+ $Y2=0
cc_347 N_A_500_392#_c_326_n N_RESET_B_c_659_n 0.00511381f $X=3.94 $Y=1.635 $X2=0
+ $Y2=0
cc_348 N_A_500_392#_c_349_n N_RESET_B_c_659_n 0.024703f $X=2.915 $Y=2.052 $X2=0
+ $Y2=0
cc_349 N_A_500_392#_c_341_n N_RESET_B_c_659_n 0.0266841f $X=3.385 $Y=1.82 $X2=0
+ $Y2=0
cc_350 N_A_500_392#_c_347_n N_RESET_B_c_661_n 0.00152844f $X=7.25 $Y=2.28 $X2=0
+ $Y2=0
cc_351 N_A_500_392#_c_382_p N_RESET_B_c_661_n 0.0123453f $X=6.82 $Y=2.03 $X2=0
+ $Y2=0
cc_352 N_A_500_392#_c_351_n N_RESET_B_c_661_n 0.0237639f $X=7.205 $Y=2.03 $X2=0
+ $Y2=0
cc_353 N_A_500_392#_c_328_n N_A_705_463#_M1002_g 0.0261676f $X=6.045 $Y=1.085
+ $X2=0 $Y2=0
cc_354 N_A_500_392#_c_336_n N_A_705_463#_M1002_g 0.0128398f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_355 N_A_500_392#_c_400_p N_A_705_463#_M1002_g 6.89487e-19 $X=6.17 $Y=0.9
+ $X2=0 $Y2=0
cc_356 N_A_500_392#_c_371_p N_A_705_463#_M1002_g 2.33891e-19 $X=6.255 $Y=1.065
+ $X2=0 $Y2=0
cc_357 N_A_500_392#_c_330_n N_A_705_463#_c_854_n 0.0123428f $X=6.12 $Y=1.16
+ $X2=0 $Y2=0
cc_358 N_A_500_392#_c_348_n N_A_705_463#_c_870_n 0.00177991f $X=3.462 $Y=2.21
+ $X2=0 $Y2=0
cc_359 N_A_500_392#_c_326_n N_A_705_463#_c_855_n 0.00263818f $X=3.94 $Y=1.635
+ $X2=0 $Y2=0
cc_360 N_A_500_392#_c_331_n N_A_705_463#_c_855_n 0.00935232f $X=4.05 $Y=1.09
+ $X2=0 $Y2=0
cc_361 N_A_500_392#_c_332_n N_A_705_463#_c_855_n 0.00354155f $X=4.05 $Y=1.24
+ $X2=0 $Y2=0
cc_362 N_A_500_392#_c_334_n N_A_705_463#_c_855_n 0.0317578f $X=4.35 $Y=0.34
+ $X2=0 $Y2=0
cc_363 N_A_500_392#_c_326_n N_A_705_463#_c_856_n 0.00575936f $X=3.94 $Y=1.635
+ $X2=0 $Y2=0
cc_364 N_A_500_392#_c_327_n N_A_705_463#_c_856_n 0.00639358f $X=4.015 $Y=1.56
+ $X2=0 $Y2=0
cc_365 N_A_500_392#_c_348_n N_A_705_463#_c_856_n 5.44904e-19 $X=3.462 $Y=2.21
+ $X2=0 $Y2=0
cc_366 N_A_500_392#_c_331_n N_A_705_463#_c_856_n 0.00254473f $X=4.05 $Y=1.09
+ $X2=0 $Y2=0
cc_367 N_A_500_392#_c_332_n N_A_705_463#_c_856_n 0.00590609f $X=4.05 $Y=1.24
+ $X2=0 $Y2=0
cc_368 N_A_500_392#_c_349_n N_A_319_392#_M1030_g 0.00867095f $X=2.915 $Y=2.052
+ $X2=0 $Y2=0
cc_369 N_A_500_392#_c_341_n N_A_319_392#_M1030_g 4.53138e-19 $X=3.385 $Y=1.82
+ $X2=0 $Y2=0
cc_370 N_A_500_392#_c_340_n N_A_319_392#_c_981_n 0.00671343f $X=2.862 $Y=0.34
+ $X2=0 $Y2=0
cc_371 N_A_500_392#_c_342_n N_A_319_392#_c_981_n 0.00489626f $X=3.052 $Y=1.205
+ $X2=0 $Y2=0
cc_372 N_A_500_392#_c_345_n N_A_319_392#_c_992_n 0.0219381f $X=3.462 $Y=2.123
+ $X2=0 $Y2=0
cc_373 N_A_500_392#_c_349_n N_A_319_392#_c_992_n 0.0105467f $X=2.915 $Y=2.052
+ $X2=0 $Y2=0
cc_374 N_A_500_392#_c_341_n N_A_319_392#_c_992_n 0.0129859f $X=3.385 $Y=1.82
+ $X2=0 $Y2=0
cc_375 N_A_500_392#_c_348_n N_A_319_392#_c_993_n 0.0103742f $X=3.462 $Y=2.21
+ $X2=0 $Y2=0
cc_376 N_A_500_392#_c_325_n N_A_319_392#_c_982_n 0.0250228f $X=3.462 $Y=1.985
+ $X2=0 $Y2=0
cc_377 N_A_500_392#_c_327_n N_A_319_392#_c_982_n 0.00530535f $X=4.015 $Y=1.56
+ $X2=0 $Y2=0
cc_378 N_A_500_392#_c_341_n N_A_319_392#_c_982_n 0.00439047f $X=3.385 $Y=1.82
+ $X2=0 $Y2=0
cc_379 N_A_500_392#_c_343_n N_A_319_392#_c_982_n 0.00304316f $X=3.052 $Y=1.39
+ $X2=0 $Y2=0
cc_380 N_A_500_392#_c_325_n N_A_319_392#_c_983_n 0.0249579f $X=3.462 $Y=1.985
+ $X2=0 $Y2=0
cc_381 N_A_500_392#_c_349_n N_A_319_392#_c_983_n 0.00475108f $X=2.915 $Y=2.052
+ $X2=0 $Y2=0
cc_382 N_A_500_392#_c_333_n N_A_319_392#_c_983_n 0.0103033f $X=3.067 $Y=1.575
+ $X2=0 $Y2=0
cc_383 N_A_500_392#_c_340_n N_A_319_392#_c_983_n 0.00550214f $X=2.862 $Y=0.34
+ $X2=0 $Y2=0
cc_384 N_A_500_392#_c_341_n N_A_319_392#_c_983_n 0.00840174f $X=3.385 $Y=1.82
+ $X2=0 $Y2=0
cc_385 N_A_500_392#_c_342_n N_A_319_392#_c_983_n 0.00298161f $X=3.052 $Y=1.205
+ $X2=0 $Y2=0
cc_386 N_A_500_392#_c_343_n N_A_319_392#_c_983_n 0.00724742f $X=3.052 $Y=1.39
+ $X2=0 $Y2=0
cc_387 N_A_500_392#_c_331_n N_A_319_392#_M1013_g 0.0129436f $X=4.05 $Y=1.09
+ $X2=0 $Y2=0
cc_388 N_A_500_392#_c_332_n N_A_319_392#_M1013_g 0.00530535f $X=4.05 $Y=1.24
+ $X2=0 $Y2=0
cc_389 N_A_500_392#_c_334_n N_A_319_392#_M1013_g 0.00330666f $X=4.35 $Y=0.34
+ $X2=0 $Y2=0
cc_390 N_A_500_392#_c_340_n N_A_319_392#_M1013_g 0.00563626f $X=2.862 $Y=0.34
+ $X2=0 $Y2=0
cc_391 N_A_500_392#_c_348_n N_A_319_392#_c_996_n 0.00274475f $X=3.462 $Y=2.21
+ $X2=0 $Y2=0
cc_392 N_A_500_392#_c_326_n N_A_319_392#_c_998_n 0.00408019f $X=3.94 $Y=1.635
+ $X2=0 $Y2=0
cc_393 N_A_500_392#_c_348_n N_A_319_392#_c_998_n 0.0127077f $X=3.462 $Y=2.21
+ $X2=0 $Y2=0
cc_394 N_A_500_392#_c_347_n N_A_319_392#_c_1000_n 0.002647f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_395 N_A_500_392#_c_347_n N_A_319_392#_M1012_g 0.0194051f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_396 N_A_500_392#_c_339_n N_A_319_392#_M1012_g 0.0042093f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_397 N_A_500_392#_c_382_p N_A_319_392#_M1012_g 0.00216411f $X=6.82 $Y=2.03
+ $X2=0 $Y2=0
cc_398 N_A_500_392#_c_347_n N_A_319_392#_c_985_n 0.00720172f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_399 N_A_500_392#_c_338_n N_A_319_392#_c_985_n 0.0103797f $X=6.645 $Y=1.065
+ $X2=0 $Y2=0
cc_400 N_A_500_392#_c_339_n N_A_319_392#_c_985_n 0.0123591f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_401 N_A_500_392#_c_351_n N_A_319_392#_c_985_n 0.00746766f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_402 N_A_500_392#_c_329_n N_A_319_392#_c_986_n 0.0103797f $X=6.48 $Y=1.16
+ $X2=0 $Y2=0
cc_403 N_A_500_392#_c_337_n N_A_319_392#_c_986_n 0.00126209f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_404 N_A_500_392#_c_339_n N_A_319_392#_c_986_n 8.31237e-19 $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_405 N_A_500_392#_c_337_n N_A_319_392#_M1032_g 0.00116888f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_406 N_A_500_392#_c_338_n N_A_319_392#_M1032_g 0.0216896f $X=6.645 $Y=1.065
+ $X2=0 $Y2=0
cc_407 N_A_500_392#_c_339_n N_A_319_392#_M1032_g 0.00159607f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_408 N_A_500_392#_M1029_d N_A_319_392#_c_1018_n 0.00286138f $X=2.625 $Y=0.595
+ $X2=0 $Y2=0
cc_409 N_A_500_392#_c_340_n N_A_319_392#_c_1018_n 0.00942134f $X=2.862 $Y=0.34
+ $X2=0 $Y2=0
cc_410 N_A_500_392#_c_342_n N_A_319_392#_c_1018_n 0.0138589f $X=3.052 $Y=1.205
+ $X2=0 $Y2=0
cc_411 N_A_500_392#_M1029_d N_A_319_392#_c_989_n 0.00180711f $X=2.625 $Y=0.595
+ $X2=0 $Y2=0
cc_412 N_A_500_392#_c_349_n N_A_319_392#_c_989_n 0.0256873f $X=2.915 $Y=2.052
+ $X2=0 $Y2=0
cc_413 N_A_500_392#_c_333_n N_A_319_392#_c_989_n 0.0124651f $X=3.067 $Y=1.575
+ $X2=0 $Y2=0
cc_414 N_A_500_392#_c_341_n N_A_319_392#_c_989_n 0.00943288f $X=3.385 $Y=1.82
+ $X2=0 $Y2=0
cc_415 N_A_500_392#_c_342_n N_A_319_392#_c_989_n 0.0196963f $X=3.052 $Y=1.205
+ $X2=0 $Y2=0
cc_416 N_A_500_392#_c_349_n N_A_319_392#_c_1007_n 0.00812144f $X=2.915 $Y=2.052
+ $X2=0 $Y2=0
cc_417 N_A_500_392#_c_347_n N_A_1482_48#_c_1174_n 0.0212122f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_418 N_A_500_392#_c_351_n N_A_1482_48#_c_1174_n 4.05192e-19 $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_419 N_A_500_392#_c_347_n N_A_1482_48#_c_1182_n 0.0335632f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_420 N_A_500_392#_c_336_n N_A_1224_74#_M1004_d 0.00392413f $X=6.085 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_421 N_A_500_392#_c_400_p N_A_1224_74#_M1004_d 0.00564702f $X=6.17 $Y=0.9
+ $X2=-0.19 $Y2=-0.245
cc_422 N_A_500_392#_c_337_n N_A_1224_74#_M1004_d 0.00471261f $X=6.65 $Y=1.065
+ $X2=-0.19 $Y2=-0.245
cc_423 N_A_500_392#_c_339_n N_A_1224_74#_M1012_d 0.00321319f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_424 N_A_500_392#_c_382_p N_A_1224_74#_M1012_d 0.00528653f $X=6.82 $Y=2.03
+ $X2=0 $Y2=0
cc_425 N_A_500_392#_c_351_n N_A_1224_74#_M1012_d 0.00213077f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_426 N_A_500_392#_c_328_n N_A_1224_74#_c_1297_n 0.00722906f $X=6.045 $Y=1.085
+ $X2=0 $Y2=0
cc_427 N_A_500_392#_c_336_n N_A_1224_74#_c_1297_n 0.013434f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_428 N_A_500_392#_c_337_n N_A_1224_74#_c_1297_n 0.0317086f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_429 N_A_500_392#_c_338_n N_A_1224_74#_c_1297_n 0.00506999f $X=6.645 $Y=1.065
+ $X2=0 $Y2=0
cc_430 N_A_500_392#_c_347_n N_A_1224_74#_c_1301_n 0.0215946f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_431 N_A_500_392#_c_382_p N_A_1224_74#_c_1301_n 0.00944134f $X=6.82 $Y=2.03
+ $X2=0 $Y2=0
cc_432 N_A_500_392#_c_351_n N_A_1224_74#_c_1301_n 0.0346045f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_433 N_A_500_392#_c_337_n N_A_1224_74#_c_1278_n 0.0278616f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_434 N_A_500_392#_c_338_n N_A_1224_74#_c_1278_n 9.55385e-19 $X=6.645 $Y=1.065
+ $X2=0 $Y2=0
cc_435 N_A_500_392#_c_339_n N_A_1224_74#_c_1278_n 0.0146057f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_436 N_A_500_392#_c_347_n N_A_1224_74#_c_1279_n 0.00534955f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_437 N_A_500_392#_c_351_n N_A_1224_74#_c_1279_n 0.00761315f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_438 N_A_500_392#_c_347_n N_A_1224_74#_c_1280_n 4.21127e-19 $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_439 N_A_500_392#_c_339_n N_A_1224_74#_c_1280_n 0.0133634f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_440 N_A_500_392#_c_351_n N_A_1224_74#_c_1280_n 0.00832552f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_441 N_A_500_392#_c_347_n N_A_1224_74#_c_1281_n 0.005245f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_442 N_A_500_392#_c_339_n N_A_1224_74#_c_1281_n 0.00741853f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_443 N_A_500_392#_c_351_n N_A_1224_74#_c_1281_n 0.0242903f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_444 N_A_500_392#_c_347_n N_VPWR_c_1497_n 0.00349642f $X=7.25 $Y=2.28 $X2=0
+ $Y2=0
cc_445 N_A_500_392#_c_347_n N_VPWR_c_1482_n 0.00489211f $X=7.25 $Y=2.28 $X2=0
+ $Y2=0
cc_446 N_A_500_392#_c_348_n N_VPWR_c_1482_n 9.39239e-19 $X=3.462 $Y=2.21 $X2=0
+ $Y2=0
cc_447 N_A_500_392#_M1030_d N_A_38_78#_c_1648_n 0.00662817f $X=2.5 $Y=1.96 $X2=0
+ $Y2=0
cc_448 N_A_500_392#_c_349_n N_A_38_78#_c_1648_n 0.0274349f $X=2.915 $Y=2.052
+ $X2=0 $Y2=0
cc_449 N_A_500_392#_c_341_n N_A_38_78#_c_1648_n 0.00674361f $X=3.385 $Y=1.82
+ $X2=0 $Y2=0
cc_450 N_A_500_392#_c_334_n N_A_38_78#_c_1639_n 0.0166799f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_451 N_A_500_392#_c_340_n N_A_38_78#_c_1639_n 0.0174324f $X=2.862 $Y=0.34
+ $X2=0 $Y2=0
cc_452 N_A_500_392#_c_332_n N_A_38_78#_c_1640_n 3.38135e-19 $X=4.05 $Y=1.24
+ $X2=0 $Y2=0
cc_453 N_A_500_392#_c_342_n N_A_38_78#_c_1640_n 0.0106596f $X=3.052 $Y=1.205
+ $X2=0 $Y2=0
cc_454 N_A_500_392#_c_326_n N_A_38_78#_c_1649_n 0.0029567f $X=3.94 $Y=1.635
+ $X2=0 $Y2=0
cc_455 N_A_500_392#_c_348_n N_A_38_78#_c_1649_n 0.0147646f $X=3.462 $Y=2.21
+ $X2=0 $Y2=0
cc_456 N_A_500_392#_c_341_n N_A_38_78#_c_1649_n 0.00941428f $X=3.385 $Y=1.82
+ $X2=0 $Y2=0
cc_457 N_A_500_392#_c_325_n N_A_38_78#_c_1641_n 0.010222f $X=3.462 $Y=1.985
+ $X2=0 $Y2=0
cc_458 N_A_500_392#_c_326_n N_A_38_78#_c_1641_n 0.0133559f $X=3.94 $Y=1.635
+ $X2=0 $Y2=0
cc_459 N_A_500_392#_c_327_n N_A_38_78#_c_1641_n 0.00392644f $X=4.015 $Y=1.56
+ $X2=0 $Y2=0
cc_460 N_A_500_392#_c_341_n N_A_38_78#_c_1641_n 0.034635f $X=3.385 $Y=1.82 $X2=0
+ $Y2=0
cc_461 N_A_500_392#_c_343_n N_A_38_78#_c_1641_n 0.00717504f $X=3.052 $Y=1.39
+ $X2=0 $Y2=0
cc_462 N_A_500_392#_c_325_n N_A_38_78#_c_1653_n 8.82726e-19 $X=3.462 $Y=1.985
+ $X2=0 $Y2=0
cc_463 N_A_500_392#_c_341_n N_A_38_78#_c_1653_n 0.0214811f $X=3.385 $Y=1.82
+ $X2=0 $Y2=0
cc_464 N_A_500_392#_c_341_n N_A_38_78#_c_1643_n 0.00170906f $X=3.385 $Y=1.82
+ $X2=0 $Y2=0
cc_465 N_A_500_392#_c_342_n N_A_38_78#_c_1643_n 0.0174324f $X=3.052 $Y=1.205
+ $X2=0 $Y2=0
cc_466 N_A_500_392#_c_325_n N_A_38_78#_c_1644_n 0.00452157f $X=3.462 $Y=1.985
+ $X2=0 $Y2=0
cc_467 N_A_500_392#_c_326_n N_A_38_78#_c_1644_n 7.83113e-19 $X=3.94 $Y=1.635
+ $X2=0 $Y2=0
cc_468 N_A_500_392#_c_332_n N_A_38_78#_c_1644_n 0.00147521f $X=4.05 $Y=1.24
+ $X2=0 $Y2=0
cc_469 N_A_500_392#_c_341_n N_A_38_78#_c_1644_n 0.0109562f $X=3.385 $Y=1.82
+ $X2=0 $Y2=0
cc_470 N_A_500_392#_c_343_n N_A_38_78#_c_1644_n 0.0125584f $X=3.052 $Y=1.39
+ $X2=0 $Y2=0
cc_471 N_A_500_392#_c_336_n N_VGND_M1015_d 0.00722747f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_472 N_A_500_392#_c_340_n N_VGND_c_1819_n 0.0339415f $X=2.862 $Y=0.34 $X2=0
+ $Y2=0
cc_473 N_A_500_392#_c_334_n N_VGND_c_1824_n 0.0908278f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_474 N_A_500_392#_c_336_n N_VGND_c_1824_n 0.00941435f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_475 N_A_500_392#_c_340_n N_VGND_c_1824_n 0.0339438f $X=2.862 $Y=0.34 $X2=0
+ $Y2=0
cc_476 N_A_500_392#_c_328_n N_VGND_c_1825_n 0.00320103f $X=6.045 $Y=1.085 $X2=0
+ $Y2=0
cc_477 N_A_500_392#_c_336_n N_VGND_c_1825_n 0.0163564f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_478 N_A_500_392#_c_328_n N_VGND_c_1829_n 0.00407044f $X=6.045 $Y=1.085 $X2=0
+ $Y2=0
cc_479 N_A_500_392#_c_334_n N_VGND_c_1829_n 0.0472862f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_480 N_A_500_392#_c_336_n N_VGND_c_1829_n 0.0405193f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_481 N_A_500_392#_c_340_n N_VGND_c_1829_n 0.0171833f $X=2.862 $Y=0.34 $X2=0
+ $Y2=0
cc_482 N_A_500_392#_c_334_n N_VGND_c_1832_n 0.00667783f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_483 N_A_500_392#_c_336_n N_VGND_c_1832_n 0.0245264f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_484 N_A_500_392#_c_336_n A_910_119# 0.00134207f $X=6.085 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_485 N_A_841_401#_M1033_g N_RESET_B_c_643_n 0.00973011f $X=4.475 $Y=0.805
+ $X2=0 $Y2=0
cc_486 N_A_841_401#_M1033_g N_RESET_B_M1015_g 0.0415966f $X=4.475 $Y=0.805 $X2=0
+ $Y2=0
cc_487 N_A_841_401#_c_533_n N_RESET_B_M1015_g 0.0140148f $X=5.745 $Y=1.005 $X2=0
+ $Y2=0
cc_488 N_A_841_401#_M1033_g N_RESET_B_c_646_n 0.00952315f $X=4.475 $Y=0.805
+ $X2=0 $Y2=0
cc_489 N_A_841_401#_c_531_n N_RESET_B_c_646_n 0.00524003f $X=4.465 $Y=1.65 $X2=0
+ $Y2=0
cc_490 N_A_841_401#_c_532_n N_RESET_B_c_646_n 0.0210965f $X=4.465 $Y=1.65 $X2=0
+ $Y2=0
cc_491 N_A_841_401#_c_539_n N_RESET_B_c_655_n 0.0118146f $X=4.295 $Y=2.24 $X2=0
+ $Y2=0
cc_492 N_A_841_401#_c_531_n N_RESET_B_c_648_n 0.00340449f $X=4.465 $Y=1.65 $X2=0
+ $Y2=0
cc_493 N_A_841_401#_c_533_n N_RESET_B_c_648_n 0.00175352f $X=5.745 $Y=1.005
+ $X2=0 $Y2=0
cc_494 N_A_841_401#_c_540_n N_RESET_B_c_658_n 0.0230883f $X=4.465 $Y=2.005 $X2=0
+ $Y2=0
cc_495 N_A_841_401#_c_540_n N_RESET_B_c_659_n 0.00655097f $X=4.465 $Y=2.005
+ $X2=0 $Y2=0
cc_496 N_A_841_401#_c_531_n N_RESET_B_c_659_n 0.0255411f $X=4.465 $Y=1.65 $X2=0
+ $Y2=0
cc_497 N_A_841_401#_M1017_d N_RESET_B_c_661_n 0.00313731f $X=6.165 $Y=1.735
+ $X2=0 $Y2=0
cc_498 N_A_841_401#_c_537_n N_RESET_B_c_661_n 0.0067544f $X=6.23 $Y=1.485 $X2=0
+ $Y2=0
cc_499 N_A_841_401#_c_538_n N_RESET_B_c_661_n 0.00201833f $X=5.915 $Y=1.485
+ $X2=0 $Y2=0
cc_500 N_A_841_401#_c_544_n N_RESET_B_c_661_n 0.0328549f $X=6.315 $Y=1.88 $X2=0
+ $Y2=0
cc_501 N_A_841_401#_c_533_n N_A_705_463#_M1002_g 0.011848f $X=5.745 $Y=1.005
+ $X2=0 $Y2=0
cc_502 N_A_841_401#_c_536_n N_A_705_463#_M1002_g 0.0046522f $X=5.83 $Y=1.4 $X2=0
+ $Y2=0
cc_503 N_A_841_401#_c_533_n N_A_705_463#_c_854_n 0.00506798f $X=5.745 $Y=1.005
+ $X2=0 $Y2=0
cc_504 N_A_841_401#_c_537_n N_A_705_463#_c_854_n 0.00925955f $X=6.23 $Y=1.485
+ $X2=0 $Y2=0
cc_505 N_A_841_401#_c_538_n N_A_705_463#_c_854_n 0.00867517f $X=5.915 $Y=1.485
+ $X2=0 $Y2=0
cc_506 N_A_841_401#_c_544_n N_A_705_463#_c_854_n 0.00185802f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_507 N_A_841_401#_c_544_n N_A_705_463#_c_860_n 0.00551932f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_508 N_A_841_401#_c_539_n N_A_705_463#_c_887_n 0.00751864f $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_509 N_A_841_401#_c_540_n N_A_705_463#_c_887_n 0.00160627f $X=4.465 $Y=2.005
+ $X2=0 $Y2=0
cc_510 N_A_841_401#_c_531_n N_A_705_463#_c_887_n 0.0183792f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_511 N_A_841_401#_c_540_n N_A_705_463#_c_861_n 4.44352e-19 $X=4.465 $Y=2.005
+ $X2=0 $Y2=0
cc_512 N_A_841_401#_c_531_n N_A_705_463#_c_861_n 0.025646f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_513 N_A_841_401#_c_532_n N_A_705_463#_c_861_n 0.00174091f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_514 N_A_841_401#_c_534_n N_A_705_463#_c_855_n 0.00118569f $X=4.63 $Y=1.005
+ $X2=0 $Y2=0
cc_515 N_A_841_401#_c_539_n N_A_705_463#_c_894_n 0.00995576f $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_516 N_A_841_401#_c_539_n N_A_705_463#_c_856_n 0.00179692f $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_517 N_A_841_401#_M1033_g N_A_705_463#_c_856_n 0.00126786f $X=4.475 $Y=0.805
+ $X2=0 $Y2=0
cc_518 N_A_841_401#_c_540_n N_A_705_463#_c_856_n 0.00408065f $X=4.465 $Y=2.005
+ $X2=0 $Y2=0
cc_519 N_A_841_401#_c_531_n N_A_705_463#_c_856_n 0.0796661f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_520 N_A_841_401#_c_532_n N_A_705_463#_c_856_n 0.00808319f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_521 N_A_841_401#_c_534_n N_A_705_463#_c_856_n 0.0050659f $X=4.63 $Y=1.005
+ $X2=0 $Y2=0
cc_522 N_A_841_401#_c_531_n N_A_705_463#_c_857_n 0.0144822f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_523 N_A_841_401#_c_532_n N_A_705_463#_c_857_n 4.19328e-19 $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_524 N_A_841_401#_c_533_n N_A_705_463#_c_857_n 0.0375552f $X=5.745 $Y=1.005
+ $X2=0 $Y2=0
cc_525 N_A_841_401#_c_536_n N_A_705_463#_c_857_n 0.00811118f $X=5.83 $Y=1.4
+ $X2=0 $Y2=0
cc_526 N_A_841_401#_c_538_n N_A_705_463#_c_857_n 0.0135374f $X=5.915 $Y=1.485
+ $X2=0 $Y2=0
cc_527 N_A_841_401#_c_544_n N_A_705_463#_c_857_n 0.0012591f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_528 N_A_841_401#_c_533_n N_A_705_463#_c_858_n 0.00123201f $X=5.745 $Y=1.005
+ $X2=0 $Y2=0
cc_529 N_A_841_401#_c_536_n N_A_705_463#_c_858_n 7.93674e-19 $X=5.83 $Y=1.4
+ $X2=0 $Y2=0
cc_530 N_A_841_401#_c_538_n N_A_705_463#_c_858_n 5.0886e-19 $X=5.915 $Y=1.485
+ $X2=0 $Y2=0
cc_531 N_A_841_401#_c_539_n N_A_705_463#_c_864_n 9.24612e-19 $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_532 N_A_841_401#_c_539_n N_A_319_392#_c_996_n 0.00323347f $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_533 N_A_841_401#_c_539_n N_A_319_392#_c_998_n 0.0289372f $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_534 N_A_841_401#_c_540_n N_A_319_392#_c_998_n 0.0026362f $X=4.465 $Y=2.005
+ $X2=0 $Y2=0
cc_535 N_A_841_401#_c_539_n N_A_319_392#_c_999_n 0.00996184f $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_536 N_A_841_401#_c_544_n N_A_319_392#_c_999_n 0.00262042f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_537 N_A_841_401#_c_544_n N_A_319_392#_c_1000_n 5.08057e-19 $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_538 N_A_841_401#_c_544_n N_A_319_392#_M1012_g 0.0143858f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_539 N_A_841_401#_c_537_n N_A_319_392#_c_986_n 0.00287849f $X=6.23 $Y=1.485
+ $X2=0 $Y2=0
cc_540 N_A_841_401#_c_544_n N_A_319_392#_c_986_n 0.00245265f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_541 N_A_841_401#_c_544_n N_A_1224_74#_c_1301_n 0.0217845f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_542 N_A_841_401#_c_539_n N_VPWR_c_1487_n 0.00526245f $X=4.295 $Y=2.24 $X2=0
+ $Y2=0
cc_543 N_A_841_401#_c_537_n N_VPWR_c_1488_n 0.00590731f $X=6.23 $Y=1.485 $X2=0
+ $Y2=0
cc_544 N_A_841_401#_c_538_n N_VPWR_c_1488_n 0.0111121f $X=5.915 $Y=1.485 $X2=0
+ $Y2=0
cc_545 N_A_841_401#_c_544_n N_VPWR_c_1488_n 0.0651453f $X=6.315 $Y=1.88 $X2=0
+ $Y2=0
cc_546 N_A_841_401#_c_544_n N_VPWR_c_1497_n 0.00567879f $X=6.315 $Y=1.88 $X2=0
+ $Y2=0
cc_547 N_A_841_401#_c_539_n N_VPWR_c_1482_n 9.39239e-19 $X=4.295 $Y=2.24 $X2=0
+ $Y2=0
cc_548 N_A_841_401#_c_544_n N_VPWR_c_1482_n 0.00684413f $X=6.315 $Y=1.88 $X2=0
+ $Y2=0
cc_549 N_A_841_401#_c_533_n N_VGND_M1015_d 0.00389013f $X=5.745 $Y=1.005 $X2=0
+ $Y2=0
cc_550 N_A_841_401#_c_533_n A_910_119# 0.00103428f $X=5.745 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_551 N_A_841_401#_c_534_n A_910_119# 2.36857e-19 $X=4.63 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_552 N_RESET_B_c_643_n N_A_705_463#_M1002_g 0.0226708f $X=4.79 $Y=0.18 $X2=0
+ $Y2=0
cc_553 N_RESET_B_c_648_n N_A_705_463#_M1002_g 0.00742734f $X=4.89 $Y=1.24 $X2=0
+ $Y2=0
cc_554 N_RESET_B_c_661_n N_A_705_463#_c_854_n 0.00249739f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_555 N_RESET_B_c_662_n N_A_705_463#_c_854_n 0.00116431f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_556 N_RESET_B_c_665_n N_A_705_463#_c_854_n 0.0017604f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_557 N_RESET_B_c_661_n N_A_705_463#_c_860_n 0.0069988f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_558 N_RESET_B_c_659_n N_A_705_463#_c_870_n 0.00660896f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_559 N_RESET_B_c_655_n N_A_705_463#_c_887_n 0.00433773f $X=4.93 $Y=2.24 $X2=0
+ $Y2=0
cc_560 N_RESET_B_c_659_n N_A_705_463#_c_887_n 0.0157057f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_561 N_RESET_B_c_646_n N_A_705_463#_c_861_n 0.00671367f $X=4.915 $Y=1.825
+ $X2=0 $Y2=0
cc_562 N_RESET_B_c_655_n N_A_705_463#_c_861_n 0.0015898f $X=4.93 $Y=2.24 $X2=0
+ $Y2=0
cc_563 N_RESET_B_c_658_n N_A_705_463#_c_861_n 0.0106103f $X=4.93 $Y=2.032 $X2=0
+ $Y2=0
cc_564 N_RESET_B_c_659_n N_A_705_463#_c_861_n 0.0225339f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_565 N_RESET_B_c_662_n N_A_705_463#_c_861_n 4.39853e-19 $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_566 N_RESET_B_c_664_n N_A_705_463#_c_861_n 0.00639141f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_567 N_RESET_B_c_665_n N_A_705_463#_c_861_n 0.0224281f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_568 N_RESET_B_c_655_n N_A_705_463#_c_894_n 8.10749e-19 $X=4.93 $Y=2.24 $X2=0
+ $Y2=0
cc_569 N_RESET_B_c_659_n N_A_705_463#_c_894_n 0.00372169f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_570 N_RESET_B_c_659_n N_A_705_463#_c_856_n 0.0212929f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_571 N_RESET_B_c_646_n N_A_705_463#_c_857_n 0.00724972f $X=4.915 $Y=1.825
+ $X2=0 $Y2=0
cc_572 N_RESET_B_c_659_n N_A_705_463#_c_857_n 0.00610322f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_573 N_RESET_B_c_662_n N_A_705_463#_c_857_n 0.00107679f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_574 N_RESET_B_c_664_n N_A_705_463#_c_857_n 0.00682898f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_575 N_RESET_B_c_665_n N_A_705_463#_c_857_n 0.0190365f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_576 N_RESET_B_c_646_n N_A_705_463#_c_858_n 0.0174208f $X=4.915 $Y=1.825 $X2=0
+ $Y2=0
cc_577 N_RESET_B_c_664_n N_A_705_463#_c_858_n 0.0207972f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_578 N_RESET_B_c_665_n N_A_705_463#_c_858_n 4.14991e-19 $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_579 N_RESET_B_c_655_n N_A_705_463#_c_864_n 0.00883696f $X=4.93 $Y=2.24 $X2=0
+ $Y2=0
cc_580 N_RESET_B_c_659_n N_A_705_463#_c_864_n 0.00739764f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_581 N_RESET_B_c_664_n N_A_705_463#_c_864_n 0.00865293f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_582 N_RESET_B_c_665_n N_A_705_463#_c_864_n 0.00685251f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_583 N_RESET_B_c_659_n N_A_319_392#_M1000_s 0.00116894f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_584 N_RESET_B_c_659_n N_A_319_392#_M1030_g 0.00632197f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_585 N_RESET_B_c_643_n N_A_319_392#_c_981_n 0.0103526f $X=4.79 $Y=0.18 $X2=0
+ $Y2=0
cc_586 N_RESET_B_c_659_n N_A_319_392#_c_992_n 6.78785e-19 $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_587 N_RESET_B_c_643_n N_A_319_392#_M1013_g 0.00882199f $X=4.79 $Y=0.18 $X2=0
+ $Y2=0
cc_588 N_RESET_B_c_659_n N_A_319_392#_c_998_n 0.00242159f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_589 N_RESET_B_c_655_n N_A_319_392#_c_999_n 0.010005f $X=4.93 $Y=2.24 $X2=0
+ $Y2=0
cc_590 N_RESET_B_c_661_n N_A_319_392#_M1012_g 0.0118743f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_591 N_RESET_B_c_661_n N_A_319_392#_c_985_n 3.83564e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_592 N_RESET_B_c_661_n N_A_319_392#_c_986_n 3.03408e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_593 N_RESET_B_c_649_n N_A_319_392#_c_988_n 0.00720421f $X=1.165 $Y=1.295
+ $X2=0 $Y2=0
cc_594 N_RESET_B_c_650_n N_A_319_392#_c_988_n 0.0535888f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_595 N_RESET_B_c_659_n N_A_319_392#_c_989_n 0.00305281f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_596 N_RESET_B_M1028_g N_A_319_392#_c_990_n 0.00414858f $X=0.94 $Y=0.6 $X2=0
+ $Y2=0
cc_597 N_RESET_B_c_643_n N_A_319_392#_c_990_n 0.00809322f $X=4.79 $Y=0.18 $X2=0
+ $Y2=0
cc_598 N_RESET_B_c_650_n N_A_319_392#_c_990_n 7.48694e-19 $X=1.165 $Y=1.295
+ $X2=0 $Y2=0
cc_599 N_RESET_B_c_642_n N_A_319_392#_c_1007_n 0.0024157f $X=1.097 $Y=1.908
+ $X2=0 $Y2=0
cc_600 N_RESET_B_c_652_n N_A_319_392#_c_1007_n 0.00267262f $X=0.955 $Y=2.375
+ $X2=0 $Y2=0
cc_601 N_RESET_B_c_659_n N_A_319_392#_c_1007_n 0.0312063f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_602 N_RESET_B_c_660_n N_A_319_392#_c_1007_n 0.00291288f $X=1.345 $Y=2.035
+ $X2=0 $Y2=0
cc_603 N_RESET_B_c_650_n N_A_319_392#_c_1007_n 0.0192935f $X=1.165 $Y=1.295
+ $X2=0 $Y2=0
cc_604 N_RESET_B_M1026_g N_A_1482_48#_c_1173_n 0.0196155f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_605 N_RESET_B_c_657_n N_A_1482_48#_c_1174_n 0.044692f $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_606 N_RESET_B_c_661_n N_A_1482_48#_c_1174_n 0.00564012f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_607 N_RESET_B_c_663_n N_A_1482_48#_c_1174_n 0.00149248f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_608 N_RESET_B_c_668_n N_A_1482_48#_c_1174_n 0.00190186f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_609 N_RESET_B_c_657_n N_A_1482_48#_c_1182_n 0.00623945f $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_610 N_RESET_B_M1026_g N_A_1482_48#_c_1175_n 0.0144302f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_611 N_RESET_B_c_657_n N_A_1482_48#_c_1183_n 0.00528461f $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_612 N_RESET_B_c_663_n N_A_1482_48#_c_1183_n 9.35982e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_613 N_RESET_B_c_668_n N_A_1482_48#_c_1183_n 0.0201792f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_614 N_RESET_B_M1026_g N_A_1482_48#_c_1176_n 0.00201284f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_615 N_RESET_B_M1026_g N_A_1482_48#_c_1178_n 0.00118187f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_616 N_RESET_B_M1026_g N_A_1482_48#_c_1185_n 0.00150115f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_617 N_RESET_B_c_657_n N_A_1482_48#_c_1185_n 3.55688e-19 $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_618 N_RESET_B_c_668_n N_A_1482_48#_c_1185_n 0.00823641f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_619 N_RESET_B_M1026_g N_A_1482_48#_c_1180_n 0.0401889f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_620 N_RESET_B_c_661_n N_A_1224_74#_M1012_d 0.00185339f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_621 N_RESET_B_M1026_g N_A_1224_74#_M1027_g 0.0533792f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_622 N_RESET_B_M1026_g N_A_1224_74#_c_1269_n 0.00701487f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_623 N_RESET_B_c_657_n N_A_1224_74#_c_1269_n 0.0230744f $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_624 N_RESET_B_c_668_n N_A_1224_74#_c_1269_n 3.64033e-19 $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_625 N_RESET_B_c_657_n N_A_1224_74#_c_1286_n 0.00895543f $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_626 N_RESET_B_M1026_g N_A_1224_74#_c_1271_n 0.0220605f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_627 N_RESET_B_c_661_n N_A_1224_74#_c_1301_n 0.0113671f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_628 N_RESET_B_c_661_n N_A_1224_74#_c_1279_n 0.00715094f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_629 N_RESET_B_c_661_n N_A_1224_74#_c_1280_n 0.00106639f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_630 N_RESET_B_M1026_g N_A_1224_74#_c_1281_n 0.00129569f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_631 N_RESET_B_c_657_n N_A_1224_74#_c_1281_n 0.00121033f $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_632 N_RESET_B_c_661_n N_A_1224_74#_c_1281_n 0.0226223f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_633 N_RESET_B_c_663_n N_A_1224_74#_c_1281_n 0.00270727f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_634 N_RESET_B_c_668_n N_A_1224_74#_c_1281_n 0.0230781f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_635 N_RESET_B_M1026_g N_A_1224_74#_c_1282_n 0.0108822f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_636 N_RESET_B_c_657_n N_A_1224_74#_c_1282_n 0.00436274f $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_637 N_RESET_B_c_661_n N_A_1224_74#_c_1282_n 0.00339956f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_638 N_RESET_B_c_663_n N_A_1224_74#_c_1282_n 0.00379913f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_639 N_RESET_B_c_668_n N_A_1224_74#_c_1282_n 0.0255102f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_640 N_RESET_B_M1026_g N_A_1224_74#_c_1284_n 0.00118353f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_641 N_RESET_B_c_659_n N_VPWR_M1000_d 0.00761697f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_642 N_RESET_B_c_661_n N_VPWR_M1017_s 0.00310864f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_643 N_RESET_B_c_653_n N_VPWR_c_1485_n 0.00732028f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_644 N_RESET_B_c_655_n N_VPWR_c_1487_n 0.00556482f $X=4.93 $Y=2.24 $X2=0 $Y2=0
cc_645 N_RESET_B_c_661_n N_VPWR_c_1488_n 0.0237051f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_646 N_RESET_B_c_662_n N_VPWR_c_1488_n 0.00275995f $X=5.665 $Y=2.035 $X2=0
+ $Y2=0
cc_647 N_RESET_B_c_664_n N_VPWR_c_1488_n 0.00101439f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_648 N_RESET_B_c_665_n N_VPWR_c_1488_n 0.0239958f $X=5.395 $Y=1.99 $X2=0 $Y2=0
cc_649 N_RESET_B_c_657_n N_VPWR_c_1489_n 0.0062044f $X=8.18 $Y=2.28 $X2=0 $Y2=0
cc_650 N_RESET_B_c_663_n N_VPWR_c_1489_n 0.00183431f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_651 N_RESET_B_c_668_n N_VPWR_c_1489_n 0.0174647f $X=8.135 $Y=2 $X2=0 $Y2=0
cc_652 N_RESET_B_c_657_n N_VPWR_c_1490_n 0.00454183f $X=8.18 $Y=2.28 $X2=0 $Y2=0
cc_653 N_RESET_B_c_653_n N_VPWR_c_1493_n 0.00303336f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_654 N_RESET_B_c_653_n N_VPWR_c_1482_n 0.0039334f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_655 N_RESET_B_c_655_n N_VPWR_c_1482_n 9.39239e-19 $X=4.93 $Y=2.24 $X2=0 $Y2=0
cc_656 N_RESET_B_c_657_n N_VPWR_c_1482_n 0.00489211f $X=8.18 $Y=2.28 $X2=0 $Y2=0
cc_657 N_RESET_B_M1028_g N_A_38_78#_c_1637_n 7.65322e-19 $X=0.94 $Y=0.6 $X2=0
+ $Y2=0
cc_658 N_RESET_B_c_653_n N_A_38_78#_c_1645_n 2.24915e-19 $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_659 N_RESET_B_M1028_g N_A_38_78#_c_1638_n 0.0167617f $X=0.94 $Y=0.6 $X2=0
+ $Y2=0
cc_660 N_RESET_B_c_660_n N_A_38_78#_c_1638_n 0.00199354f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_661 N_RESET_B_c_650_n N_A_38_78#_c_1638_n 0.0731888f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_662 N_RESET_B_c_652_n N_A_38_78#_c_1647_n 0.00897965f $X=0.955 $Y=2.375 $X2=0
+ $Y2=0
cc_663 N_RESET_B_c_653_n N_A_38_78#_c_1647_n 0.0112966f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_664 N_RESET_B_c_659_n N_A_38_78#_c_1647_n 0.0058487f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_665 N_RESET_B_c_660_n N_A_38_78#_c_1647_n 0.00916403f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_666 N_RESET_B_c_650_n N_A_38_78#_c_1647_n 0.0179915f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_667 N_RESET_B_c_667_n N_A_38_78#_c_1647_n 0.00293275f $X=1.165 $Y=1.975 $X2=0
+ $Y2=0
cc_668 N_RESET_B_c_659_n N_A_38_78#_c_1648_n 0.00472935f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_669 N_RESET_B_c_659_n N_A_38_78#_c_1649_n 0.0118525f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_670 N_RESET_B_c_659_n N_A_38_78#_c_1641_n 0.0132834f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_671 N_RESET_B_M1028_g N_A_38_78#_c_1642_n 8.39005e-19 $X=0.94 $Y=0.6 $X2=0
+ $Y2=0
cc_672 N_RESET_B_c_652_n N_A_38_78#_c_1651_n 0.00180915f $X=0.955 $Y=2.375 $X2=0
+ $Y2=0
cc_673 N_RESET_B_c_653_n N_A_38_78#_c_1651_n 0.00426947f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_674 N_RESET_B_c_659_n N_A_38_78#_c_1652_n 0.00420888f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_675 N_RESET_B_c_659_n N_A_38_78#_c_1669_n 0.0182491f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_676 N_RESET_B_c_659_n N_A_38_78#_c_1653_n 0.00774538f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_677 N_RESET_B_c_659_n N_A_38_78#_c_1644_n 0.00599017f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_678 N_RESET_B_M1028_g N_VGND_c_1817_n 0.00269179f $X=0.94 $Y=0.6 $X2=0 $Y2=0
cc_679 N_RESET_B_c_643_n N_VGND_c_1817_n 0.0190483f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_680 N_RESET_B_c_649_n N_VGND_c_1817_n 0.00181416f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_681 N_RESET_B_c_650_n N_VGND_c_1817_n 0.0144384f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_682 N_RESET_B_c_643_n N_VGND_c_1818_n 0.0235672f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_683 N_RESET_B_c_643_n N_VGND_c_1819_n 0.0257653f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_684 N_RESET_B_M1026_g N_VGND_c_1820_n 0.0152783f $X=8.045 $Y=0.58 $X2=0 $Y2=0
cc_685 N_RESET_B_c_644_n N_VGND_c_1823_n 0.0064002f $X=1.015 $Y=0.18 $X2=0 $Y2=0
cc_686 N_RESET_B_c_643_n N_VGND_c_1824_n 0.0561385f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_687 N_RESET_B_M1026_g N_VGND_c_1826_n 0.00383152f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_688 N_RESET_B_c_643_n N_VGND_c_1829_n 0.0943075f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_689 N_RESET_B_c_644_n N_VGND_c_1829_n 0.0113744f $X=1.015 $Y=0.18 $X2=0 $Y2=0
cc_690 N_RESET_B_M1026_g N_VGND_c_1829_n 0.0075725f $X=8.045 $Y=0.58 $X2=0 $Y2=0
cc_691 N_RESET_B_c_643_n N_VGND_c_1832_n 0.00776078f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_692 N_A_705_463#_c_870_n N_A_319_392#_c_993_n 0.00333009f $X=4.01 $Y=2.61
+ $X2=0 $Y2=0
cc_693 N_A_705_463#_c_855_n N_A_319_392#_M1013_g 0.00230849f $X=4.095 $Y=0.812
+ $X2=0 $Y2=0
cc_694 N_A_705_463#_c_856_n N_A_319_392#_M1013_g 5.83463e-19 $X=4.14 $Y=2.325
+ $X2=0 $Y2=0
cc_695 N_A_705_463#_c_870_n N_A_319_392#_c_998_n 0.00897602f $X=4.01 $Y=2.61
+ $X2=0 $Y2=0
cc_696 N_A_705_463#_c_856_n N_A_319_392#_c_998_n 0.00168289f $X=4.14 $Y=2.325
+ $X2=0 $Y2=0
cc_697 N_A_705_463#_c_860_n N_A_319_392#_c_999_n 0.0103562f $X=6.09 $Y=1.66
+ $X2=0 $Y2=0
cc_698 N_A_705_463#_c_887_n N_A_319_392#_c_999_n 0.00337238f $X=4.89 $Y=2.41
+ $X2=0 $Y2=0
cc_699 N_A_705_463#_c_894_n N_A_319_392#_c_999_n 0.00241116f $X=4.14 $Y=2.41
+ $X2=0 $Y2=0
cc_700 N_A_705_463#_c_864_n N_A_319_392#_c_999_n 0.0059408f $X=4.975 $Y=2.48
+ $X2=0 $Y2=0
cc_701 N_A_705_463#_c_860_n N_A_319_392#_c_1000_n 0.00249951f $X=6.09 $Y=1.66
+ $X2=0 $Y2=0
cc_702 N_A_705_463#_c_860_n N_A_319_392#_M1012_g 0.00575058f $X=6.09 $Y=1.66
+ $X2=0 $Y2=0
cc_703 N_A_705_463#_c_854_n N_A_319_392#_c_986_n 0.00860655f $X=6 $Y=1.54 $X2=0
+ $Y2=0
cc_704 N_A_705_463#_c_887_n N_VPWR_M1006_d 0.0084725f $X=4.89 $Y=2.41 $X2=0
+ $Y2=0
cc_705 N_A_705_463#_c_887_n N_VPWR_c_1487_n 0.0264204f $X=4.89 $Y=2.41 $X2=0
+ $Y2=0
cc_706 N_A_705_463#_c_894_n N_VPWR_c_1487_n 0.00229636f $X=4.14 $Y=2.41 $X2=0
+ $Y2=0
cc_707 N_A_705_463#_c_864_n N_VPWR_c_1487_n 0.00101701f $X=4.975 $Y=2.48 $X2=0
+ $Y2=0
cc_708 N_A_705_463#_c_854_n N_VPWR_c_1488_n 0.00446017f $X=6 $Y=1.54 $X2=0 $Y2=0
cc_709 N_A_705_463#_c_860_n N_VPWR_c_1488_n 0.0144868f $X=6.09 $Y=1.66 $X2=0
+ $Y2=0
cc_710 N_A_705_463#_c_864_n N_VPWR_c_1488_n 0.0158268f $X=4.975 $Y=2.48 $X2=0
+ $Y2=0
cc_711 N_A_705_463#_c_870_n N_VPWR_c_1495_n 0.0073432f $X=4.01 $Y=2.61 $X2=0
+ $Y2=0
cc_712 N_A_705_463#_c_894_n N_VPWR_c_1495_n 0.00408501f $X=4.14 $Y=2.41 $X2=0
+ $Y2=0
cc_713 N_A_705_463#_c_864_n N_VPWR_c_1496_n 0.00551323f $X=4.975 $Y=2.48 $X2=0
+ $Y2=0
cc_714 N_A_705_463#_c_860_n N_VPWR_c_1482_n 8.51577e-19 $X=6.09 $Y=1.66 $X2=0
+ $Y2=0
cc_715 N_A_705_463#_c_870_n N_VPWR_c_1482_n 0.0119615f $X=4.01 $Y=2.61 $X2=0
+ $Y2=0
cc_716 N_A_705_463#_c_887_n N_VPWR_c_1482_n 0.00920255f $X=4.89 $Y=2.41 $X2=0
+ $Y2=0
cc_717 N_A_705_463#_c_894_n N_VPWR_c_1482_n 0.00667121f $X=4.14 $Y=2.41 $X2=0
+ $Y2=0
cc_718 N_A_705_463#_c_864_n N_VPWR_c_1482_n 0.0117253f $X=4.975 $Y=2.48 $X2=0
+ $Y2=0
cc_719 N_A_705_463#_c_855_n N_A_38_78#_c_1639_n 0.0161825f $X=4.095 $Y=0.812
+ $X2=0 $Y2=0
cc_720 N_A_705_463#_M1023_d N_A_38_78#_c_1649_n 0.00206971f $X=3.525 $Y=2.315
+ $X2=0 $Y2=0
cc_721 N_A_705_463#_c_870_n N_A_38_78#_c_1649_n 0.0154028f $X=4.01 $Y=2.61 $X2=0
+ $Y2=0
cc_722 N_A_705_463#_c_856_n N_A_38_78#_c_1649_n 0.0120586f $X=4.14 $Y=2.325
+ $X2=0 $Y2=0
cc_723 N_A_705_463#_c_856_n N_A_38_78#_c_1641_n 0.0587849f $X=4.14 $Y=2.325
+ $X2=0 $Y2=0
cc_724 N_A_705_463#_c_856_n N_A_38_78#_c_1643_n 0.00502811f $X=4.14 $Y=2.325
+ $X2=0 $Y2=0
cc_725 N_A_705_463#_c_855_n N_A_38_78#_c_1644_n 0.0109431f $X=4.095 $Y=0.812
+ $X2=0 $Y2=0
cc_726 N_A_705_463#_c_856_n N_A_38_78#_c_1644_n 0.0131878f $X=4.14 $Y=2.325
+ $X2=0 $Y2=0
cc_727 N_A_705_463#_c_894_n A_796_463# 0.00200517f $X=4.14 $Y=2.41 $X2=-0.19
+ $Y2=-0.245
cc_728 N_A_705_463#_M1002_g N_VGND_c_1825_n 0.00320129f $X=5.455 $Y=0.69 $X2=0
+ $Y2=0
cc_729 N_A_705_463#_M1002_g N_VGND_c_1829_n 0.00402508f $X=5.455 $Y=0.69 $X2=0
+ $Y2=0
cc_730 N_A_705_463#_M1002_g N_VGND_c_1832_n 0.00397703f $X=5.455 $Y=0.69 $X2=0
+ $Y2=0
cc_731 N_A_319_392#_M1032_g N_A_1482_48#_c_1173_n 0.0495982f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_732 N_A_319_392#_M1032_g N_A_1482_48#_c_1174_n 0.0112982f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_733 N_A_319_392#_M1032_g N_A_1482_48#_c_1178_n 0.00102678f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_734 N_A_319_392#_M1032_g N_A_1224_74#_c_1297_n 0.0169263f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_735 N_A_319_392#_M1012_g N_A_1224_74#_c_1301_n 0.00382767f $X=6.54 $Y=2.235
+ $X2=0 $Y2=0
cc_736 N_A_319_392#_M1032_g N_A_1224_74#_c_1278_n 0.0221333f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_737 N_A_319_392#_c_985_n N_A_1224_74#_c_1279_n 0.00206465f $X=7.02 $Y=1.55
+ $X2=0 $Y2=0
cc_738 N_A_319_392#_M1032_g N_A_1224_74#_c_1279_n 0.0011854f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_739 N_A_319_392#_c_985_n N_A_1224_74#_c_1280_n 0.00561544f $X=7.02 $Y=1.55
+ $X2=0 $Y2=0
cc_740 N_A_319_392#_M1032_g N_A_1224_74#_c_1280_n 0.00135722f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_741 N_A_319_392#_c_985_n N_A_1224_74#_c_1281_n 3.07924e-19 $X=7.02 $Y=1.55
+ $X2=0 $Y2=0
cc_742 N_A_319_392#_M1030_g N_VPWR_c_1486_n 0.00777078f $X=2.425 $Y=2.46 $X2=0
+ $Y2=0
cc_743 N_A_319_392#_c_992_n N_VPWR_c_1486_n 0.0015647f $X=2.935 $Y=3.075 $X2=0
+ $Y2=0
cc_744 N_A_319_392#_c_994_n N_VPWR_c_1486_n 0.00232909f $X=3.01 $Y=3.15 $X2=0
+ $Y2=0
cc_745 N_A_319_392#_c_996_n N_VPWR_c_1487_n 0.00604299f $X=3.905 $Y=2.9 $X2=0
+ $Y2=0
cc_746 N_A_319_392#_c_999_n N_VPWR_c_1487_n 0.0261571f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_747 N_A_319_392#_c_999_n N_VPWR_c_1488_n 0.0213056f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_748 N_A_319_392#_c_1000_n N_VPWR_c_1488_n 0.00613773f $X=6.54 $Y=2.9 $X2=0
+ $Y2=0
cc_749 N_A_319_392#_M1012_g N_VPWR_c_1488_n 6.32588e-19 $X=6.54 $Y=2.235 $X2=0
+ $Y2=0
cc_750 N_A_319_392#_M1030_g N_VPWR_c_1495_n 0.00326216f $X=2.425 $Y=2.46 $X2=0
+ $Y2=0
cc_751 N_A_319_392#_c_994_n N_VPWR_c_1495_n 0.0448843f $X=3.01 $Y=3.15 $X2=0
+ $Y2=0
cc_752 N_A_319_392#_c_999_n N_VPWR_c_1496_n 0.0315528f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_753 N_A_319_392#_c_999_n N_VPWR_c_1497_n 0.0193014f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_754 N_A_319_392#_M1030_g N_VPWR_c_1482_n 0.00423492f $X=2.425 $Y=2.46 $X2=0
+ $Y2=0
cc_755 N_A_319_392#_c_993_n N_VPWR_c_1482_n 0.0235991f $X=3.815 $Y=3.15 $X2=0
+ $Y2=0
cc_756 N_A_319_392#_c_994_n N_VPWR_c_1482_n 0.00688635f $X=3.01 $Y=3.15 $X2=0
+ $Y2=0
cc_757 N_A_319_392#_c_999_n N_VPWR_c_1482_n 0.0775234f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_758 N_A_319_392#_c_1005_n N_VPWR_c_1482_n 0.00512307f $X=3.905 $Y=3.15 $X2=0
+ $Y2=0
cc_759 N_A_319_392#_c_990_n N_A_38_78#_c_1638_n 0.0101177f $X=1.92 $Y=0.867
+ $X2=0 $Y2=0
cc_760 N_A_319_392#_c_1007_n N_A_38_78#_c_1647_n 0.00319492f $X=1.555 $Y=2.057
+ $X2=0 $Y2=0
cc_761 N_A_319_392#_M1030_g N_A_38_78#_c_1648_n 0.0131699f $X=2.425 $Y=2.46
+ $X2=0 $Y2=0
cc_762 N_A_319_392#_c_992_n N_A_38_78#_c_1648_n 0.0130681f $X=2.935 $Y=3.075
+ $X2=0 $Y2=0
cc_763 N_A_319_392#_M1013_g N_A_38_78#_c_1639_n 0.00375823f $X=3.585 $Y=0.805
+ $X2=0 $Y2=0
cc_764 N_A_319_392#_c_982_n N_A_38_78#_c_1640_n 0.00370387f $X=3.51 $Y=1.275
+ $X2=0 $Y2=0
cc_765 N_A_319_392#_M1013_g N_A_38_78#_c_1640_n 0.0056506f $X=3.585 $Y=0.805
+ $X2=0 $Y2=0
cc_766 N_A_319_392#_c_998_n N_A_38_78#_c_1649_n 0.00397085f $X=3.905 $Y=2.81
+ $X2=0 $Y2=0
cc_767 N_A_319_392#_c_983_n N_A_38_78#_c_1641_n 0.00102542f $X=3.145 $Y=1.275
+ $X2=0 $Y2=0
cc_768 N_A_319_392#_M1000_s N_A_38_78#_c_1652_n 0.00803591f $X=1.595 $Y=1.96
+ $X2=0 $Y2=0
cc_769 N_A_319_392#_c_1007_n N_A_38_78#_c_1652_n 0.0203078f $X=1.555 $Y=2.057
+ $X2=0 $Y2=0
cc_770 N_A_319_392#_c_992_n N_A_38_78#_c_1653_n 0.00810868f $X=2.935 $Y=3.075
+ $X2=0 $Y2=0
cc_771 N_A_319_392#_c_993_n N_A_38_78#_c_1653_n 0.00444409f $X=3.815 $Y=3.15
+ $X2=0 $Y2=0
cc_772 N_A_319_392#_c_982_n N_A_38_78#_c_1643_n 0.00108086f $X=3.51 $Y=1.275
+ $X2=0 $Y2=0
cc_773 N_A_319_392#_M1013_g N_A_38_78#_c_1643_n 0.00186734f $X=3.585 $Y=0.805
+ $X2=0 $Y2=0
cc_774 N_A_319_392#_c_982_n N_A_38_78#_c_1644_n 0.0151742f $X=3.51 $Y=1.275
+ $X2=0 $Y2=0
cc_775 N_A_319_392#_c_1018_n N_VGND_M1001_d 0.00948826f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_776 N_A_319_392#_c_990_n N_VGND_c_1817_n 0.0178351f $X=1.92 $Y=0.867 $X2=0
+ $Y2=0
cc_777 N_A_319_392#_c_990_n N_VGND_c_1818_n 0.0088414f $X=1.92 $Y=0.867 $X2=0
+ $Y2=0
cc_778 N_A_319_392#_c_981_n N_VGND_c_1819_n 0.00249513f $X=2.55 $Y=1.41 $X2=0
+ $Y2=0
cc_779 N_A_319_392#_c_1018_n N_VGND_c_1819_n 0.0257093f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_780 N_A_319_392#_M1032_g N_VGND_c_1820_n 0.00154981f $X=7.095 $Y=0.58 $X2=0
+ $Y2=0
cc_781 N_A_319_392#_M1032_g N_VGND_c_1825_n 0.00309049f $X=7.095 $Y=0.58 $X2=0
+ $Y2=0
cc_782 N_A_319_392#_c_981_n N_VGND_c_1829_n 8.51577e-19 $X=2.55 $Y=1.41 $X2=0
+ $Y2=0
cc_783 N_A_319_392#_M1032_g N_VGND_c_1829_n 0.0040628f $X=7.095 $Y=0.58 $X2=0
+ $Y2=0
cc_784 N_A_319_392#_c_990_n N_VGND_c_1829_n 0.0121021f $X=1.92 $Y=0.867 $X2=0
+ $Y2=0
cc_785 N_A_1482_48#_c_1175_n N_A_1224_74#_M1027_g 0.0108008f $X=8.485 $Y=0.985
+ $X2=0 $Y2=0
cc_786 N_A_1482_48#_c_1176_n N_A_1224_74#_M1027_g 0.0132755f $X=8.65 $Y=0.58
+ $X2=0 $Y2=0
cc_787 N_A_1482_48#_c_1177_n N_A_1224_74#_M1027_g 0.00584201f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_788 N_A_1482_48#_c_1179_n N_A_1224_74#_M1027_g 0.0045388f $X=8.727 $Y=0.985
+ $X2=0 $Y2=0
cc_789 N_A_1482_48#_c_1183_n N_A_1224_74#_c_1269_n 0.00705834f $X=8.555 $Y=2.335
+ $X2=0 $Y2=0
cc_790 N_A_1482_48#_c_1177_n N_A_1224_74#_c_1269_n 0.00407488f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_791 N_A_1482_48#_c_1185_n N_A_1224_74#_c_1269_n 0.0144908f $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_792 N_A_1482_48#_c_1183_n N_A_1224_74#_c_1286_n 0.0115505f $X=8.555 $Y=2.335
+ $X2=0 $Y2=0
cc_793 N_A_1482_48#_c_1177_n N_A_1224_74#_c_1270_n 0.0256662f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_794 N_A_1482_48#_c_1185_n N_A_1224_74#_c_1270_n 0.00384268f $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_795 N_A_1482_48#_c_1185_n N_A_1224_74#_c_1271_n 4.86873e-19 $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_796 N_A_1482_48#_c_1179_n N_A_1224_74#_c_1271_n 0.00795f $X=8.727 $Y=0.985
+ $X2=0 $Y2=0
cc_797 N_A_1482_48#_c_1183_n N_A_1224_74#_c_1272_n 5.60188e-19 $X=8.555 $Y=2.335
+ $X2=0 $Y2=0
cc_798 N_A_1482_48#_c_1177_n N_A_1224_74#_c_1272_n 0.00210772f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_799 N_A_1482_48#_c_1185_n N_A_1224_74#_c_1272_n 0.00185013f $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_800 N_A_1482_48#_c_1176_n N_A_1224_74#_M1009_g 0.00122775f $X=8.65 $Y=0.58
+ $X2=0 $Y2=0
cc_801 N_A_1482_48#_c_1177_n N_A_1224_74#_M1009_g 0.00251042f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_802 N_A_1482_48#_c_1173_n N_A_1224_74#_c_1297_n 0.0012657f $X=7.485 $Y=0.9
+ $X2=0 $Y2=0
cc_803 N_A_1482_48#_c_1182_n N_A_1224_74#_c_1301_n 0.00944193f $X=7.67 $Y=2.28
+ $X2=0 $Y2=0
cc_804 N_A_1482_48#_c_1173_n N_A_1224_74#_c_1278_n 0.00230939f $X=7.485 $Y=0.9
+ $X2=0 $Y2=0
cc_805 N_A_1482_48#_c_1174_n N_A_1224_74#_c_1278_n 0.00111943f $X=7.67 $Y=2.19
+ $X2=0 $Y2=0
cc_806 N_A_1482_48#_c_1178_n N_A_1224_74#_c_1278_n 0.0162835f $X=7.595 $Y=0.985
+ $X2=0 $Y2=0
cc_807 N_A_1482_48#_c_1178_n N_A_1224_74#_c_1279_n 0.00432309f $X=7.595 $Y=0.985
+ $X2=0 $Y2=0
cc_808 N_A_1482_48#_c_1180_n N_A_1224_74#_c_1279_n 0.00127859f $X=7.67 $Y=1.065
+ $X2=0 $Y2=0
cc_809 N_A_1482_48#_c_1174_n N_A_1224_74#_c_1281_n 0.0153989f $X=7.67 $Y=2.19
+ $X2=0 $Y2=0
cc_810 N_A_1482_48#_c_1182_n N_A_1224_74#_c_1281_n 0.00481867f $X=7.67 $Y=2.28
+ $X2=0 $Y2=0
cc_811 N_A_1482_48#_c_1174_n N_A_1224_74#_c_1282_n 0.00617973f $X=7.67 $Y=2.19
+ $X2=0 $Y2=0
cc_812 N_A_1482_48#_c_1175_n N_A_1224_74#_c_1282_n 0.0246405f $X=8.485 $Y=0.985
+ $X2=0 $Y2=0
cc_813 N_A_1482_48#_c_1178_n N_A_1224_74#_c_1282_n 0.00601156f $X=7.595 $Y=0.985
+ $X2=0 $Y2=0
cc_814 N_A_1482_48#_c_1174_n N_A_1224_74#_c_1283_n 0.0053332f $X=7.67 $Y=2.19
+ $X2=0 $Y2=0
cc_815 N_A_1482_48#_c_1178_n N_A_1224_74#_c_1283_n 0.0125972f $X=7.595 $Y=0.985
+ $X2=0 $Y2=0
cc_816 N_A_1482_48#_c_1180_n N_A_1224_74#_c_1283_n 6.55449e-19 $X=7.67 $Y=1.065
+ $X2=0 $Y2=0
cc_817 N_A_1482_48#_c_1175_n N_A_1224_74#_c_1284_n 0.00997859f $X=8.485 $Y=0.985
+ $X2=0 $Y2=0
cc_818 N_A_1482_48#_c_1177_n N_A_1224_74#_c_1284_n 0.0233867f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_819 N_A_1482_48#_c_1185_n N_A_1224_74#_c_1284_n 0.0116759f $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_820 N_A_1482_48#_c_1179_n N_A_1224_74#_c_1284_n 0.0109402f $X=8.727 $Y=0.985
+ $X2=0 $Y2=0
cc_821 N_A_1482_48#_c_1185_n N_VPWR_M1020_d 0.00365297f $X=8.885 $Y=1.85 $X2=0
+ $Y2=0
cc_822 N_A_1482_48#_c_1182_n N_VPWR_c_1489_n 0.00610146f $X=7.67 $Y=2.28 $X2=0
+ $Y2=0
cc_823 N_A_1482_48#_c_1183_n N_VPWR_c_1489_n 0.00131777f $X=8.555 $Y=2.335 $X2=0
+ $Y2=0
cc_824 N_A_1482_48#_c_1183_n N_VPWR_c_1490_n 0.00646407f $X=8.555 $Y=2.335 $X2=0
+ $Y2=0
cc_825 N_A_1482_48#_c_1183_n N_VPWR_c_1491_n 0.0463782f $X=8.555 $Y=2.335 $X2=0
+ $Y2=0
cc_826 N_A_1482_48#_c_1185_n N_VPWR_c_1491_n 0.012936f $X=8.885 $Y=1.85 $X2=0
+ $Y2=0
cc_827 N_A_1482_48#_c_1182_n N_VPWR_c_1497_n 0.00405364f $X=7.67 $Y=2.28 $X2=0
+ $Y2=0
cc_828 N_A_1482_48#_c_1182_n N_VPWR_c_1482_n 0.00489211f $X=7.67 $Y=2.28 $X2=0
+ $Y2=0
cc_829 N_A_1482_48#_c_1183_n N_VPWR_c_1482_n 0.011426f $X=8.555 $Y=2.335 $X2=0
+ $Y2=0
cc_830 N_A_1482_48#_c_1177_n N_Q_N_c_1770_n 0.018767f $X=8.885 $Y=1.765 $X2=0
+ $Y2=0
cc_831 N_A_1482_48#_c_1185_n N_Q_N_c_1770_n 0.00158159f $X=8.885 $Y=1.85 $X2=0
+ $Y2=0
cc_832 N_A_1482_48#_c_1185_n N_Q_N_c_1773_n 0.00456533f $X=8.885 $Y=1.85 $X2=0
+ $Y2=0
cc_833 N_A_1482_48#_c_1173_n N_VGND_c_1820_n 0.0147674f $X=7.485 $Y=0.9 $X2=0
+ $Y2=0
cc_834 N_A_1482_48#_c_1175_n N_VGND_c_1820_n 0.0137782f $X=8.485 $Y=0.985 $X2=0
+ $Y2=0
cc_835 N_A_1482_48#_c_1176_n N_VGND_c_1820_n 0.0110441f $X=8.65 $Y=0.58 $X2=0
+ $Y2=0
cc_836 N_A_1482_48#_c_1178_n N_VGND_c_1820_n 0.0129689f $X=7.595 $Y=0.985 $X2=0
+ $Y2=0
cc_837 N_A_1482_48#_c_1180_n N_VGND_c_1820_n 0.00131228f $X=7.67 $Y=1.065 $X2=0
+ $Y2=0
cc_838 N_A_1482_48#_c_1176_n N_VGND_c_1821_n 0.0454165f $X=8.65 $Y=0.58 $X2=0
+ $Y2=0
cc_839 N_A_1482_48#_c_1177_n N_VGND_c_1821_n 0.00455872f $X=8.885 $Y=1.765 $X2=0
+ $Y2=0
cc_840 N_A_1482_48#_c_1179_n N_VGND_c_1821_n 0.0145003f $X=8.727 $Y=0.985 $X2=0
+ $Y2=0
cc_841 N_A_1482_48#_c_1173_n N_VGND_c_1825_n 0.00383152f $X=7.485 $Y=0.9 $X2=0
+ $Y2=0
cc_842 N_A_1482_48#_c_1176_n N_VGND_c_1826_n 0.0215384f $X=8.65 $Y=0.58 $X2=0
+ $Y2=0
cc_843 N_A_1482_48#_c_1173_n N_VGND_c_1829_n 0.0075725f $X=7.485 $Y=0.9 $X2=0
+ $Y2=0
cc_844 N_A_1482_48#_c_1176_n N_VGND_c_1829_n 0.0177458f $X=8.65 $Y=0.58 $X2=0
+ $Y2=0
cc_845 N_A_1224_74#_M1008_g N_A_2026_424#_M1005_g 0.0197956f $X=10.515 $Y=0.645
+ $X2=0 $Y2=0
cc_846 N_A_1224_74#_c_1275_n N_A_2026_424#_c_1433_n 0.00994164f $X=10.5 $Y=1.955
+ $X2=0 $Y2=0
cc_847 N_A_1224_74#_c_1289_n N_A_2026_424#_c_1433_n 0.00588428f $X=10.5 $Y=2.045
+ $X2=0 $Y2=0
cc_848 N_A_1224_74#_c_1277_n N_A_2026_424#_c_1433_n 0.0214662f $X=10.5 $Y=1.43
+ $X2=0 $Y2=0
cc_849 N_A_1224_74#_c_1274_n N_A_2026_424#_c_1434_n 0.00517977f $X=10.41 $Y=1.43
+ $X2=0 $Y2=0
cc_850 N_A_1224_74#_M1008_g N_A_2026_424#_c_1434_n 0.0146713f $X=10.515 $Y=0.645
+ $X2=0 $Y2=0
cc_851 N_A_1224_74#_c_1277_n N_A_2026_424#_c_1434_n 6.73726e-19 $X=10.5 $Y=1.43
+ $X2=0 $Y2=0
cc_852 N_A_1224_74#_c_1275_n N_A_2026_424#_c_1435_n 0.0112992f $X=10.5 $Y=1.955
+ $X2=0 $Y2=0
cc_853 N_A_1224_74#_c_1289_n N_A_2026_424#_c_1435_n 0.0166377f $X=10.5 $Y=2.045
+ $X2=0 $Y2=0
cc_854 N_A_1224_74#_c_1275_n N_A_2026_424#_c_1436_n 0.00782285f $X=10.5 $Y=1.955
+ $X2=0 $Y2=0
cc_855 N_A_1224_74#_c_1277_n N_A_2026_424#_c_1436_n 0.0139388f $X=10.5 $Y=1.43
+ $X2=0 $Y2=0
cc_856 N_A_1224_74#_c_1274_n N_A_2026_424#_c_1437_n 0.0166486f $X=10.41 $Y=1.43
+ $X2=0 $Y2=0
cc_857 N_A_1224_74#_c_1275_n N_A_2026_424#_c_1437_n 7.34008e-19 $X=10.5 $Y=1.955
+ $X2=0 $Y2=0
cc_858 N_A_1224_74#_c_1277_n N_A_2026_424#_c_1437_n 8.33355e-19 $X=10.5 $Y=1.43
+ $X2=0 $Y2=0
cc_859 N_A_1224_74#_c_1301_n N_VPWR_c_1489_n 0.0264538f $X=7.495 $Y=2.53 $X2=0
+ $Y2=0
cc_860 N_A_1224_74#_c_1281_n N_VPWR_c_1489_n 0.0021468f $X=7.58 $Y=2.365 $X2=0
+ $Y2=0
cc_861 N_A_1224_74#_c_1286_n N_VPWR_c_1490_n 0.00393528f $X=8.63 $Y=2.28 $X2=0
+ $Y2=0
cc_862 N_A_1224_74#_c_1269_n N_VPWR_c_1491_n 0.0013401f $X=8.63 $Y=2.19 $X2=0
+ $Y2=0
cc_863 N_A_1224_74#_c_1286_n N_VPWR_c_1491_n 0.00764221f $X=8.63 $Y=2.28 $X2=0
+ $Y2=0
cc_864 N_A_1224_74#_c_1270_n N_VPWR_c_1491_n 0.00151008f $X=9.055 $Y=1.43 $X2=0
+ $Y2=0
cc_865 N_A_1224_74#_c_1272_n N_VPWR_c_1491_n 0.00556331f $X=9.145 $Y=1.765 $X2=0
+ $Y2=0
cc_866 N_A_1224_74#_c_1275_n N_VPWR_c_1492_n 0.00204674f $X=10.5 $Y=1.955 $X2=0
+ $Y2=0
cc_867 N_A_1224_74#_c_1289_n N_VPWR_c_1492_n 0.00449437f $X=10.5 $Y=2.045 $X2=0
+ $Y2=0
cc_868 N_A_1224_74#_c_1301_n N_VPWR_c_1497_n 0.0159863f $X=7.495 $Y=2.53 $X2=0
+ $Y2=0
cc_869 N_A_1224_74#_c_1272_n N_VPWR_c_1498_n 0.00461464f $X=9.145 $Y=1.765 $X2=0
+ $Y2=0
cc_870 N_A_1224_74#_c_1289_n N_VPWR_c_1498_n 0.00445665f $X=10.5 $Y=2.045 $X2=0
+ $Y2=0
cc_871 N_A_1224_74#_c_1286_n N_VPWR_c_1482_n 0.00489211f $X=8.63 $Y=2.28 $X2=0
+ $Y2=0
cc_872 N_A_1224_74#_c_1272_n N_VPWR_c_1482_n 0.00918106f $X=9.145 $Y=1.765 $X2=0
+ $Y2=0
cc_873 N_A_1224_74#_c_1289_n N_VPWR_c_1482_n 0.00862405f $X=10.5 $Y=2.045 $X2=0
+ $Y2=0
cc_874 N_A_1224_74#_c_1301_n N_VPWR_c_1482_n 0.0282176f $X=7.495 $Y=2.53 $X2=0
+ $Y2=0
cc_875 N_A_1224_74#_c_1301_n A_1465_471# 0.00449141f $X=7.495 $Y=2.53 $X2=-0.19
+ $Y2=-0.245
cc_876 N_A_1224_74#_c_1272_n N_Q_N_c_1770_n 0.0044298f $X=9.145 $Y=1.765 $X2=0
+ $Y2=0
cc_877 N_A_1224_74#_M1009_g N_Q_N_c_1770_n 0.0191689f $X=9.44 $Y=0.74 $X2=0
+ $Y2=0
cc_878 N_A_1224_74#_c_1274_n N_Q_N_c_1770_n 0.0449729f $X=10.41 $Y=1.43 $X2=0
+ $Y2=0
cc_879 N_A_1224_74#_c_1275_n N_Q_N_c_1770_n 0.0010753f $X=10.5 $Y=1.955 $X2=0
+ $Y2=0
cc_880 N_A_1224_74#_c_1272_n N_Q_N_c_1773_n 0.014297f $X=9.145 $Y=1.765 $X2=0
+ $Y2=0
cc_881 N_A_1224_74#_c_1289_n N_Q_N_c_1773_n 0.00385512f $X=10.5 $Y=2.045 $X2=0
+ $Y2=0
cc_882 N_A_1224_74#_M1027_g N_VGND_c_1820_n 0.0014914f $X=8.435 $Y=0.58 $X2=0
+ $Y2=0
cc_883 N_A_1224_74#_c_1297_n N_VGND_c_1820_n 0.0120929f $X=6.99 $Y=0.565 $X2=0
+ $Y2=0
cc_884 N_A_1224_74#_M1027_g N_VGND_c_1821_n 0.00378178f $X=8.435 $Y=0.58 $X2=0
+ $Y2=0
cc_885 N_A_1224_74#_c_1272_n N_VGND_c_1821_n 0.00633828f $X=9.145 $Y=1.765 $X2=0
+ $Y2=0
cc_886 N_A_1224_74#_M1009_g N_VGND_c_1821_n 0.017876f $X=9.44 $Y=0.74 $X2=0
+ $Y2=0
cc_887 N_A_1224_74#_M1008_g N_VGND_c_1822_n 0.00770628f $X=10.515 $Y=0.645 $X2=0
+ $Y2=0
cc_888 N_A_1224_74#_c_1297_n N_VGND_c_1825_n 0.0242914f $X=6.99 $Y=0.565 $X2=0
+ $Y2=0
cc_889 N_A_1224_74#_M1027_g N_VGND_c_1826_n 0.00434272f $X=8.435 $Y=0.58 $X2=0
+ $Y2=0
cc_890 N_A_1224_74#_M1009_g N_VGND_c_1827_n 0.00383152f $X=9.44 $Y=0.74 $X2=0
+ $Y2=0
cc_891 N_A_1224_74#_M1008_g N_VGND_c_1827_n 0.00461464f $X=10.515 $Y=0.645 $X2=0
+ $Y2=0
cc_892 N_A_1224_74#_M1027_g N_VGND_c_1829_n 0.00825979f $X=8.435 $Y=0.58 $X2=0
+ $Y2=0
cc_893 N_A_1224_74#_M1009_g N_VGND_c_1829_n 0.00762539f $X=9.44 $Y=0.74 $X2=0
+ $Y2=0
cc_894 N_A_1224_74#_M1008_g N_VGND_c_1829_n 0.00914043f $X=10.515 $Y=0.645 $X2=0
+ $Y2=0
cc_895 N_A_1224_74#_c_1297_n N_VGND_c_1829_n 0.02509f $X=6.99 $Y=0.565 $X2=0
+ $Y2=0
cc_896 N_A_2026_424#_c_1433_n N_VPWR_c_1492_n 0.00610705f $X=11.015 $Y=1.765
+ $X2=0 $Y2=0
cc_897 N_A_2026_424#_c_1435_n N_VPWR_c_1492_n 0.0542643f $X=10.275 $Y=2.27 $X2=0
+ $Y2=0
cc_898 N_A_2026_424#_c_1436_n N_VPWR_c_1492_n 0.0235211f $X=10.965 $Y=1.465
+ $X2=0 $Y2=0
cc_899 N_A_2026_424#_c_1435_n N_VPWR_c_1498_n 0.0108068f $X=10.275 $Y=2.27 $X2=0
+ $Y2=0
cc_900 N_A_2026_424#_c_1433_n N_VPWR_c_1499_n 0.00445602f $X=11.015 $Y=1.765
+ $X2=0 $Y2=0
cc_901 N_A_2026_424#_c_1433_n N_VPWR_c_1482_n 0.00861048f $X=11.015 $Y=1.765
+ $X2=0 $Y2=0
cc_902 N_A_2026_424#_c_1435_n N_VPWR_c_1482_n 0.00906421f $X=10.275 $Y=2.27
+ $X2=0 $Y2=0
cc_903 N_A_2026_424#_c_1434_n N_Q_N_c_1770_n 0.0605318f $X=10.3 $Y=0.64 $X2=0
+ $Y2=0
cc_904 N_A_2026_424#_c_1435_n N_Q_N_c_1770_n 0.0894769f $X=10.275 $Y=2.27 $X2=0
+ $Y2=0
cc_905 N_A_2026_424#_c_1437_n N_Q_N_c_1770_n 0.0205307f $X=10.315 $Y=1.465 $X2=0
+ $Y2=0
cc_906 N_A_2026_424#_M1005_g Q 0.00795463f $X=11.015 $Y=0.74 $X2=0 $Y2=0
cc_907 N_A_2026_424#_M1005_g Q 0.00263483f $X=11.015 $Y=0.74 $X2=0 $Y2=0
cc_908 N_A_2026_424#_c_1433_n Q 0.00169664f $X=11.015 $Y=1.765 $X2=0 $Y2=0
cc_909 N_A_2026_424#_c_1436_n Q 0.00233746f $X=10.965 $Y=1.465 $X2=0 $Y2=0
cc_910 N_A_2026_424#_c_1433_n Q 0.00408255f $X=11.015 $Y=1.765 $X2=0 $Y2=0
cc_911 N_A_2026_424#_c_1436_n Q 0.00140951f $X=10.965 $Y=1.465 $X2=0 $Y2=0
cc_912 N_A_2026_424#_c_1433_n Q 0.0109295f $X=11.015 $Y=1.765 $X2=0 $Y2=0
cc_913 N_A_2026_424#_M1005_g N_Q_c_1796_n 0.00406947f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_914 N_A_2026_424#_c_1433_n N_Q_c_1796_n 0.0126603f $X=11.015 $Y=1.765 $X2=0
+ $Y2=0
cc_915 N_A_2026_424#_c_1436_n N_Q_c_1796_n 0.0262113f $X=10.965 $Y=1.465 $X2=0
+ $Y2=0
cc_916 N_A_2026_424#_M1005_g N_VGND_c_1822_n 0.00357902f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_917 N_A_2026_424#_c_1433_n N_VGND_c_1822_n 0.00218979f $X=11.015 $Y=1.765
+ $X2=0 $Y2=0
cc_918 N_A_2026_424#_c_1434_n N_VGND_c_1822_n 0.0295846f $X=10.3 $Y=0.64 $X2=0
+ $Y2=0
cc_919 N_A_2026_424#_c_1436_n N_VGND_c_1822_n 0.0215504f $X=10.965 $Y=1.465
+ $X2=0 $Y2=0
cc_920 N_A_2026_424#_c_1434_n N_VGND_c_1827_n 0.011066f $X=10.3 $Y=0.64 $X2=0
+ $Y2=0
cc_921 N_A_2026_424#_M1005_g N_VGND_c_1828_n 0.00434272f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_922 N_A_2026_424#_M1005_g N_VGND_c_1829_n 0.00824463f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_923 N_A_2026_424#_c_1434_n N_VGND_c_1829_n 0.00915947f $X=10.3 $Y=0.64 $X2=0
+ $Y2=0
cc_924 N_VPWR_c_1484_n N_A_38_78#_c_1645_n 0.0231787f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_925 N_VPWR_c_1485_n N_A_38_78#_c_1645_n 0.00940122f $X=1.18 $Y=2.835 $X2=0
+ $Y2=0
cc_926 N_VPWR_c_1493_n N_A_38_78#_c_1645_n 0.0122114f $X=1.015 $Y=3.33 $X2=0
+ $Y2=0
cc_927 N_VPWR_c_1482_n N_A_38_78#_c_1645_n 0.0101411f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_928 N_VPWR_M1022_d N_A_38_78#_c_1647_n 0.00272596f $X=1.03 $Y=2.54 $X2=0
+ $Y2=0
cc_929 N_VPWR_c_1485_n N_A_38_78#_c_1647_n 0.0213829f $X=1.18 $Y=2.835 $X2=0
+ $Y2=0
cc_930 N_VPWR_c_1493_n N_A_38_78#_c_1647_n 0.00162049f $X=1.015 $Y=3.33 $X2=0
+ $Y2=0
cc_931 N_VPWR_c_1494_n N_A_38_78#_c_1647_n 0.00275677f $X=2.025 $Y=3.33 $X2=0
+ $Y2=0
cc_932 N_VPWR_c_1482_n N_A_38_78#_c_1647_n 0.00892716f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_933 N_VPWR_M1000_d N_A_38_78#_c_1648_n 0.00538932f $X=2.04 $Y=1.96 $X2=0
+ $Y2=0
cc_934 N_VPWR_c_1486_n N_A_38_78#_c_1648_n 0.0166706f $X=2.19 $Y=2.835 $X2=0
+ $Y2=0
cc_935 N_VPWR_c_1494_n N_A_38_78#_c_1648_n 7.47605e-19 $X=2.025 $Y=3.33 $X2=0
+ $Y2=0
cc_936 N_VPWR_c_1495_n N_A_38_78#_c_1648_n 0.00915743f $X=4.44 $Y=3.33 $X2=0
+ $Y2=0
cc_937 N_VPWR_c_1482_n N_A_38_78#_c_1648_n 0.0193758f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_938 N_VPWR_c_1484_n N_A_38_78#_c_1651_n 0.00766412f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_939 N_VPWR_c_1493_n N_A_38_78#_c_1651_n 4.31008e-19 $X=1.015 $Y=3.33 $X2=0
+ $Y2=0
cc_940 N_VPWR_c_1482_n N_A_38_78#_c_1651_n 0.00120957f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_941 N_VPWR_c_1494_n N_A_38_78#_c_1652_n 0.00568973f $X=2.025 $Y=3.33 $X2=0
+ $Y2=0
cc_942 N_VPWR_c_1482_n N_A_38_78#_c_1652_n 0.011076f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_943 N_VPWR_c_1495_n N_A_38_78#_c_1653_n 0.00493758f $X=4.44 $Y=3.33 $X2=0
+ $Y2=0
cc_944 N_VPWR_c_1482_n N_A_38_78#_c_1653_n 0.00718941f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_945 N_VPWR_c_1491_n Q_N 0.00163554f $X=8.92 $Y=2.27 $X2=0 $Y2=0
cc_946 N_VPWR_c_1492_n Q_N 3.35434e-19 $X=10.79 $Y=1.985 $X2=0 $Y2=0
cc_947 N_VPWR_c_1498_n Q_N 0.0313273f $X=10.61 $Y=3.33 $X2=0 $Y2=0
cc_948 N_VPWR_c_1482_n Q_N 0.0254862f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_949 N_VPWR_c_1492_n Q 0.0456259f $X=10.79 $Y=1.985 $X2=0 $Y2=0
cc_950 N_VPWR_c_1499_n Q 0.0159324f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_951 N_VPWR_c_1482_n Q 0.0131546f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_952 N_A_38_78#_c_1637_n A_125_78# 0.00236678f $X=0.69 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_953 N_A_38_78#_c_1637_n N_VGND_c_1817_n 0.00157034f $X=0.69 $Y=0.745 $X2=0
+ $Y2=0
cc_954 N_A_38_78#_c_1642_n N_VGND_c_1817_n 0.00465719f $X=0.335 $Y=0.6 $X2=0
+ $Y2=0
cc_955 N_A_38_78#_c_1637_n N_VGND_c_1823_n 0.00520932f $X=0.69 $Y=0.745 $X2=0
+ $Y2=0
cc_956 N_A_38_78#_c_1642_n N_VGND_c_1823_n 0.0131067f $X=0.335 $Y=0.6 $X2=0
+ $Y2=0
cc_957 N_A_38_78#_c_1637_n N_VGND_c_1829_n 0.0102476f $X=0.69 $Y=0.745 $X2=0
+ $Y2=0
cc_958 N_A_38_78#_c_1642_n N_VGND_c_1829_n 0.0117869f $X=0.335 $Y=0.6 $X2=0
+ $Y2=0
cc_959 N_Q_N_c_1770_n N_VGND_c_1821_n 0.0296698f $X=9.725 $Y=0.515 $X2=0 $Y2=0
cc_960 N_Q_N_c_1773_n N_VGND_c_1821_n 0.00437693f $X=9.37 $Y=1.985 $X2=0 $Y2=0
cc_961 N_Q_N_c_1770_n N_VGND_c_1827_n 0.0173129f $X=9.725 $Y=0.515 $X2=0 $Y2=0
cc_962 N_Q_N_c_1770_n N_VGND_c_1829_n 0.0143301f $X=9.725 $Y=0.515 $X2=0 $Y2=0
cc_963 Q N_VGND_c_1822_n 0.0312622f $X=11.195 $Y=0.47 $X2=0 $Y2=0
cc_964 Q N_VGND_c_1828_n 0.0163488f $X=11.195 $Y=0.47 $X2=0 $Y2=0
cc_965 Q N_VGND_c_1829_n 0.0134757f $X=11.195 $Y=0.47 $X2=0 $Y2=0
