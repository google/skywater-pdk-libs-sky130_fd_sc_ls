* File: sky130_fd_sc_ls__dlrtp_2.spice
* Created: Fri Aug 28 13:19:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dlrtp_2.pex.spice"
.subckt sky130_fd_sc_ls__dlrtp_2  VNB VPB D GATE RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_D_M1006_g N_A_27_392#_M1006_s VNB NSHORT L=0.15 W=0.55
+ AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1019 N_A_235_74#_M1019_d N_GATE_M1019_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1021_d N_A_235_74#_M1021_g N_A_347_98#_M1021_s VNB NSHORT L=0.15
+ W=0.74 AD=0.205216 AS=0.2701 PD=1.59797 PS=2.21 NRD=36.048 NRS=12.972 M=1
+ R=4.93333 SA=75000.3 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1000 A_568_74# N_A_27_392#_M1000_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.177484 PD=0.88 PS=1.38203 NRD=12.18 NRS=15.936 M=1 R=4.26667
+ SA=75000.8 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1001 N_A_646_74#_M1001_d N_A_347_98#_M1001_g A_568_74# VNB NSHORT L=0.15
+ W=0.64 AD=0.194158 AS=0.0768 PD=1.42491 PS=0.88 NRD=16.872 NRS=12.18 M=1
+ R=4.26667 SA=75001.2 SB=75001 A=0.096 P=1.58 MULT=1
MM1015 A_784_81# N_A_235_74#_M1015_g N_A_646_74#_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.127417 PD=0.66 PS=0.935094 NRD=18.564 NRS=48.564 M=1
+ R=2.8 SA=75001.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_832_55#_M1016_g A_784_81# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 A_1060_74# N_A_646_74#_M1011_g N_A_832_55#_M1011_s VNB NSHORT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_RESET_B_M1003_g A_1060_74# VNB NSHORT L=0.15 W=0.74
+ AD=0.1628 AS=0.0888 PD=1.18 PS=0.98 NRD=14.592 NRS=10.536 M=1 R=4.93333
+ SA=75000.6 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1004 N_Q_M1004_d N_A_832_55#_M1004_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1073 AS=0.1628 PD=1.03 PS=1.18 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1013 N_Q_M1004_d N_A_832_55#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1073 AS=0.2553 PD=1.03 PS=2.17 NRD=1.62 NRS=9.72 M=1 R=4.93333 SA=75001.6
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1012 N_VPWR_M1012_d N_D_M1012_g N_A_27_392#_M1012_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.23945 AS=0.2478 PD=1.6 PS=2.27 NRD=53.9386 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1009 N_A_235_74#_M1009_d N_GATE_M1009_g N_VPWR_M1012_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.23945 PD=2.27 PS=1.6 NRD=2.3443 NRS=53.9386 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1017 N_VPWR_M1017_d N_A_235_74#_M1017_g N_A_347_98#_M1017_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.222623 AS=0.2478 PD=1.4563 PS=2.27 NRD=49.25 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1010 A_565_392# N_A_27_392#_M1010_g N_VPWR_M1017_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.265027 PD=1.27 PS=1.7337 NRD=15.7403 NRS=18.6953 M=1 R=6.66667
+ SA=75000.7 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1008 N_A_646_74#_M1008_d N_A_235_74#_M1008_g A_565_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.234366 AS=0.135 PD=1.9507 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75001.2 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1018 A_756_508# N_A_347_98#_M1018_g N_A_646_74#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.11235 AS=0.0984338 PD=0.955 PS=0.819296 NRD=99.6623 NRS=46.886 M=1
+ R=2.8 SA=75001.6 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_832_55#_M1005_g A_756_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.125618 AS=0.11235 PD=0.968182 PS=0.955 NRD=75.0373 NRS=99.6623 M=1 R=2.8
+ SA=75002.3 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1007 N_A_832_55#_M1007_d N_A_646_74#_M1007_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.334982 PD=1.42 PS=2.58182 NRD=1.7533 NRS=37.8043 M=1
+ R=7.46667 SA=75001.3 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1014_d N_RESET_B_M1014_g N_A_832_55#_M1007_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1002 N_Q_M1002_d N_A_832_55#_M1002_g N_VPWR_M1014_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1764 AS=0.224 PD=1.435 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.3 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1020 N_Q_M1002_d N_A_832_55#_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1764 AS=0.3696 PD=1.435 PS=2.9 NRD=4.3931 NRS=7.8997 M=1 R=7.46667
+ SA=75002.7 SB=75000.3 A=0.168 P=2.54 MULT=1
DX22_noxref VNB VPB NWDIODE A=14.0988 P=18.88
c_1045 A_784_81# 0 1.78997e-19 $X=3.92 $Y=0.405
*
.include "sky130_fd_sc_ls__dlrtp_2.pxi.spice"
*
.ends
*
*
