* File: sky130_fd_sc_ls__mux2i_4.spice
* Created: Fri Aug 28 13:30:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__mux2i_4.pex.spice"
.subckt sky130_fd_sc_ls__mux2i_4  VNB VPB A1 A0 S Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* S	S
* A0	A0
* A1	A1
* VPB	VPB
* VNB	VNB
MM1011 N_A_114_85#_M1011_d N_A1_M1011_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1012 N_A_114_85#_M1011_d N_A1_M1012_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1032 N_A_114_85#_M1032_d N_A1_M1032_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.13505 AS=0.1036 PD=1.105 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1034 N_A_114_85#_M1032_d N_A1_M1034_g N_Y_M1034_s VNB NSHORT L=0.15 W=0.74
+ AD=0.13505 AS=0.1036 PD=1.105 PS=1.02 NRD=13.776 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75002 A=0.111 P=1.78 MULT=1
MM1004 N_A_475_85#_M1004_d N_A0_M1004_g N_Y_M1034_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1027 N_A_475_85#_M1004_d N_A0_M1027_g N_Y_M1027_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.12025 PD=1.09 PS=1.065 NRD=0 NRS=3.24 M=1 R=4.93333 SA=75002.5
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1028 N_A_475_85#_M1028_d N_A0_M1028_g N_Y_M1027_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.12025 PD=1.02 PS=1.065 NRD=0 NRS=4.044 M=1 R=4.93333 SA=75003
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1031 N_A_475_85#_M1028_d N_A0_M1031_g N_Y_M1031_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_475_85#_M1006_d N_A_1030_268#_M1006_g N_VGND_M1006_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.36 PD=1.02 PS=2.83 NRD=0 NRS=69.96 M=1 R=4.93333
+ SA=75000.3 SB=75003.9 A=0.111 P=1.78 MULT=1
MM1007 N_A_475_85#_M1006_d N_A_1030_268#_M1007_g N_VGND_M1007_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.20315 PD=1.02 PS=1.49 NRD=0 NRS=35.592 M=1
+ R=4.93333 SA=75000.7 SB=75003.5 A=0.111 P=1.78 MULT=1
MM1021 N_A_475_85#_M1021_d N_A_1030_268#_M1021_g N_VGND_M1007_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.20315 PD=1.02 PS=1.49 NRD=0 NRS=35.592 M=1
+ R=4.93333 SA=75001.2 SB=75003.3 A=0.111 P=1.78 MULT=1
MM1024 N_A_475_85#_M1021_d N_A_1030_268#_M1024_g N_VGND_M1024_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.1036 AS=0.19615 PD=1.02 PS=1.41 NRD=0 NRS=34.056 M=1
+ R=4.93333 SA=75001.6 SB=75002.9 A=0.111 P=1.78 MULT=1
MM1005 N_A_114_85#_M1005_d N_S_M1005_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.19615 PD=1.02 PS=1.41 NRD=0 NRS=34.056 M=1 R=4.93333 SA=75002.2
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1009 N_A_114_85#_M1005_d N_S_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1887 PD=1.02 PS=1.25 NRD=0 NRS=18.648 M=1 R=4.93333 SA=75002.6
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1019 N_A_114_85#_M1019_d N_S_M1019_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1887 PD=1.02 PS=1.25 NRD=0 NRS=18.648 M=1 R=4.93333 SA=75003.3
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1022 N_A_114_85#_M1019_d N_S_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.7
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1013 N_A_1030_268#_M1013_d N_S_M1013_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2627 AS=0.1295 PD=2.19 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75004.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A1_M1000_g N_A_116_368#_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.6 A=0.168 P=2.54 MULT=1
MM1014 N_Y_M1014_d N_A1_M1014_g N_A_116_368#_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1015 N_Y_M1014_d N_A1_M1015_g N_A_116_368#_M1015_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1025 N_Y_M1025_d N_A1_M1025_g N_A_116_368#_M1015_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1736 AS=0.168 PD=1.43 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1001 N_A_478_368#_M1001_d N_A0_M1001_g N_Y_M1025_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1904 AS=0.1736 PD=1.46 PS=1.43 NRD=8.7862 NRS=3.5066 M=1 R=7.46667
+ SA=75002 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1010 N_A_478_368#_M1001_d N_A0_M1010_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1904 AS=0.196 PD=1.46 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.5 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1020 N_A_478_368#_M1020_d N_A0_M1020_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1029 N_A_478_368#_M1020_d N_A0_M1029_g N_Y_M1029_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.3864 PD=1.47 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.5 SB=75000.3 A=0.168 P=2.54 MULT=1
MM1002 N_A_116_368#_M1002_d N_A_1030_268#_M1002_g N_VPWR_M1002_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.7504 PD=1.42 PS=3.58 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.6 SB=75004.3 A=0.168 P=2.54 MULT=1
MM1018 N_A_116_368#_M1002_d N_A_1030_268#_M1018_g N_VPWR_M1018_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75001 SB=75003.9 A=0.168 P=2.54 MULT=1
MM1023 N_A_116_368#_M1023_d N_A_1030_268#_M1023_g N_VPWR_M1018_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.2128 AS=0.168 PD=1.5 PS=1.42 NRD=4.3931 NRS=1.7533 M=1
+ R=7.46667 SA=75001.5 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1030 N_A_116_368#_M1023_d N_A_1030_268#_M1030_g N_VPWR_M1030_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.2128 AS=0.196 PD=1.5 PS=1.47 NRD=13.1793 NRS=1.7533 M=1
+ R=7.46667 SA=75002 SB=75002.9 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1030_s N_S_M1003_g N_A_478_368#_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1008_d N_S_M1008_g N_A_478_368#_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1008_d N_S_M1016_g N_A_478_368#_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75001.4 A=0.168 P=2.54 MULT=1
MM1033 N_VPWR_M1033_d N_S_M1033_g N_A_478_368#_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2128 AS=0.168 PD=1.68571 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004 SB=75000.9 A=0.168 P=2.54 MULT=1
MM1017 N_A_1030_268#_M1017_d N_S_M1017_g N_VPWR_M1033_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.126 AS=0.1596 PD=1.14 PS=1.26429 NRD=2.3443 NRS=15.2281 M=1 R=5.6
+ SA=75004.5 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1026 N_A_1030_268#_M1017_d N_S_M1026_g N_VPWR_M1026_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.126 AS=0.2478 PD=1.14 PS=2.27 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75004.9 SB=75000.2 A=0.126 P=1.98 MULT=1
DX35_noxref VNB VPB NWDIODE A=19.4556 P=24.64
*
.include "sky130_fd_sc_ls__mux2i_4.pxi.spice"
*
.ends
*
*
