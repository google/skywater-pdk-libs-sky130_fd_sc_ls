* File: sky130_fd_sc_ls__decaphe_2.spice
* Created: Fri Aug 28 13:12:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__decaphe_2.pex.spice"
.subckt sky130_fd_sc_ls__decaphe_2  VNB VPB VGND VPWR
* 
* VPWR	VPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1000 N_VPWR_M1000_s N_VGND_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.17 W=1.255
+ AD=0.3263 AS=0.3263 PD=3.03 PS=3.03 NRD=0 NRS=0 M=1 R=7.38235 SA=85000.2
+ SB=85000.2 A=0.21335 P=2.85 MULT=1
DX1_noxref VNB VPB NWDIODE A=2.4924 P=6.4
*
.include "sky130_fd_sc_ls__decaphe_2.pxi.spice"
*
.ends
*
*
