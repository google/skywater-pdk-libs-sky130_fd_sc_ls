* File: sky130_fd_sc_ls__a221oi_2.spice
* Created: Fri Aug 28 12:53:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a221oi_2.pex.spice"
.subckt sky130_fd_sc_ls__a221oi_2  VNB VPB C1 B1 B2 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1015 N_Y_M1015_d N_C1_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.111 PD=2.01 PS=1.04 NRD=0 NRS=1.62 M=1 R=4.93333 SA=75000.2
+ SB=75004.7 A=0.111 P=1.78 MULT=1
MM1019 N_Y_M1019_d N_C1_M1019_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.111 PD=1.02 PS=1.04 NRD=0 NRS=1.62 M=1 R=4.93333 SA=75000.6
+ SB=75004.3 A=0.111 P=1.78 MULT=1
MM1003 N_A_293_74#_M1003_d N_B1_M1003_g N_Y_M1019_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1184 AS=0.1036 PD=1.06 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75003.8 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_B2_M1001_g N_A_293_74#_M1003_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1443 AS=0.1184 PD=1.13 PS=1.06 NRD=5.664 NRS=6.48 M=1 R=4.93333
+ SA=75001.5 SB=75003.4 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1001_d N_B2_M1008_g N_A_293_74#_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1443 AS=0.1036 PD=1.13 PS=1.02 NRD=12.156 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1014 N_A_293_74#_M1008_s N_B1_M1014_g N_Y_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1184 PD=1.02 PS=1.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1014_s N_A1_M1006_g N_A_675_74#_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1184 AS=0.2479 PD=1.06 PS=1.41 NRD=6.48 NRS=0 M=1 R=4.93333 SA=75003
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1005 N_A_675_74#_M1006_s N_A2_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2479 AS=0.1295 PD=1.41 PS=1.09 NRD=0 NRS=4.86 M=1 R=4.93333 SA=75003.8
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_A_675_74#_M1007_d N_A2_M1007_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=6.48 M=1 R=4.93333 SA=75004.3
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1012 N_Y_M1012_d N_A1_M1012_g N_A_675_74#_M1007_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_Y_M1016_d N_C1_M1016_g N_A_29_368#_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1017 N_Y_M1016_d N_C1_M1017_g N_A_29_368#_M1017_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75002 A=0.168 P=2.54 MULT=1
MM1000 N_A_294_368#_M1000_d N_B1_M1000_g N_A_29_368#_M1017_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.1848 AS=0.168 PD=1.45 PS=1.42 NRD=4.3931 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1011 N_A_29_368#_M1011_d N_B2_M1011_g N_A_294_368#_M1000_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.1848 PD=1.42 PS=1.45 NRD=1.7533 NRS=4.3931 M=1 R=7.46667
+ SA=75001.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1018 N_A_29_368#_M1011_d N_B2_M1018_g N_A_294_368#_M1018_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1002 N_A_294_368#_M1018_s N_B1_M1002_g N_A_29_368#_M1002_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1004 N_A_294_368#_M1004_d N_A1_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1009_d N_A2_M1009_g N_A_294_368#_M1004_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1010 N_VPWR_M1009_d N_A2_M1010_g N_A_294_368#_M1010_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1013 N_A_294_368#_M1010_s N_A1_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ls__a221oi_2.pxi.spice"
*
.ends
*
*
