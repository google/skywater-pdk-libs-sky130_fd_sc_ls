* File: sky130_fd_sc_ls__a21bo_1.pxi.spice
* Created: Wed Sep  2 10:47:52 2020
* 
x_PM_SKY130_FD_SC_LS__A21BO_1%A2 N_A2_c_74_n N_A2_c_75_n N_A2_c_80_n
+ N_A2_M1004_g N_A2_M1001_g N_A2_c_77_n A2 N_A2_c_78_n
+ PM_SKY130_FD_SC_LS__A21BO_1%A2
x_PM_SKY130_FD_SC_LS__A21BO_1%A1 N_A1_M1007_g N_A1_c_107_n N_A1_M1008_g A1
+ PM_SKY130_FD_SC_LS__A21BO_1%A1
x_PM_SKY130_FD_SC_LS__A21BO_1%A_272_110# N_A_272_110#_M1006_s
+ N_A_272_110#_M1005_s N_A_272_110#_c_142_n N_A_272_110#_M1003_g
+ N_A_272_110#_c_143_n N_A_272_110#_c_152_n N_A_272_110#_M1000_g
+ N_A_272_110#_c_144_n N_A_272_110#_c_145_n N_A_272_110#_c_146_n
+ N_A_272_110#_c_147_n N_A_272_110#_c_148_n N_A_272_110#_c_155_n
+ N_A_272_110#_c_149_n N_A_272_110#_c_150_n
+ PM_SKY130_FD_SC_LS__A21BO_1%A_272_110#
x_PM_SKY130_FD_SC_LS__A21BO_1%B1_N N_B1_N_c_208_n N_B1_N_M1005_g N_B1_N_M1006_g
+ B1_N PM_SKY130_FD_SC_LS__A21BO_1%B1_N
x_PM_SKY130_FD_SC_LS__A21BO_1%A_194_136# N_A_194_136#_M1007_d
+ N_A_194_136#_M1000_d N_A_194_136#_M1002_g N_A_194_136#_c_241_n
+ N_A_194_136#_M1009_g N_A_194_136#_c_242_n N_A_194_136#_c_262_n
+ N_A_194_136#_c_252_n N_A_194_136#_c_246_n N_A_194_136#_c_247_n
+ N_A_194_136#_c_248_n N_A_194_136#_c_249_n N_A_194_136#_c_243_n
+ N_A_194_136#_c_244_n PM_SKY130_FD_SC_LS__A21BO_1%A_194_136#
x_PM_SKY130_FD_SC_LS__A21BO_1%A_34_392# N_A_34_392#_M1004_s N_A_34_392#_M1008_d
+ N_A_34_392#_c_323_n N_A_34_392#_c_324_n N_A_34_392#_c_325_n
+ N_A_34_392#_c_326_n N_A_34_392#_c_327_n PM_SKY130_FD_SC_LS__A21BO_1%A_34_392#
x_PM_SKY130_FD_SC_LS__A21BO_1%VPWR N_VPWR_M1004_d N_VPWR_M1005_d N_VPWR_c_354_n
+ N_VPWR_c_355_n VPWR N_VPWR_c_356_n N_VPWR_c_357_n N_VPWR_c_353_n
+ N_VPWR_c_359_n N_VPWR_c_360_n PM_SKY130_FD_SC_LS__A21BO_1%VPWR
x_PM_SKY130_FD_SC_LS__A21BO_1%X N_X_M1002_d N_X_M1009_d N_X_c_391_n N_X_c_392_n
+ X X X X N_X_c_393_n PM_SKY130_FD_SC_LS__A21BO_1%X
x_PM_SKY130_FD_SC_LS__A21BO_1%VGND N_VGND_M1001_s N_VGND_M1003_d N_VGND_M1006_d
+ N_VGND_c_416_n N_VGND_c_417_n N_VGND_c_418_n N_VGND_c_419_n N_VGND_c_420_n
+ N_VGND_c_421_n N_VGND_c_422_n N_VGND_c_423_n VGND N_VGND_c_424_n
+ N_VGND_c_425_n N_VGND_c_426_n N_VGND_c_427_n PM_SKY130_FD_SC_LS__A21BO_1%VGND
cc_1 VNB N_A2_c_74_n 0.00824473f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.485
cc_2 VNB N_A2_c_75_n 0.0144971f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.795
cc_3 VNB N_A2_M1001_g 0.0108761f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1
cc_4 VNB N_A2_c_77_n 0.0711591f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=0.405
cc_5 VNB N_A2_c_78_n 0.0087821f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.405
cc_6 VNB N_A1_M1007_g 0.0190091f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.885
cc_7 VNB N_A1_c_107_n 0.0161762f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.46
cc_8 VNB A1 0.00835686f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1
cc_9 VNB N_A_272_110#_c_142_n 0.0179505f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.395
cc_10 VNB N_A_272_110#_c_143_n 0.00637459f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=0.405
cc_11 VNB N_A_272_110#_c_144_n 0.0182102f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.405
cc_12 VNB N_A_272_110#_c_145_n 0.00578316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_272_110#_c_146_n 0.00108341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_272_110#_c_147_n 0.006464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_272_110#_c_148_n 0.0492722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_272_110#_c_149_n 0.00458865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_272_110#_c_150_n 0.0306579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_N_c_208_n 0.0401678f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.485
cc_19 VNB N_B1_N_M1006_g 0.0340384f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.57
cc_20 VNB B1_N 0.00383465f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1
cc_21 VNB N_A_194_136#_M1002_g 0.0293029f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1
cc_22 VNB N_A_194_136#_c_241_n 0.0353214f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=0.405
cc_23 VNB N_A_194_136#_c_242_n 0.00491491f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.405
cc_24 VNB N_A_194_136#_c_243_n 0.0025844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_194_136#_c_244_n 0.00483797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_353_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_391_n 0.0285266f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1
cc_28 VNB N_X_c_392_n 0.0179941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_393_n 0.0251251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_416_n 0.015592f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=0.405
cc_31 VNB N_VGND_c_417_n 0.0314912f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.405
cc_32 VNB N_VGND_c_418_n 0.0085077f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.405
cc_33 VNB N_VGND_c_419_n 0.0252027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_420_n 0.0179973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_421_n 0.00311272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_422_n 0.0294344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_423_n 0.00413547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_424_n 0.0209588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_425_n 0.0216364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_426_n 0.243723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_427_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_A2_c_75_n 0.0112012f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.795
cc_43 VPB N_A2_c_80_n 0.0297875f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.885
cc_44 VPB N_A1_c_107_n 0.0335282f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=2.46
cc_45 VPB A1 0.00514464f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1
cc_46 VPB N_A_272_110#_c_143_n 0.00753824f $X=-0.19 $Y=1.66 $X2=0.46 $Y2=0.405
cc_47 VPB N_A_272_110#_c_152_n 0.0258564f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_48 VPB N_A_272_110#_c_146_n 0.0102106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_272_110#_c_148_n 0.0171171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_272_110#_c_155_n 0.0131545f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_B1_N_c_208_n 0.0281918f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.485
cc_52 VPB N_A_194_136#_c_241_n 0.0288543f $X=-0.19 $Y=1.66 $X2=0.46 $Y2=0.405
cc_53 VPB N_A_194_136#_c_246_n 6.9775e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_194_136#_c_247_n 0.00251211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_194_136#_c_248_n 0.0323224f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_194_136#_c_249_n 0.00179604f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_194_136#_c_243_n 0.00615429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_34_392#_c_323_n 0.013293f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.395
cc_59 VPB N_A_34_392#_c_324_n 0.0360166f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1
cc_60 VPB N_A_34_392#_c_325_n 0.00382599f $X=-0.19 $Y=1.66 $X2=0.46 $Y2=0.405
cc_61 VPB N_A_34_392#_c_326_n 0.00293494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_34_392#_c_327_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.405
cc_63 VPB N_VPWR_c_354_n 0.00835244f $X=-0.19 $Y=1.66 $X2=0.46 $Y2=0.405
cc_64 VPB N_VPWR_c_355_n 0.0171686f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.405
cc_65 VPB N_VPWR_c_356_n 0.0608614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_357_n 0.0188734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_353_n 0.107436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_359_n 0.0243021f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_360_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB X 0.0131928f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.405
cc_71 VPB X 0.0443399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_X_c_393_n 0.00755811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 N_A2_c_77_n N_A1_M1007_g 0.0362809f $X=0.46 $Y=0.405 $X2=0 $Y2=0
cc_74 N_A2_c_74_n N_A1_c_107_n 0.0362809f $X=0.52 $Y=1.485 $X2=0 $Y2=0
cc_75 N_A2_c_75_n N_A1_c_107_n 0.00512744f $X=0.52 $Y=1.795 $X2=0 $Y2=0
cc_76 N_A2_c_80_n N_A1_c_107_n 0.0172837f $X=0.52 $Y=1.885 $X2=0 $Y2=0
cc_77 N_A2_c_74_n A1 0.0100513f $X=0.52 $Y=1.485 $X2=0 $Y2=0
cc_78 N_A2_M1001_g N_A_194_136#_c_242_n 3.74963e-19 $X=0.535 $Y=1 $X2=0 $Y2=0
cc_79 N_A2_M1001_g N_A_194_136#_c_252_n 4.60392e-19 $X=0.535 $Y=1 $X2=0 $Y2=0
cc_80 N_A2_c_80_n N_A_34_392#_c_323_n 0.0017173f $X=0.52 $Y=1.885 $X2=0 $Y2=0
cc_81 N_A2_c_80_n N_A_34_392#_c_324_n 0.0106338f $X=0.52 $Y=1.885 $X2=0 $Y2=0
cc_82 N_A2_c_80_n N_A_34_392#_c_325_n 0.0165078f $X=0.52 $Y=1.885 $X2=0 $Y2=0
cc_83 N_A2_c_80_n N_A_34_392#_c_327_n 6.36743e-19 $X=0.52 $Y=1.885 $X2=0 $Y2=0
cc_84 N_A2_c_80_n N_VPWR_c_354_n 0.00507786f $X=0.52 $Y=1.885 $X2=0 $Y2=0
cc_85 N_A2_c_80_n N_VPWR_c_353_n 0.00861479f $X=0.52 $Y=1.885 $X2=0 $Y2=0
cc_86 N_A2_c_80_n N_VPWR_c_359_n 0.00445602f $X=0.52 $Y=1.885 $X2=0 $Y2=0
cc_87 N_A2_M1001_g N_VGND_c_416_n 0.00907665f $X=0.535 $Y=1 $X2=0 $Y2=0
cc_88 N_A2_c_77_n N_VGND_c_416_n 0.0105624f $X=0.46 $Y=0.405 $X2=0 $Y2=0
cc_89 N_A2_c_78_n N_VGND_c_416_n 0.0300105f $X=0.27 $Y=0.405 $X2=0 $Y2=0
cc_90 N_A2_c_74_n N_VGND_c_419_n 0.00110067f $X=0.52 $Y=1.485 $X2=0 $Y2=0
cc_91 N_A2_M1001_g N_VGND_c_419_n 0.0211774f $X=0.535 $Y=1 $X2=0 $Y2=0
cc_92 N_A2_c_77_n N_VGND_c_419_n 0.00158926f $X=0.46 $Y=0.405 $X2=0 $Y2=0
cc_93 N_A2_c_78_n N_VGND_c_419_n 0.0223651f $X=0.27 $Y=0.405 $X2=0 $Y2=0
cc_94 N_A2_c_77_n N_VGND_c_420_n 0.0108f $X=0.46 $Y=0.405 $X2=0 $Y2=0
cc_95 N_A2_c_78_n N_VGND_c_420_n 0.0215843f $X=0.27 $Y=0.405 $X2=0 $Y2=0
cc_96 N_A2_c_77_n N_VGND_c_426_n 0.0124008f $X=0.46 $Y=0.405 $X2=0 $Y2=0
cc_97 N_A2_c_78_n N_VGND_c_426_n 0.0110944f $X=0.27 $Y=0.405 $X2=0 $Y2=0
cc_98 N_A1_M1007_g N_A_272_110#_c_142_n 0.0158982f $X=0.895 $Y=1 $X2=0 $Y2=0
cc_99 N_A1_c_107_n N_A_272_110#_c_143_n 0.00517498f $X=1 $Y=1.885 $X2=0 $Y2=0
cc_100 N_A1_c_107_n N_A_272_110#_c_152_n 0.00877946f $X=1 $Y=1.885 $X2=0 $Y2=0
cc_101 N_A1_c_107_n N_A_272_110#_c_145_n 0.0201051f $X=1 $Y=1.885 $X2=0 $Y2=0
cc_102 A1 N_A_272_110#_c_145_n 0.00311702f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_103 N_A1_M1007_g N_A_194_136#_c_242_n 0.00522309f $X=0.895 $Y=1 $X2=0 $Y2=0
cc_104 N_A1_M1007_g N_A_194_136#_c_252_n 0.00304397f $X=0.895 $Y=1 $X2=0 $Y2=0
cc_105 N_A1_c_107_n N_A_194_136#_c_252_n 0.00444086f $X=1 $Y=1.885 $X2=0 $Y2=0
cc_106 A1 N_A_194_136#_c_252_n 0.0278432f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_107 N_A1_M1007_g N_A_194_136#_c_243_n 2.19497e-19 $X=0.895 $Y=1 $X2=0 $Y2=0
cc_108 A1 N_A_194_136#_c_243_n 0.020131f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_109 N_A1_c_107_n N_A_34_392#_c_324_n 6.36743e-19 $X=1 $Y=1.885 $X2=0 $Y2=0
cc_110 N_A1_c_107_n N_A_34_392#_c_325_n 0.0149383f $X=1 $Y=1.885 $X2=0 $Y2=0
cc_111 A1 N_A_34_392#_c_325_n 0.0305802f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_112 N_A1_c_107_n N_A_34_392#_c_326_n 0.00237082f $X=1 $Y=1.885 $X2=0 $Y2=0
cc_113 A1 N_A_34_392#_c_326_n 0.0221184f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_114 N_A1_c_107_n N_A_34_392#_c_327_n 0.0104821f $X=1 $Y=1.885 $X2=0 $Y2=0
cc_115 N_A1_c_107_n N_VPWR_c_354_n 0.00507786f $X=1 $Y=1.885 $X2=0 $Y2=0
cc_116 N_A1_c_107_n N_VPWR_c_356_n 0.00445602f $X=1 $Y=1.885 $X2=0 $Y2=0
cc_117 N_A1_c_107_n N_VPWR_c_353_n 0.0085802f $X=1 $Y=1.885 $X2=0 $Y2=0
cc_118 N_A1_M1007_g N_VGND_c_416_n 0.00320336f $X=0.895 $Y=1 $X2=0 $Y2=0
cc_119 N_A1_M1007_g N_VGND_c_417_n 5.76731e-19 $X=0.895 $Y=1 $X2=0 $Y2=0
cc_120 N_A1_M1007_g N_VGND_c_419_n 8.05577e-19 $X=0.895 $Y=1 $X2=0 $Y2=0
cc_121 A1 N_VGND_c_419_n 0.00551077f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_122 N_A1_M1007_g N_VGND_c_424_n 0.0037378f $X=0.895 $Y=1 $X2=0 $Y2=0
cc_123 N_A1_M1007_g N_VGND_c_426_n 0.00454494f $X=0.895 $Y=1 $X2=0 $Y2=0
cc_124 N_A_272_110#_c_146_n N_B1_N_c_208_n 0.00256654f $X=2.08 $Y=1.605
+ $X2=-0.19 $Y2=-0.245
cc_125 N_A_272_110#_c_147_n N_B1_N_c_208_n 0.00126721f $X=2.08 $Y=1.265
+ $X2=-0.19 $Y2=-0.245
cc_126 N_A_272_110#_c_148_n N_B1_N_c_208_n 0.0210311f $X=2.08 $Y=1.265 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A_272_110#_c_155_n N_B1_N_c_208_n 0.00595754f $X=2.53 $Y=1.985
+ $X2=-0.19 $Y2=-0.245
cc_128 N_A_272_110#_c_150_n N_B1_N_c_208_n 0.00121279f $X=2.555 $Y=0.645
+ $X2=-0.19 $Y2=-0.245
cc_129 N_A_272_110#_c_147_n N_B1_N_M1006_g 4.83119e-19 $X=2.08 $Y=1.265 $X2=0
+ $Y2=0
cc_130 N_A_272_110#_c_148_n N_B1_N_M1006_g 0.00321701f $X=2.08 $Y=1.265 $X2=0
+ $Y2=0
cc_131 N_A_272_110#_c_149_n N_B1_N_M1006_g 0.00406543f $X=2.08 $Y=1.1 $X2=0
+ $Y2=0
cc_132 N_A_272_110#_c_150_n N_B1_N_M1006_g 0.0118322f $X=2.555 $Y=0.645 $X2=0
+ $Y2=0
cc_133 N_A_272_110#_c_147_n B1_N 0.0193295f $X=2.08 $Y=1.265 $X2=0 $Y2=0
cc_134 N_A_272_110#_c_148_n B1_N 0.00169009f $X=2.08 $Y=1.265 $X2=0 $Y2=0
cc_135 N_A_272_110#_c_155_n B1_N 0.00986955f $X=2.53 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_272_110#_c_150_n B1_N 0.0139046f $X=2.555 $Y=0.645 $X2=0 $Y2=0
cc_137 N_A_272_110#_c_150_n N_A_194_136#_M1002_g 2.74584e-19 $X=2.555 $Y=0.645
+ $X2=0 $Y2=0
cc_138 N_A_272_110#_c_155_n N_A_194_136#_c_241_n 2.23035e-19 $X=2.53 $Y=1.985
+ $X2=0 $Y2=0
cc_139 N_A_272_110#_c_142_n N_A_194_136#_c_242_n 0.00263456f $X=1.435 $Y=1.395
+ $X2=0 $Y2=0
cc_140 N_A_272_110#_c_142_n N_A_194_136#_c_262_n 0.0186854f $X=1.435 $Y=1.395
+ $X2=0 $Y2=0
cc_141 N_A_272_110#_c_147_n N_A_194_136#_c_262_n 0.014001f $X=2.08 $Y=1.265
+ $X2=0 $Y2=0
cc_142 N_A_272_110#_c_148_n N_A_194_136#_c_262_n 0.00145776f $X=2.08 $Y=1.265
+ $X2=0 $Y2=0
cc_143 N_A_272_110#_c_144_n N_A_194_136#_c_246_n 4.53459e-19 $X=1.915 $Y=1.47
+ $X2=0 $Y2=0
cc_144 N_A_272_110#_c_146_n N_A_194_136#_c_246_n 0.00694643f $X=2.08 $Y=1.605
+ $X2=0 $Y2=0
cc_145 N_A_272_110#_c_152_n N_A_194_136#_c_247_n 4.43985e-19 $X=1.45 $Y=1.885
+ $X2=0 $Y2=0
cc_146 N_A_272_110#_M1005_s N_A_194_136#_c_248_n 0.0114482f $X=2.405 $Y=1.84
+ $X2=0 $Y2=0
cc_147 N_A_272_110#_c_144_n N_A_194_136#_c_248_n 0.00128732f $X=1.915 $Y=1.47
+ $X2=0 $Y2=0
cc_148 N_A_272_110#_c_146_n N_A_194_136#_c_248_n 0.0202781f $X=2.08 $Y=1.605
+ $X2=0 $Y2=0
cc_149 N_A_272_110#_c_148_n N_A_194_136#_c_248_n 0.0014957f $X=2.08 $Y=1.265
+ $X2=0 $Y2=0
cc_150 N_A_272_110#_c_155_n N_A_194_136#_c_248_n 0.0296882f $X=2.53 $Y=1.985
+ $X2=0 $Y2=0
cc_151 N_A_272_110#_c_155_n N_A_194_136#_c_249_n 0.0101888f $X=2.53 $Y=1.985
+ $X2=0 $Y2=0
cc_152 N_A_272_110#_c_142_n N_A_194_136#_c_243_n 0.00286167f $X=1.435 $Y=1.395
+ $X2=0 $Y2=0
cc_153 N_A_272_110#_c_143_n N_A_194_136#_c_243_n 0.00676459f $X=1.45 $Y=1.795
+ $X2=0 $Y2=0
cc_154 N_A_272_110#_c_152_n N_A_194_136#_c_243_n 0.00272187f $X=1.45 $Y=1.885
+ $X2=0 $Y2=0
cc_155 N_A_272_110#_c_144_n N_A_194_136#_c_243_n 0.0121573f $X=1.915 $Y=1.47
+ $X2=0 $Y2=0
cc_156 N_A_272_110#_c_146_n N_A_194_136#_c_243_n 0.0449041f $X=2.08 $Y=1.605
+ $X2=0 $Y2=0
cc_157 N_A_272_110#_c_148_n N_A_194_136#_c_243_n 0.00189136f $X=2.08 $Y=1.265
+ $X2=0 $Y2=0
cc_158 N_A_272_110#_c_152_n N_A_34_392#_c_326_n 0.00292913f $X=1.45 $Y=1.885
+ $X2=0 $Y2=0
cc_159 N_A_272_110#_c_152_n N_A_34_392#_c_327_n 0.00926234f $X=1.45 $Y=1.885
+ $X2=0 $Y2=0
cc_160 N_A_272_110#_c_152_n N_VPWR_c_356_n 0.00445602f $X=1.45 $Y=1.885 $X2=0
+ $Y2=0
cc_161 N_A_272_110#_c_152_n N_VPWR_c_353_n 0.00863237f $X=1.45 $Y=1.885 $X2=0
+ $Y2=0
cc_162 N_A_272_110#_c_150_n N_X_c_391_n 0.00129386f $X=2.555 $Y=0.645 $X2=0
+ $Y2=0
cc_163 N_A_272_110#_c_142_n N_VGND_c_417_n 0.00848694f $X=1.435 $Y=1.395 $X2=0
+ $Y2=0
cc_164 N_A_272_110#_c_144_n N_VGND_c_417_n 0.00271372f $X=1.915 $Y=1.47 $X2=0
+ $Y2=0
cc_165 N_A_272_110#_c_150_n N_VGND_c_417_n 0.0378925f $X=2.555 $Y=0.645 $X2=0
+ $Y2=0
cc_166 N_A_272_110#_c_150_n N_VGND_c_418_n 0.0223843f $X=2.555 $Y=0.645 $X2=0
+ $Y2=0
cc_167 N_A_272_110#_c_150_n N_VGND_c_422_n 0.028291f $X=2.555 $Y=0.645 $X2=0
+ $Y2=0
cc_168 N_A_272_110#_c_142_n N_VGND_c_424_n 0.00322089f $X=1.435 $Y=1.395 $X2=0
+ $Y2=0
cc_169 N_A_272_110#_c_142_n N_VGND_c_426_n 0.00381775f $X=1.435 $Y=1.395 $X2=0
+ $Y2=0
cc_170 N_A_272_110#_c_150_n N_VGND_c_426_n 0.0235701f $X=2.555 $Y=0.645 $X2=0
+ $Y2=0
cc_171 N_B1_N_M1006_g N_A_194_136#_M1002_g 0.0242832f $X=2.77 $Y=0.645 $X2=0
+ $Y2=0
cc_172 B1_N N_A_194_136#_M1002_g 8.42001e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_173 N_B1_N_c_208_n N_A_194_136#_c_241_n 0.0462257f $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_174 B1_N N_A_194_136#_c_241_n 8.4674e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_175 N_B1_N_c_208_n N_A_194_136#_c_248_n 0.0212461f $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_176 N_B1_N_c_208_n N_A_194_136#_c_249_n 0.00859635f $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_B1_N_c_208_n N_A_194_136#_c_244_n 0.00150548f $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_178 B1_N N_A_194_136#_c_244_n 0.0131032f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_179 N_B1_N_c_208_n N_VPWR_c_355_n 0.00641581f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_180 N_B1_N_c_208_n N_VPWR_c_356_n 0.00402388f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_181 N_B1_N_c_208_n N_VPWR_c_353_n 0.00462577f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_182 N_B1_N_M1006_g N_X_c_391_n 0.00118491f $X=2.77 $Y=0.645 $X2=0 $Y2=0
cc_183 N_B1_N_M1006_g N_VGND_c_418_n 0.00360765f $X=2.77 $Y=0.645 $X2=0 $Y2=0
cc_184 N_B1_N_M1006_g N_VGND_c_422_n 0.00433162f $X=2.77 $Y=0.645 $X2=0 $Y2=0
cc_185 N_B1_N_M1006_g N_VGND_c_426_n 0.00822133f $X=2.77 $Y=0.645 $X2=0 $Y2=0
cc_186 N_A_194_136#_c_262_n N_A_34_392#_c_326_n 0.0015886f $X=1.575 $Y=1.195
+ $X2=0 $Y2=0
cc_187 N_A_194_136#_c_246_n N_A_34_392#_c_326_n 0.00701355f $X=1.667 $Y=2.032
+ $X2=0 $Y2=0
cc_188 N_A_194_136#_c_247_n N_A_34_392#_c_327_n 0.0206684f $X=1.675 $Y=2.46
+ $X2=0 $Y2=0
cc_189 N_A_194_136#_c_248_n N_VPWR_M1005_d 0.0110254f $X=3.085 $Y=2.325 $X2=0
+ $Y2=0
cc_190 N_A_194_136#_c_249_n N_VPWR_M1005_d 0.00490214f $X=3.17 $Y=2.24 $X2=0
+ $Y2=0
cc_191 N_A_194_136#_c_241_n N_VPWR_c_355_n 0.0124058f $X=3.29 $Y=1.765 $X2=0
+ $Y2=0
cc_192 N_A_194_136#_c_248_n N_VPWR_c_355_n 0.022613f $X=3.085 $Y=2.325 $X2=0
+ $Y2=0
cc_193 N_A_194_136#_c_247_n N_VPWR_c_356_n 0.00816563f $X=1.675 $Y=2.46 $X2=0
+ $Y2=0
cc_194 N_A_194_136#_c_241_n N_VPWR_c_357_n 0.00413917f $X=3.29 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A_194_136#_c_241_n N_VPWR_c_353_n 0.00821361f $X=3.29 $Y=1.765 $X2=0
+ $Y2=0
cc_196 N_A_194_136#_c_247_n N_VPWR_c_353_n 0.0067588f $X=1.675 $Y=2.46 $X2=0
+ $Y2=0
cc_197 N_A_194_136#_M1002_g N_X_c_391_n 0.00764773f $X=3.245 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A_194_136#_M1002_g N_X_c_392_n 0.00524476f $X=3.245 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A_194_136#_c_241_n N_X_c_392_n 7.28954e-19 $X=3.29 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A_194_136#_c_244_n N_X_c_392_n 0.00908321f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_201 N_A_194_136#_c_241_n X 0.0089135f $X=3.29 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A_194_136#_c_249_n X 0.0303104f $X=3.17 $Y=2.24 $X2=0 $Y2=0
cc_203 N_A_194_136#_c_248_n X 0.0136806f $X=3.085 $Y=2.325 $X2=0 $Y2=0
cc_204 N_A_194_136#_M1002_g N_X_c_393_n 0.00431388f $X=3.245 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A_194_136#_c_241_n N_X_c_393_n 0.00986012f $X=3.29 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A_194_136#_c_249_n N_X_c_393_n 0.00520007f $X=3.17 $Y=2.24 $X2=0 $Y2=0
cc_207 N_A_194_136#_c_244_n N_X_c_393_n 0.0248017f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_208 N_A_194_136#_c_262_n N_VGND_M1003_d 0.00401902f $X=1.575 $Y=1.195 $X2=0
+ $Y2=0
cc_209 N_A_194_136#_c_243_n N_VGND_M1003_d 7.55995e-19 $X=1.667 $Y=1.94 $X2=0
+ $Y2=0
cc_210 N_A_194_136#_c_242_n N_VGND_c_416_n 0.00758818f $X=1.13 $Y=0.805 $X2=0
+ $Y2=0
cc_211 N_A_194_136#_c_242_n N_VGND_c_417_n 0.0109353f $X=1.13 $Y=0.805 $X2=0
+ $Y2=0
cc_212 N_A_194_136#_c_262_n N_VGND_c_417_n 0.0169764f $X=1.575 $Y=1.195 $X2=0
+ $Y2=0
cc_213 N_A_194_136#_M1002_g N_VGND_c_418_n 0.00359027f $X=3.245 $Y=0.74 $X2=0
+ $Y2=0
cc_214 N_A_194_136#_c_244_n N_VGND_c_418_n 0.00117839f $X=3.25 $Y=1.485 $X2=0
+ $Y2=0
cc_215 N_A_194_136#_c_242_n N_VGND_c_419_n 4.90416e-19 $X=1.13 $Y=0.805 $X2=0
+ $Y2=0
cc_216 N_A_194_136#_c_252_n N_VGND_c_419_n 0.00604662f $X=1.315 $Y=1.195 $X2=0
+ $Y2=0
cc_217 N_A_194_136#_c_242_n N_VGND_c_424_n 0.00697694f $X=1.13 $Y=0.805 $X2=0
+ $Y2=0
cc_218 N_A_194_136#_M1002_g N_VGND_c_425_n 0.00434272f $X=3.245 $Y=0.74 $X2=0
+ $Y2=0
cc_219 N_A_194_136#_M1002_g N_VGND_c_426_n 0.00824739f $X=3.245 $Y=0.74 $X2=0
+ $Y2=0
cc_220 N_A_194_136#_c_242_n N_VGND_c_426_n 0.0108859f $X=1.13 $Y=0.805 $X2=0
+ $Y2=0
cc_221 N_A_34_392#_c_325_n N_VPWR_M1004_d 0.00279158f $X=1.06 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_222 N_A_34_392#_c_324_n N_VPWR_c_354_n 0.0455206f $X=0.295 $Y=2.815 $X2=0
+ $Y2=0
cc_223 N_A_34_392#_c_325_n N_VPWR_c_354_n 0.016109f $X=1.06 $Y=2.035 $X2=0 $Y2=0
cc_224 N_A_34_392#_c_327_n N_VPWR_c_354_n 0.0455206f $X=1.225 $Y=2.815 $X2=0
+ $Y2=0
cc_225 N_A_34_392#_c_327_n N_VPWR_c_356_n 0.014552f $X=1.225 $Y=2.815 $X2=0
+ $Y2=0
cc_226 N_A_34_392#_c_324_n N_VPWR_c_353_n 0.0120466f $X=0.295 $Y=2.815 $X2=0
+ $Y2=0
cc_227 N_A_34_392#_c_327_n N_VPWR_c_353_n 0.0119791f $X=1.225 $Y=2.815 $X2=0
+ $Y2=0
cc_228 N_A_34_392#_c_324_n N_VPWR_c_359_n 0.0145938f $X=0.295 $Y=2.815 $X2=0
+ $Y2=0
cc_229 N_A_34_392#_c_323_n N_VGND_c_419_n 0.0114724f $X=0.295 $Y=2.12 $X2=0
+ $Y2=0
cc_230 N_A_34_392#_c_325_n N_VGND_c_419_n 6.30365e-19 $X=1.06 $Y=2.035 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_355_n X 0.0273968f $X=3.065 $Y=2.745 $X2=0 $Y2=0
cc_232 N_VPWR_c_357_n X 0.0144126f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_233 N_VPWR_c_353_n X 0.0119295f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_234 N_X_c_391_n N_VGND_c_418_n 0.021263f $X=3.46 $Y=0.515 $X2=0 $Y2=0
cc_235 N_X_c_391_n N_VGND_c_425_n 0.0203646f $X=3.46 $Y=0.515 $X2=0 $Y2=0
cc_236 N_X_c_391_n N_VGND_c_426_n 0.0167997f $X=3.46 $Y=0.515 $X2=0 $Y2=0
cc_237 N_VGND_c_419_n A_122_136# 0.0015121f $X=0.32 $Y=1.09 $X2=-0.19 $Y2=-0.245
