* File: sky130_fd_sc_ls__einvn_1.pxi.spice
* Created: Fri Aug 28 13:23:26 2020
* 
x_PM_SKY130_FD_SC_LS__EINVN_1%A_22_46# N_A_22_46#_M1004_s N_A_22_46#_M1005_s
+ N_A_22_46#_c_42_n N_A_22_46#_c_43_n N_A_22_46#_M1000_g N_A_22_46#_c_44_n
+ N_A_22_46#_c_45_n N_A_22_46#_c_75_p N_A_22_46#_c_46_n N_A_22_46#_c_47_n
+ N_A_22_46#_c_50_n N_A_22_46#_c_48_n PM_SKY130_FD_SC_LS__EINVN_1%A_22_46#
x_PM_SKY130_FD_SC_LS__EINVN_1%TE_B N_TE_B_c_85_n N_TE_B_M1005_g N_TE_B_c_86_n
+ N_TE_B_M1004_g N_TE_B_c_87_n N_TE_B_c_92_n N_TE_B_M1003_g TE_B N_TE_B_c_89_n
+ PM_SKY130_FD_SC_LS__EINVN_1%TE_B
x_PM_SKY130_FD_SC_LS__EINVN_1%A N_A_c_129_n N_A_M1002_g N_A_c_130_n N_A_M1001_g
+ A N_A_c_131_n PM_SKY130_FD_SC_LS__EINVN_1%A
x_PM_SKY130_FD_SC_LS__EINVN_1%VPWR N_VPWR_M1005_d N_VPWR_c_160_n VPWR
+ N_VPWR_c_161_n N_VPWR_c_162_n N_VPWR_c_159_n N_VPWR_c_164_n
+ PM_SKY130_FD_SC_LS__EINVN_1%VPWR
x_PM_SKY130_FD_SC_LS__EINVN_1%Z N_Z_M1002_d N_Z_M1001_d N_Z_c_185_n N_Z_c_183_n
+ N_Z_c_184_n Z Z PM_SKY130_FD_SC_LS__EINVN_1%Z
x_PM_SKY130_FD_SC_LS__EINVN_1%VGND N_VGND_M1004_d N_VGND_c_205_n VGND
+ N_VGND_c_206_n N_VGND_c_207_n N_VGND_c_208_n N_VGND_c_209_n
+ PM_SKY130_FD_SC_LS__EINVN_1%VGND
cc_1 VNB N_A_22_46#_c_42_n 0.0464381f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=0.35
cc_2 VNB N_A_22_46#_c_43_n 0.0137421f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=0.425
cc_3 VNB N_A_22_46#_c_44_n 0.0189997f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=0.92
cc_4 VNB N_A_22_46#_c_45_n 0.0201391f $X=-0.19 $Y=-0.245 $X2=0.195 $Y2=1.93
cc_5 VNB N_A_22_46#_c_46_n 0.066973f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.395
cc_6 VNB N_A_22_46#_c_47_n 0.0247124f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.085
cc_7 VNB N_A_22_46#_c_48_n 0.0199392f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.395
cc_8 VNB N_TE_B_c_85_n 0.0295297f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.9
cc_9 VNB N_TE_B_c_86_n 0.019244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_TE_B_c_87_n 0.0161663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB TE_B 0.00343606f $X=-0.19 $Y=-0.245 $X2=0.195 $Y2=1.93
cc_12 VNB N_TE_B_c_89_n 0.00549215f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.395
cc_13 VNB N_A_c_129_n 0.0207146f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.9
cc_14 VNB N_A_c_130_n 0.0311384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_c_131_n 0.00786651f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=0.425
cc_16 VNB N_VPWR_c_159_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=0.395
cc_17 VNB N_Z_c_183_n 0.0228045f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=0.87
cc_18 VNB N_Z_c_184_n 0.0420195f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=0.56
cc_19 VNB N_VGND_c_205_n 0.0100327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_206_n 0.0257484f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=0.87
cc_21 VNB N_VGND_c_207_n 0.0344986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_208_n 0.169809f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=0.395
cc_23 VNB N_VGND_c_209_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VPB N_A_22_46#_c_45_n 0.0140148f $X=-0.19 $Y=1.66 $X2=0.195 $Y2=1.93
cc_25 VPB N_A_22_46#_c_50_n 0.046307f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.075
cc_26 VPB N_TE_B_c_85_n 0.0418316f $X=-0.19 $Y=1.66 $X2=0.455 $Y2=0.9
cc_27 VPB N_TE_B_c_87_n 0.0175905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_28 VPB N_TE_B_c_92_n 0.0172282f $X=-0.19 $Y=1.66 $X2=1.255 $Y2=0.35
cc_29 VPB TE_B 0.0016346f $X=-0.19 $Y=1.66 $X2=0.195 $Y2=1.93
cc_30 VPB N_TE_B_c_89_n 9.38834e-19 $X=-0.19 $Y=1.66 $X2=0.615 $Y2=0.395
cc_31 VPB N_A_c_130_n 0.0311811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_A_c_131_n 0.00689703f $X=-0.19 $Y=1.66 $X2=1.33 $Y2=0.425
cc_33 VPB N_VPWR_c_160_n 0.0216517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_161_n 0.0304179f $X=-0.19 $Y=1.66 $X2=1.33 $Y2=0.87
cc_35 VPB N_VPWR_c_162_n 0.0341405f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_159_n 0.0801174f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=0.395
cc_37 VPB N_VPWR_c_164_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_Z_c_185_n 0.0146645f $X=-0.19 $Y=1.66 $X2=1.33 $Y2=0.425
cc_39 VPB N_Z_c_183_n 0.0140697f $X=-0.19 $Y=1.66 $X2=1.33 $Y2=0.87
cc_40 VPB Z 0.0401493f $X=-0.19 $Y=1.66 $X2=0.195 $Y2=1.93
cc_41 N_A_22_46#_c_45_n N_TE_B_c_85_n 0.00666373f $X=0.195 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_42 N_A_22_46#_c_47_n N_TE_B_c_85_n 0.00671511f $X=0.605 $Y=1.085 $X2=-0.19
+ $Y2=-0.245
cc_43 N_A_22_46#_c_50_n N_TE_B_c_85_n 0.0131248f $X=0.555 $Y=2.075 $X2=-0.19
+ $Y2=-0.245
cc_44 N_A_22_46#_c_42_n N_TE_B_c_86_n 0.00493939f $X=1.255 $Y=0.35 $X2=0 $Y2=0
cc_45 N_A_22_46#_c_43_n N_TE_B_c_86_n 0.0115742f $X=1.33 $Y=0.425 $X2=0 $Y2=0
cc_46 N_A_22_46#_c_44_n N_TE_B_c_86_n 0.00482005f $X=0.44 $Y=0.92 $X2=0 $Y2=0
cc_47 N_A_22_46#_c_45_n N_TE_B_c_86_n 0.00404556f $X=0.195 $Y=1.93 $X2=0 $Y2=0
cc_48 N_A_22_46#_c_47_n N_TE_B_c_86_n 0.00379808f $X=0.605 $Y=1.085 $X2=0 $Y2=0
cc_49 N_A_22_46#_c_48_n N_TE_B_c_86_n 0.0023126f $X=0.78 $Y=0.395 $X2=0 $Y2=0
cc_50 N_A_22_46#_c_43_n N_TE_B_c_87_n 0.00986428f $X=1.33 $Y=0.425 $X2=0 $Y2=0
cc_51 N_A_22_46#_c_43_n TE_B 0.00122005f $X=1.33 $Y=0.425 $X2=0 $Y2=0
cc_52 N_A_22_46#_c_45_n N_TE_B_c_89_n 0.0256401f $X=0.195 $Y=1.93 $X2=0 $Y2=0
cc_53 N_A_22_46#_c_47_n N_TE_B_c_89_n 0.022249f $X=0.605 $Y=1.085 $X2=0 $Y2=0
cc_54 N_A_22_46#_c_50_n N_TE_B_c_89_n 0.0174267f $X=0.555 $Y=2.075 $X2=0 $Y2=0
cc_55 N_A_22_46#_c_42_n N_A_c_129_n 0.0253488f $X=1.255 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_56 N_A_22_46#_c_43_n N_A_c_130_n 0.0253488f $X=1.33 $Y=0.425 $X2=0 $Y2=0
cc_57 N_A_22_46#_c_43_n N_A_c_131_n 4.88499e-19 $X=1.33 $Y=0.425 $X2=0 $Y2=0
cc_58 N_A_22_46#_c_50_n N_VPWR_c_160_n 0.0428227f $X=0.555 $Y=2.075 $X2=0 $Y2=0
cc_59 N_A_22_46#_c_50_n N_VPWR_c_161_n 0.00514082f $X=0.555 $Y=2.075 $X2=0 $Y2=0
cc_60 N_A_22_46#_c_50_n N_VPWR_c_159_n 0.00896853f $X=0.555 $Y=2.075 $X2=0 $Y2=0
cc_61 N_A_22_46#_c_43_n N_Z_c_184_n 0.0019742f $X=1.33 $Y=0.425 $X2=0 $Y2=0
cc_62 N_A_22_46#_c_42_n N_VGND_c_205_n 0.0256607f $X=1.255 $Y=0.35 $X2=0 $Y2=0
cc_63 N_A_22_46#_c_43_n N_VGND_c_205_n 0.016172f $X=1.33 $Y=0.425 $X2=0 $Y2=0
cc_64 N_A_22_46#_c_44_n N_VGND_c_205_n 0.0419197f $X=0.44 $Y=0.92 $X2=0 $Y2=0
cc_65 N_A_22_46#_c_75_p N_VGND_c_205_n 0.0248316f $X=0.615 $Y=0.395 $X2=0 $Y2=0
cc_66 N_A_22_46#_c_48_n N_VGND_c_205_n 0.00277657f $X=0.78 $Y=0.395 $X2=0 $Y2=0
cc_67 N_A_22_46#_c_42_n N_VGND_c_206_n 0.00502076f $X=1.255 $Y=0.35 $X2=0 $Y2=0
cc_68 N_A_22_46#_c_75_p N_VGND_c_206_n 0.0454726f $X=0.615 $Y=0.395 $X2=0 $Y2=0
cc_69 N_A_22_46#_c_46_n N_VGND_c_206_n 0.0116198f $X=0.615 $Y=0.395 $X2=0 $Y2=0
cc_70 N_A_22_46#_c_42_n N_VGND_c_207_n 0.0045897f $X=1.255 $Y=0.35 $X2=0 $Y2=0
cc_71 N_A_22_46#_c_42_n N_VGND_c_208_n 0.0093352f $X=1.255 $Y=0.35 $X2=0 $Y2=0
cc_72 N_A_22_46#_c_75_p N_VGND_c_208_n 0.0228727f $X=0.615 $Y=0.395 $X2=0 $Y2=0
cc_73 N_A_22_46#_c_46_n N_VGND_c_208_n 0.0114391f $X=0.615 $Y=0.395 $X2=0 $Y2=0
cc_74 N_A_22_46#_c_48_n N_VGND_c_208_n 0.00394079f $X=0.78 $Y=0.395 $X2=0 $Y2=0
cc_75 N_TE_B_c_87_n N_A_c_130_n 0.00859903f $X=1.225 $Y=1.685 $X2=0 $Y2=0
cc_76 N_TE_B_c_92_n N_A_c_130_n 0.058129f $X=1.315 $Y=1.765 $X2=0 $Y2=0
cc_77 TE_B N_A_c_130_n 0.0013061f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_78 N_TE_B_c_85_n N_A_c_131_n 5.88986e-19 $X=0.78 $Y=1.845 $X2=0 $Y2=0
cc_79 N_TE_B_c_86_n N_A_c_131_n 0.001417f $X=0.82 $Y=1.43 $X2=0 $Y2=0
cc_80 N_TE_B_c_87_n N_A_c_131_n 0.00125263f $X=1.225 $Y=1.685 $X2=0 $Y2=0
cc_81 TE_B N_A_c_131_n 0.0229497f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_82 N_TE_B_c_85_n N_VPWR_c_160_n 0.00881142f $X=0.78 $Y=1.845 $X2=0 $Y2=0
cc_83 N_TE_B_c_87_n N_VPWR_c_160_n 0.00408348f $X=1.225 $Y=1.685 $X2=0 $Y2=0
cc_84 N_TE_B_c_92_n N_VPWR_c_160_n 0.0219159f $X=1.315 $Y=1.765 $X2=0 $Y2=0
cc_85 TE_B N_VPWR_c_160_n 0.0120168f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_86 N_TE_B_c_89_n N_VPWR_c_160_n 0.0120133f $X=1.085 $Y=1.605 $X2=0 $Y2=0
cc_87 N_TE_B_c_85_n N_VPWR_c_161_n 0.00339865f $X=0.78 $Y=1.845 $X2=0 $Y2=0
cc_88 N_TE_B_c_92_n N_VPWR_c_162_n 0.00413917f $X=1.315 $Y=1.765 $X2=0 $Y2=0
cc_89 N_TE_B_c_85_n N_VPWR_c_159_n 0.00431146f $X=0.78 $Y=1.845 $X2=0 $Y2=0
cc_90 N_TE_B_c_92_n N_VPWR_c_159_n 0.00817532f $X=1.315 $Y=1.765 $X2=0 $Y2=0
cc_91 N_TE_B_c_92_n N_Z_c_185_n 0.00310499f $X=1.315 $Y=1.765 $X2=0 $Y2=0
cc_92 N_TE_B_c_86_n N_VGND_c_205_n 0.00300331f $X=0.82 $Y=1.43 $X2=0 $Y2=0
cc_93 N_TE_B_c_87_n N_VGND_c_205_n 0.00162249f $X=1.225 $Y=1.685 $X2=0 $Y2=0
cc_94 N_TE_B_c_89_n N_VGND_c_205_n 0.0285478f $X=1.085 $Y=1.605 $X2=0 $Y2=0
cc_95 N_A_c_130_n N_VPWR_c_160_n 0.00347662f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A_c_130_n N_VPWR_c_162_n 0.00411612f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A_c_130_n N_VPWR_c_159_n 0.00752013f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A_c_130_n N_Z_c_185_n 0.0064962f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_c_131_n N_Z_c_185_n 0.015552f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_100 N_A_c_129_n N_Z_c_183_n 0.00337861f $X=1.72 $Y=1.35 $X2=0 $Y2=0
cc_101 N_A_c_130_n N_Z_c_183_n 0.0104829f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_c_131_n N_Z_c_183_n 0.0332868f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_103 N_A_c_129_n N_Z_c_184_n 0.0126824f $X=1.72 $Y=1.35 $X2=0 $Y2=0
cc_104 N_A_c_130_n N_Z_c_184_n 0.0012398f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A_c_131_n N_Z_c_184_n 0.0145144f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_106 N_A_c_130_n Z 0.0147462f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A_c_129_n N_VGND_c_205_n 0.00292024f $X=1.72 $Y=1.35 $X2=0 $Y2=0
cc_108 N_A_c_129_n N_VGND_c_207_n 0.00467453f $X=1.72 $Y=1.35 $X2=0 $Y2=0
cc_109 N_A_c_129_n N_VGND_c_208_n 0.00505379f $X=1.72 $Y=1.35 $X2=0 $Y2=0
cc_110 N_VPWR_c_160_n N_Z_c_185_n 0.032773f $X=1.09 $Y=2.115 $X2=0 $Y2=0
cc_111 N_VPWR_c_162_n Z 0.0243207f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_112 N_VPWR_c_159_n Z 0.0200272f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_113 N_Z_c_184_n N_VGND_c_205_n 0.0230605f $X=1.935 $Y=0.645 $X2=0 $Y2=0
cc_114 N_Z_c_184_n N_VGND_c_207_n 0.0157999f $X=1.935 $Y=0.645 $X2=0 $Y2=0
cc_115 N_Z_c_184_n N_VGND_c_208_n 0.0184123f $X=1.935 $Y=0.645 $X2=0 $Y2=0
