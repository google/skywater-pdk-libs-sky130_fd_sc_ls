* NGSPICE file created from sky130_fd_sc_ls__nand4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
M1000 VPWR A_N a_27_158# VPB phighvt w=840000u l=150000u
+  ad=5.0862e+12p pd=2.218e+07u as=2.52e+11p ps=2.28e+06u
M1001 a_225_74# B a_656_74# VNB nshort w=740000u l=150000u
+  ad=1.01295e+12p pd=1.022e+07u as=8.399e+11p ps=8.19e+06u
M1002 a_225_74# a_27_158# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1003 Y B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=2.2512e+12p pd=1.298e+07u as=0p ps=0u
M1004 VPWR D Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_1025_158# D VGND VNB nshort w=740000u l=150000u
+  ad=1.0287e+12p pd=1.022e+07u as=6.9465e+11p ps=6.36e+06u
M1006 a_1025_158# C a_656_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_656_74# B a_225_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_27_158# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_225_74# a_27_158# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR C Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1025_158# C a_656_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1025_158# D VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND D a_1025_158# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_225_74# B a_656_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_27_158# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_656_74# B a_225_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_158# A_N VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A_N a_27_158# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=1.962e+11p ps=2.05e+06u
M1021 Y a_27_158# a_225_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y D VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y a_27_158# a_225_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_656_74# C a_1025_158# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_656_74# C a_1025_158# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND D a_1025_158# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

