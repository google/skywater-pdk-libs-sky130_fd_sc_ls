* File: sky130_fd_sc_ls__einvn_8.pex.spice
* Created: Wed Sep  2 11:06:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__EINVN_8%A_126_74# 1 2 7 8 9 11 12 14 16 17 19 21 22
+ 24 26 27 29 31 32 34 36 37 39 41 42 44 46 48 49 50 51 52 53 54 57 63 64 69
c152 64 0 3.46022e-20 $X=1.19 $Y=0.49
c153 57 0 1.57621e-19 $X=0.78 $Y=1.985
c154 42 0 1.6104e-19 $X=4.9 $Y=1.26
c155 8 0 1.9459e-20 $X=1.355 $Y=1.26
r156 69 72 6.39005 $w=7.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=1.17
+ $X2=0.985 $Y2=1.335
r157 69 71 0.778307 $w=7.38e-07 $l=4e-08 $layer=LI1_cond $X=0.985 $Y=1.17
+ $X2=0.985 $Y2=1.13
r158 69 70 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.19
+ $Y=1.17 $X2=1.19 $Y2=1.17
r159 67 71 10.9789 $w=6.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.02 $Y=0.515
+ $X2=1.02 $Y2=1.13
r160 64 70 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=1.19 $Y=0.49
+ $X2=1.19 $Y2=1.17
r161 63 67 0.446298 $w=6.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.02 $Y=0.49
+ $X2=1.02 $Y2=0.515
r162 63 64 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.19
+ $Y=0.49 $X2=1.19 $Y2=0.49
r163 57 59 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.78 $Y=1.985
+ $X2=0.78 $Y2=2.815
r164 57 72 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=0.78 $Y=1.985
+ $X2=0.78 $Y2=1.335
r165 47 70 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.19 $Y=1.185
+ $X2=1.19 $Y2=1.17
r166 44 46 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.975 $Y=1.185
+ $X2=4.975 $Y2=0.74
r167 43 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.62 $Y=1.26
+ $X2=4.545 $Y2=1.26
r168 42 44 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.9 $Y=1.26
+ $X2=4.975 $Y2=1.185
r169 42 43 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.9 $Y=1.26
+ $X2=4.62 $Y2=1.26
r170 39 54 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.545 $Y=1.185
+ $X2=4.545 $Y2=1.26
r171 39 41 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.545 $Y=1.185
+ $X2=4.545 $Y2=0.74
r172 38 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.19 $Y=1.26
+ $X2=4.115 $Y2=1.26
r173 37 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.47 $Y=1.26
+ $X2=4.545 $Y2=1.26
r174 37 38 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.47 $Y=1.26
+ $X2=4.19 $Y2=1.26
r175 34 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.115 $Y=1.185
+ $X2=4.115 $Y2=1.26
r176 34 36 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.115 $Y=1.185
+ $X2=4.115 $Y2=0.74
r177 33 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.69 $Y=1.26
+ $X2=3.615 $Y2=1.26
r178 32 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.04 $Y=1.26
+ $X2=4.115 $Y2=1.26
r179 32 33 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.04 $Y=1.26
+ $X2=3.69 $Y2=1.26
r180 29 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.615 $Y=1.185
+ $X2=3.615 $Y2=1.26
r181 29 31 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.615 $Y=1.185
+ $X2=3.615 $Y2=0.74
r182 28 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.26 $Y=1.26
+ $X2=3.185 $Y2=1.26
r183 27 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.54 $Y=1.26
+ $X2=3.615 $Y2=1.26
r184 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.54 $Y=1.26
+ $X2=3.26 $Y2=1.26
r185 24 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.185 $Y=1.185
+ $X2=3.185 $Y2=1.26
r186 24 26 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.185 $Y=1.185
+ $X2=3.185 $Y2=0.74
r187 23 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.76 $Y=1.26
+ $X2=2.685 $Y2=1.26
r188 22 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.11 $Y=1.26
+ $X2=3.185 $Y2=1.26
r189 22 23 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.11 $Y=1.26
+ $X2=2.76 $Y2=1.26
r190 19 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.685 $Y=1.185
+ $X2=2.685 $Y2=1.26
r191 19 21 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.685 $Y=1.185
+ $X2=2.685 $Y2=0.74
r192 18 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.33 $Y=1.26
+ $X2=2.255 $Y2=1.26
r193 17 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.61 $Y=1.26
+ $X2=2.685 $Y2=1.26
r194 17 18 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.61 $Y=1.26
+ $X2=2.33 $Y2=1.26
r195 14 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.255 $Y=1.185
+ $X2=2.255 $Y2=1.26
r196 14 16 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.255 $Y=1.185
+ $X2=2.255 $Y2=0.74
r197 13 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.9 $Y=1.26
+ $X2=1.825 $Y2=1.26
r198 12 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.18 $Y=1.26
+ $X2=2.255 $Y2=1.26
r199 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.18 $Y=1.26
+ $X2=1.9 $Y2=1.26
r200 9 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.825 $Y=1.185
+ $X2=1.825 $Y2=1.26
r201 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.825 $Y=1.185
+ $X2=1.825 $Y2=0.74
r202 8 47 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.355 $Y=1.26
+ $X2=1.19 $Y2=1.185
r203 7 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.75 $Y=1.26
+ $X2=1.825 $Y2=1.26
r204 7 8 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.75 $Y=1.26
+ $X2=1.355 $Y2=1.26
r205 2 59 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.84 $X2=0.78 $Y2=2.815
r206 2 57 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.84 $X2=0.78 $Y2=1.985
r207 1 67 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.63
+ $Y=0.37 $X2=0.77 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__EINVN_8%TE_B 3 5 7 8 10 12 13 15 17 18 20 22 23 25
+ 27 28 30 32 33 35 37 38 40 42 43 45 47 48 49 50 51 52 53 54 55
c168 55 0 1.9459e-20 $X=0.24 $Y=1.295
c169 54 0 1.61579e-19 $X=4.415 $Y=1.67
c170 52 0 1.73215e-20 $X=3.465 $Y=1.67
c171 48 0 1.57621e-19 $X=1.565 $Y=1.67
c172 43 0 1.48702e-19 $X=4.875 $Y=1.65
c173 40 0 5.7999e-20 $X=4.415 $Y=1.765
r174 58 60 17.5187 $w=5.09e-07 $l=1.85e-07 $layer=POLY_cond $X=0.375 $Y=1.465
+ $X2=0.375 $Y2=1.65
r175 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r176 55 59 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.465
r177 45 47 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.965 $Y=1.765
+ $X2=4.965 $Y2=2.4
r178 44 54 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=4.505 $Y=1.65
+ $X2=4.415 $Y2=1.67
r179 43 45 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=4.875 $Y=1.65
+ $X2=4.965 $Y2=1.765
r180 43 44 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.875 $Y=1.65
+ $X2=4.505 $Y2=1.65
r181 40 54 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=4.415 $Y=1.765
+ $X2=4.415 $Y2=1.67
r182 40 42 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.415 $Y=1.765
+ $X2=4.415 $Y2=2.4
r183 39 53 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=4.055 $Y=1.65
+ $X2=3.965 $Y2=1.67
r184 38 54 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=4.325 $Y=1.65
+ $X2=4.415 $Y2=1.67
r185 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.325 $Y=1.65
+ $X2=4.055 $Y2=1.65
r186 35 53 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=3.965 $Y=1.765
+ $X2=3.965 $Y2=1.67
r187 35 37 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.965 $Y=1.765
+ $X2=3.965 $Y2=2.4
r188 34 52 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=3.555 $Y=1.65
+ $X2=3.465 $Y2=1.67
r189 33 53 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=3.875 $Y=1.65
+ $X2=3.965 $Y2=1.67
r190 33 34 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.875 $Y=1.65
+ $X2=3.555 $Y2=1.65
r191 30 52 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=3.465 $Y=1.765
+ $X2=3.465 $Y2=1.67
r192 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.465 $Y=1.765
+ $X2=3.465 $Y2=2.4
r193 29 51 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=3.105 $Y=1.65
+ $X2=3.015 $Y2=1.67
r194 28 52 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=3.375 $Y=1.65
+ $X2=3.465 $Y2=1.67
r195 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.375 $Y=1.65
+ $X2=3.105 $Y2=1.65
r196 25 51 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=3.015 $Y=1.765
+ $X2=3.015 $Y2=1.67
r197 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.015 $Y=1.765
+ $X2=3.015 $Y2=2.4
r198 24 50 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=2.605 $Y=1.65
+ $X2=2.515 $Y2=1.67
r199 23 51 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=2.925 $Y=1.65
+ $X2=3.015 $Y2=1.67
r200 23 24 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.925 $Y=1.65
+ $X2=2.605 $Y2=1.65
r201 20 50 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=2.515 $Y=1.765
+ $X2=2.515 $Y2=1.67
r202 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.515 $Y=1.765
+ $X2=2.515 $Y2=2.4
r203 19 49 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=2.155 $Y=1.65
+ $X2=2.065 $Y2=1.67
r204 18 50 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=2.425 $Y=1.65
+ $X2=2.515 $Y2=1.67
r205 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.425 $Y=1.65
+ $X2=2.155 $Y2=1.65
r206 15 49 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=2.065 $Y=1.765
+ $X2=2.065 $Y2=1.67
r207 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.065 $Y=1.765
+ $X2=2.065 $Y2=2.4
r208 14 48 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=1.655 $Y=1.65
+ $X2=1.565 $Y2=1.67
r209 13 49 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=1.975 $Y=1.65
+ $X2=2.065 $Y2=1.67
r210 13 14 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.975 $Y=1.65
+ $X2=1.655 $Y2=1.65
r211 10 48 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=1.565 $Y=1.765
+ $X2=1.565 $Y2=1.67
r212 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.565 $Y=1.765
+ $X2=1.565 $Y2=2.4
r213 9 60 31.8593 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.645 $Y=1.65
+ $X2=0.375 $Y2=1.65
r214 8 48 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=1.475 $Y=1.65
+ $X2=1.565 $Y2=1.67
r215 8 9 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=1.475 $Y=1.65
+ $X2=0.645 $Y2=1.65
r216 5 60 37.4241 $w=5.09e-07 $l=2.30434e-07 $layer=POLY_cond $X=0.555 $Y=1.765
+ $X2=0.375 $Y2=1.65
r217 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.555 $Y=1.765
+ $X2=0.555 $Y2=2.4
r218 1 58 42.1589 $w=5.09e-07 $l=2.49199e-07 $layer=POLY_cond $X=0.555 $Y=1.3
+ $X2=0.375 $Y2=1.465
r219 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.555 $Y=1.3
+ $X2=0.555 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__EINVN_8%A 3 5 7 10 12 14 17 19 21 24 26 28 31 33 35
+ 38 40 42 45 47 49 50 52 55 57 58 59 60 61 87
c159 87 0 1.18608e-19 $X=8.615 $Y=1.557
c160 31 0 1.56455e-19 $X=7.195 $Y=0.74
c161 12 0 1.68675e-19 $X=5.865 $Y=1.765
c162 10 0 1.47232e-19 $X=5.835 $Y=0.74
r163 87 88 1.31694 $w=3.66e-07 $l=1e-08 $layer=POLY_cond $X=8.615 $Y=1.557
+ $X2=8.625 $Y2=1.557
r164 85 87 9.87705 $w=3.66e-07 $l=7.5e-08 $layer=POLY_cond $X=8.54 $Y=1.557
+ $X2=8.615 $Y2=1.557
r165 85 86 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=8.54
+ $Y=1.515 $X2=8.54 $Y2=1.515
r166 83 85 49.3852 $w=3.66e-07 $l=3.75e-07 $layer=POLY_cond $X=8.165 $Y=1.557
+ $X2=8.54 $Y2=1.557
r167 82 83 14.4863 $w=3.66e-07 $l=1.1e-07 $layer=POLY_cond $X=8.055 $Y=1.557
+ $X2=8.165 $Y2=1.557
r168 81 82 44.776 $w=3.66e-07 $l=3.4e-07 $layer=POLY_cond $X=7.715 $Y=1.557
+ $X2=8.055 $Y2=1.557
r169 80 81 11.8525 $w=3.66e-07 $l=9e-08 $layer=POLY_cond $X=7.625 $Y=1.557
+ $X2=7.715 $Y2=1.557
r170 79 80 47.4098 $w=3.66e-07 $l=3.6e-07 $layer=POLY_cond $X=7.265 $Y=1.557
+ $X2=7.625 $Y2=1.557
r171 78 79 9.21858 $w=3.66e-07 $l=7e-08 $layer=POLY_cond $X=7.195 $Y=1.557
+ $X2=7.265 $Y2=1.557
r172 77 78 50.0437 $w=3.66e-07 $l=3.8e-07 $layer=POLY_cond $X=6.815 $Y=1.557
+ $X2=7.195 $Y2=1.557
r173 76 77 15.8033 $w=3.66e-07 $l=1.2e-07 $layer=POLY_cond $X=6.695 $Y=1.557
+ $X2=6.815 $Y2=1.557
r174 75 76 50.0437 $w=3.66e-07 $l=3.8e-07 $layer=POLY_cond $X=6.315 $Y=1.557
+ $X2=6.695 $Y2=1.557
r175 74 75 6.5847 $w=3.66e-07 $l=5e-08 $layer=POLY_cond $X=6.265 $Y=1.557
+ $X2=6.315 $Y2=1.557
r176 72 74 13.8279 $w=3.66e-07 $l=1.05e-07 $layer=POLY_cond $X=6.16 $Y=1.557
+ $X2=6.265 $Y2=1.557
r177 72 73 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=6.16
+ $Y=1.515 $X2=6.16 $Y2=1.515
r178 70 72 38.8497 $w=3.66e-07 $l=2.95e-07 $layer=POLY_cond $X=5.865 $Y=1.557
+ $X2=6.16 $Y2=1.557
r179 69 70 3.95082 $w=3.66e-07 $l=3e-08 $layer=POLY_cond $X=5.835 $Y=1.557
+ $X2=5.865 $Y2=1.557
r180 68 69 55.3115 $w=3.66e-07 $l=4.2e-07 $layer=POLY_cond $X=5.415 $Y=1.557
+ $X2=5.835 $Y2=1.557
r181 67 68 1.31694 $w=3.66e-07 $l=1e-08 $layer=POLY_cond $X=5.405 $Y=1.557
+ $X2=5.415 $Y2=1.557
r182 61 86 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=8.54 $Y2=1.565
r183 60 86 3.75214 $w=4.28e-07 $l=1.4e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.54 $Y2=1.565
r184 59 60 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=8.4 $Y2=1.565
r185 58 59 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.92 $Y2=1.565
r186 57 58 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r187 57 73 21.4408 $w=4.28e-07 $l=8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.16 $Y2=1.565
r188 53 88 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.625 $Y=1.35
+ $X2=8.625 $Y2=1.557
r189 53 55 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.625 $Y=1.35
+ $X2=8.625 $Y2=0.74
r190 50 87 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.615 $Y=1.765
+ $X2=8.615 $Y2=1.557
r191 50 52 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.615 $Y=1.765
+ $X2=8.615 $Y2=2.4
r192 47 83 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.165 $Y=1.765
+ $X2=8.165 $Y2=1.557
r193 47 49 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.165 $Y=1.765
+ $X2=8.165 $Y2=2.4
r194 43 82 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.055 $Y=1.35
+ $X2=8.055 $Y2=1.557
r195 43 45 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.055 $Y=1.35
+ $X2=8.055 $Y2=0.74
r196 40 81 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.715 $Y=1.765
+ $X2=7.715 $Y2=1.557
r197 40 42 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.715 $Y=1.765
+ $X2=7.715 $Y2=2.4
r198 36 80 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.625 $Y=1.35
+ $X2=7.625 $Y2=1.557
r199 36 38 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.625 $Y=1.35
+ $X2=7.625 $Y2=0.74
r200 33 79 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.265 $Y=1.765
+ $X2=7.265 $Y2=1.557
r201 33 35 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.265 $Y=1.765
+ $X2=7.265 $Y2=2.4
r202 29 78 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.195 $Y=1.35
+ $X2=7.195 $Y2=1.557
r203 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.195 $Y=1.35
+ $X2=7.195 $Y2=0.74
r204 26 77 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.815 $Y=1.765
+ $X2=6.815 $Y2=1.557
r205 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.815 $Y=1.765
+ $X2=6.815 $Y2=2.4
r206 22 76 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.695 $Y=1.35
+ $X2=6.695 $Y2=1.557
r207 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.695 $Y=1.35
+ $X2=6.695 $Y2=0.74
r208 19 75 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.315 $Y=1.765
+ $X2=6.315 $Y2=1.557
r209 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.315 $Y=1.765
+ $X2=6.315 $Y2=2.4
r210 15 74 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.265 $Y=1.35
+ $X2=6.265 $Y2=1.557
r211 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.265 $Y=1.35
+ $X2=6.265 $Y2=0.74
r212 12 70 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.865 $Y=1.765
+ $X2=5.865 $Y2=1.557
r213 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.865 $Y=1.765
+ $X2=5.865 $Y2=2.4
r214 8 69 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.835 $Y=1.35
+ $X2=5.835 $Y2=1.557
r215 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.835 $Y=1.35
+ $X2=5.835 $Y2=0.74
r216 5 68 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.415 $Y=1.765
+ $X2=5.415 $Y2=1.557
r217 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.415 $Y=1.765
+ $X2=5.415 $Y2=2.4
r218 1 67 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.405 $Y=1.35
+ $X2=5.405 $Y2=1.557
r219 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.405 $Y=1.35
+ $X2=5.405 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__EINVN_8%VPWR 1 2 3 4 5 16 18 24 28 32 36 40 44 48 50
+ 52 62 63 69 72 75 78
r106 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r107 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r108 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r109 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r110 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r111 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r112 62 63 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r113 60 63 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=8.88 $Y2=3.33
r114 59 62 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=8.88 $Y2=3.33
r115 59 60 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r116 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=4.69 $Y2=3.33
r117 57 59 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=5.04 $Y2=3.33
r118 56 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r119 56 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r120 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r121 53 66 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r122 53 55 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r123 52 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.625 $Y=3.33
+ $X2=1.79 $Y2=3.33
r124 52 55 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=1.625 $Y=3.33
+ $X2=0.72 $Y2=3.33
r125 50 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r126 50 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.6 $Y2=3.33
r127 50 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r128 46 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.69 $Y=3.245
+ $X2=4.69 $Y2=3.33
r129 46 48 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=4.69 $Y=3.245
+ $X2=4.69 $Y2=2.455
r130 45 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=3.69 $Y2=3.33
r131 44 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=4.69 $Y2=3.33
r132 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=3.855 $Y2=3.33
r133 40 43 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=3.69 $Y=2.09
+ $X2=3.69 $Y2=2.815
r134 38 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=3.245
+ $X2=3.69 $Y2=3.33
r135 38 43 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.69 $Y=3.245
+ $X2=3.69 $Y2=2.815
r136 37 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=3.33
+ $X2=2.74 $Y2=3.33
r137 36 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=3.33
+ $X2=3.69 $Y2=3.33
r138 36 37 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.525 $Y=3.33
+ $X2=2.905 $Y2=3.33
r139 32 35 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=2.74 $Y=2.09
+ $X2=2.74 $Y2=2.815
r140 30 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=3.245
+ $X2=2.74 $Y2=3.33
r141 30 35 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.74 $Y=3.245
+ $X2=2.74 $Y2=2.815
r142 29 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=1.79 $Y2=3.33
r143 28 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=3.33
+ $X2=2.74 $Y2=3.33
r144 28 29 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.575 $Y=3.33
+ $X2=1.955 $Y2=3.33
r145 24 27 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=1.79 $Y=2.09
+ $X2=1.79 $Y2=2.815
r146 22 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=3.245
+ $X2=1.79 $Y2=3.33
r147 22 27 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.79 $Y=3.245
+ $X2=1.79 $Y2=2.815
r148 18 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r149 16 66 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r150 16 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r151 5 48 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=4.49
+ $Y=1.84 $X2=4.69 $Y2=2.455
r152 4 43 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.54
+ $Y=1.84 $X2=3.69 $Y2=2.815
r153 4 40 400 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_PDIFF $count=1 $X=3.54
+ $Y=1.84 $X2=3.69 $Y2=2.09
r154 3 35 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=1.84 $X2=2.74 $Y2=2.815
r155 3 32 400 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=1.84 $X2=2.74 $Y2=2.09
r156 2 27 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.64
+ $Y=1.84 $X2=1.79 $Y2=2.815
r157 2 24 400 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_PDIFF $count=1 $X=1.64
+ $Y=1.84 $X2=1.79 $Y2=2.09
r158 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r159 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__EINVN_8%A_239_368# 1 2 3 4 5 6 7 8 9 30 34 35 38 42
+ 46 50 54 56 58 61 62 63 66 68 72 74 78 80 84 88 89 90 98 99 100
c173 90 0 1.66023e-19 $X=4.26 $Y=1.75
c174 56 0 4.28201e-20 $X=5.025 $Y=2.035
c175 50 0 6.65594e-20 $X=4.025 $Y=1.75
r176 94 95 1.20266 $w=4.68e-07 $l=5e-09 $layer=LI1_cond $X=4.26 $Y=2.115
+ $X2=4.26 $Y2=2.12
r177 92 94 2.03588 $w=4.68e-07 $l=8e-08 $layer=LI1_cond $X=4.26 $Y=2.035
+ $X2=4.26 $Y2=2.115
r178 90 92 7.25282 $w=4.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.26 $Y=1.75
+ $X2=4.26 $Y2=2.035
r179 84 87 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=8.88 $Y=2.115
+ $X2=8.88 $Y2=2.815
r180 82 87 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=8.88 $Y=2.905
+ $X2=8.88 $Y2=2.815
r181 81 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.025 $Y=2.99
+ $X2=7.94 $Y2=2.99
r182 80 82 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.755 $Y=2.99
+ $X2=8.88 $Y2=2.905
r183 80 81 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=8.755 $Y=2.99
+ $X2=8.025 $Y2=2.99
r184 76 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.94 $Y=2.905
+ $X2=7.94 $Y2=2.99
r185 76 78 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=7.94 $Y=2.905
+ $X2=7.94 $Y2=2.455
r186 75 99 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.125 $Y=2.99
+ $X2=7.04 $Y2=2.99
r187 74 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.855 $Y=2.99
+ $X2=7.94 $Y2=2.99
r188 74 75 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.855 $Y=2.99
+ $X2=7.125 $Y2=2.99
r189 70 99 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.04 $Y=2.905
+ $X2=7.04 $Y2=2.99
r190 70 72 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=7.04 $Y=2.905
+ $X2=7.04 $Y2=2.455
r191 69 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=2.99
+ $X2=6.09 $Y2=2.99
r192 68 99 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.955 $Y=2.99
+ $X2=7.04 $Y2=2.99
r193 68 69 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.955 $Y=2.99
+ $X2=6.255 $Y2=2.99
r194 64 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.09 $Y=2.905
+ $X2=6.09 $Y2=2.99
r195 64 66 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.09 $Y=2.905
+ $X2=6.09 $Y2=2.455
r196 62 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.925 $Y=2.99
+ $X2=6.09 $Y2=2.99
r197 62 63 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.925 $Y=2.99
+ $X2=5.355 $Y2=2.99
r198 59 63 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.19 $Y=2.905
+ $X2=5.355 $Y2=2.99
r199 59 61 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.19 $Y=2.905
+ $X2=5.19 $Y2=2.815
r200 58 97 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=2.12 $X2=5.19
+ $Y2=2.035
r201 58 61 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.19 $Y=2.12
+ $X2=5.19 $Y2=2.815
r202 57 92 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=4.495 $Y=2.035
+ $X2=4.26 $Y2=2.035
r203 56 97 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.025 $Y=2.035
+ $X2=5.19 $Y2=2.035
r204 56 57 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.025 $Y=2.035
+ $X2=4.495 $Y2=2.035
r205 54 95 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.19 $Y=2.815
+ $X2=4.19 $Y2=2.12
r206 51 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.325 $Y=1.75
+ $X2=3.2 $Y2=1.75
r207 50 90 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=4.025 $Y=1.75
+ $X2=4.26 $Y2=1.75
r208 50 51 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.025 $Y=1.75
+ $X2=3.325 $Y2=1.75
r209 46 48 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=3.2 $Y=2.115 $X2=3.2
+ $Y2=2.815
r210 44 89 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=1.835
+ $X2=3.2 $Y2=1.75
r211 44 46 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=3.2 $Y=1.835
+ $X2=3.2 $Y2=2.115
r212 43 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.375 $Y=1.75
+ $X2=2.25 $Y2=1.75
r213 42 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.075 $Y=1.75
+ $X2=3.2 $Y2=1.75
r214 42 43 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.075 $Y=1.75
+ $X2=2.375 $Y2=1.75
r215 38 40 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=2.25 $Y=2.115
+ $X2=2.25 $Y2=2.815
r216 36 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.25 $Y=1.835
+ $X2=2.25 $Y2=1.75
r217 36 38 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=2.25 $Y=1.835
+ $X2=2.25 $Y2=2.115
r218 34 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.125 $Y=1.75
+ $X2=2.25 $Y2=1.75
r219 34 35 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.125 $Y=1.75
+ $X2=1.425 $Y2=1.75
r220 30 32 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=1.3 $Y=2.115 $X2=1.3
+ $Y2=2.815
r221 28 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.3 $Y=1.835
+ $X2=1.425 $Y2=1.75
r222 28 30 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=1.3 $Y=1.835
+ $X2=1.3 $Y2=2.115
r223 9 87 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.69
+ $Y=1.84 $X2=8.84 $Y2=2.815
r224 9 84 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=8.69
+ $Y=1.84 $X2=8.84 $Y2=2.115
r225 8 78 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=7.79
+ $Y=1.84 $X2=7.94 $Y2=2.455
r226 7 72 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=6.89
+ $Y=1.84 $X2=7.04 $Y2=2.455
r227 6 66 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=5.94
+ $Y=1.84 $X2=6.09 $Y2=2.455
r228 5 97 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=5.04
+ $Y=1.84 $X2=5.19 $Y2=2.115
r229 5 61 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.04
+ $Y=1.84 $X2=5.19 $Y2=2.815
r230 4 94 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=1.84 $X2=4.19 $Y2=2.115
r231 4 54 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=1.84 $X2=4.19 $Y2=2.815
r232 3 48 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.09
+ $Y=1.84 $X2=3.24 $Y2=2.815
r233 3 46 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.09
+ $Y=1.84 $X2=3.24 $Y2=2.115
r234 2 40 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.14
+ $Y=1.84 $X2=2.29 $Y2=2.815
r235 2 38 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.14
+ $Y=1.84 $X2=2.29 $Y2=2.115
r236 1 32 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=1.195
+ $Y=1.84 $X2=1.34 $Y2=2.815
r237 1 30 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=1.195
+ $Y=1.84 $X2=1.34 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__EINVN_8%Z 1 2 3 4 5 6 7 8 25 26 28 31 35 39 41 43 47
+ 51 53 57 63 64 66 69 70 72 73 75 77 78
c121 70 0 1.47232e-19 $X=6.645 $Y=0.975
c122 64 0 1.68675e-19 $X=5.59 $Y=1.665
c123 63 0 1.53018e-19 $X=5.455 $Y=1.665
c124 26 0 1.1822e-19 $X=5.59 $Y=1.55
r125 68 70 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.48 $Y=0.975
+ $X2=6.645 $Y2=0.975
r126 68 69 4.83878 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.48 $Y=0.975
+ $X2=6.315 $Y2=0.975
r127 63 78 20.7941 $w=2.28e-07 $l=4.15e-07 $layer=LI1_cond $X=5.455 $Y=1.665
+ $X2=5.04 $Y2=1.665
r128 63 64 1.18299 $w=2.3e-07 $l=1.35e-07 $layer=LI1_cond $X=5.455 $Y=1.665
+ $X2=5.59 $Y2=1.665
r129 55 57 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=8.34 $Y=1.01
+ $X2=8.34 $Y2=0.78
r130 54 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.655 $Y=2.035
+ $X2=7.49 $Y2=2.035
r131 53 77 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.225 $Y=2.035
+ $X2=8.39 $Y2=2.035
r132 53 54 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.225 $Y=2.035
+ $X2=7.655 $Y2=2.035
r133 52 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.495 $Y=1.095
+ $X2=7.41 $Y2=1.095
r134 51 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.175 $Y=1.095
+ $X2=8.34 $Y2=1.01
r135 51 52 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.175 $Y=1.095
+ $X2=7.495 $Y2=1.095
r136 45 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.41 $Y=1.01
+ $X2=7.41 $Y2=1.095
r137 45 47 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.41 $Y=1.01
+ $X2=7.41 $Y2=0.78
r138 44 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.755 $Y=2.035
+ $X2=6.59 $Y2=2.035
r139 43 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.325 $Y=2.035
+ $X2=7.49 $Y2=2.035
r140 43 44 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.325 $Y=2.035
+ $X2=6.755 $Y2=2.035
r141 41 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.325 $Y=1.095
+ $X2=7.41 $Y2=1.095
r142 41 70 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.325 $Y=1.095
+ $X2=6.645 $Y2=1.095
r143 37 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.59 $Y=2.12
+ $X2=6.59 $Y2=2.035
r144 37 39 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=6.59 $Y=2.12
+ $X2=6.59 $Y2=2.615
r145 36 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.725 $Y=2.035
+ $X2=5.64 $Y2=2.035
r146 35 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.425 $Y=2.035
+ $X2=6.59 $Y2=2.035
r147 35 36 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.425 $Y=2.035
+ $X2=5.725 $Y2=2.035
r148 34 62 2.99957 $w=3.6e-07 $l=1.35e-07 $layer=LI1_cond $X=5.725 $Y=0.95
+ $X2=5.59 $Y2=0.95
r149 34 69 18.8873 $w=3.58e-07 $l=5.9e-07 $layer=LI1_cond $X=5.725 $Y=0.95
+ $X2=6.315 $Y2=0.95
r150 29 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.64 $Y=2.12
+ $X2=5.64 $Y2=2.035
r151 29 31 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.64 $Y=2.12
+ $X2=5.64 $Y2=2.57
r152 28 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.64 $Y=1.95
+ $X2=5.64 $Y2=2.035
r153 27 64 5.35987 $w=2.2e-07 $l=1.3775e-07 $layer=LI1_cond $X=5.64 $Y=1.78
+ $X2=5.59 $Y2=1.665
r154 27 28 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.64 $Y=1.78
+ $X2=5.64 $Y2=1.95
r155 26 64 5.35987 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=5.59 $Y=1.55
+ $X2=5.59 $Y2=1.665
r156 25 62 3.99943 $w=2.7e-07 $l=1.8e-07 $layer=LI1_cond $X=5.59 $Y=1.13
+ $X2=5.59 $Y2=0.95
r157 25 26 17.9269 $w=2.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.59 $Y=1.13
+ $X2=5.59 $Y2=1.55
r158 8 77 300 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=2 $X=8.24
+ $Y=1.84 $X2=8.39 $Y2=2.035
r159 7 75 300 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=2 $X=7.34
+ $Y=1.84 $X2=7.49 $Y2=2.035
r160 6 72 600 $w=1.7e-07 $l=2.81069e-07 $layer=licon1_PDIFF $count=1 $X=6.39
+ $Y=1.84 $X2=6.59 $Y2=2.035
r161 6 39 600 $w=1.7e-07 $l=8.69267e-07 $layer=licon1_PDIFF $count=1 $X=6.39
+ $Y=1.84 $X2=6.59 $Y2=2.615
r162 5 66 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.49
+ $Y=1.84 $X2=5.64 $Y2=1.985
r163 5 31 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=5.49
+ $Y=1.84 $X2=5.64 $Y2=2.57
r164 4 57 182 $w=1.7e-07 $l=5.04182e-07 $layer=licon1_NDIFF $count=1 $X=8.13
+ $Y=0.37 $X2=8.34 $Y2=0.78
r165 3 47 182 $w=1.7e-07 $l=4.74868e-07 $layer=licon1_NDIFF $count=1 $X=7.27
+ $Y=0.37 $X2=7.41 $Y2=0.78
r166 2 68 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=6.34
+ $Y=0.37 $X2=6.48 $Y2=0.91
r167 1 62 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.48
+ $Y=0.37 $X2=5.62 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LS__EINVN_8%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 43 44 46 47 48 70 71
c108 71 0 3.46022e-20 $X=8.88 $Y=0
r109 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r110 70 71 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r111 68 71 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=8.88
+ $Y2=0
r112 67 70 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=8.88
+ $Y2=0
r113 67 68 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r114 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r115 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r116 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r117 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r118 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r119 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r120 53 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r121 52 55 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r122 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r123 50 74 4.61231 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=0.505 $Y=0
+ $X2=0.252 $Y2=0
r124 50 52 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.505 $Y=0
+ $X2=0.72 $Y2=0
r125 48 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r126 48 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r127 48 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r128 46 64 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.595 $Y=0 $X2=4.56
+ $Y2=0
r129 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.595 $Y=0 $X2=4.76
+ $Y2=0
r130 45 67 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.925 $Y=0
+ $X2=5.04 $Y2=0
r131 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.925 $Y=0 $X2=4.76
+ $Y2=0
r132 43 61 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.6
+ $Y2=0
r133 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.83
+ $Y2=0
r134 42 64 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=4.56
+ $Y2=0
r135 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=3.83
+ $Y2=0
r136 40 58 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.64
+ $Y2=0
r137 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.9
+ $Y2=0
r138 39 61 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.065 $Y=0 $X2=3.6
+ $Y2=0
r139 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.065 $Y=0 $X2=2.9
+ $Y2=0
r140 37 55 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.68 $Y2=0
r141 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2
+ $Y2=0
r142 36 58 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.125 $Y=0
+ $X2=2.64 $Y2=0
r143 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=2
+ $Y2=0
r144 32 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.76 $Y=0.085
+ $X2=4.76 $Y2=0
r145 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.76 $Y=0.085
+ $X2=4.76 $Y2=0.515
r146 28 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.83 $Y=0.085
+ $X2=3.83 $Y2=0
r147 28 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.83 $Y=0.085
+ $X2=3.83 $Y2=0.515
r148 24 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=0.085 $X2=2.9
+ $Y2=0
r149 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.9 $Y=0.085
+ $X2=2.9 $Y2=0.515
r150 20 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0
r151 20 22 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0.515
r152 16 74 3.15387 $w=3.3e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.34 $Y=0.085
+ $X2=0.252 $Y2=0
r153 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.34 $Y=0.085
+ $X2=0.34 $Y2=0.515
r154 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.62
+ $Y=0.37 $X2=4.76 $Y2=0.515
r155 4 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.69
+ $Y=0.37 $X2=3.83 $Y2=0.515
r156 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.76
+ $Y=0.37 $X2=2.9 $Y2=0.515
r157 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.9
+ $Y=0.37 $X2=2.04 $Y2=0.515
r158 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.195
+ $Y=0.37 $X2=0.34 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__EINVN_8%A_293_74# 1 2 3 4 5 6 7 8 9 30 32 33 36 38
+ 42 44 48 50 52 55 56 60 64 66 70 72 73 74 77 83
c165 70 0 1.18608e-19 $X=8.84 $Y=0.515
c166 56 0 1.56455e-19 $X=6.815 $Y=0.427
r167 79 81 8.13695 $w=3.28e-07 $l=2.33e-07 $layer=LI1_cond $X=6.98 $Y=0.427
+ $X2=6.98 $Y2=0.66
r168 77 79 3.03826 $w=3.28e-07 $l=8.7e-08 $layer=LI1_cond $X=6.98 $Y=0.34
+ $X2=6.98 $Y2=0.427
r169 68 70 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=8.84 $Y=0.425
+ $X2=8.84 $Y2=0.515
r170 67 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.005 $Y=0.34
+ $X2=7.84 $Y2=0.34
r171 66 68 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.675 $Y=0.34
+ $X2=8.84 $Y2=0.425
r172 66 67 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.675 $Y=0.34
+ $X2=8.005 $Y2=0.34
r173 62 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.84 $Y=0.425
+ $X2=7.84 $Y2=0.34
r174 62 64 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=7.84 $Y=0.425
+ $X2=7.84 $Y2=0.66
r175 61 77 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.145 $Y=0.34
+ $X2=6.98 $Y2=0.34
r176 60 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.675 $Y=0.34
+ $X2=7.84 $Y2=0.34
r177 60 61 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.675 $Y=0.34
+ $X2=7.145 $Y2=0.34
r178 57 76 2.60071 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.275 $Y=0.427
+ $X2=5.19 $Y2=0.427
r179 57 59 25.8882 $w=3.43e-07 $l=7.75e-07 $layer=LI1_cond $X=5.275 $Y=0.427
+ $X2=6.05 $Y2=0.427
r180 56 79 0.462083 $w=3.45e-07 $l=1.65e-07 $layer=LI1_cond $X=6.815 $Y=0.427
+ $X2=6.98 $Y2=0.427
r181 56 59 25.5542 $w=3.43e-07 $l=7.65e-07 $layer=LI1_cond $X=6.815 $Y=0.427
+ $X2=6.05 $Y2=0.427
r182 53 55 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.19 $Y=1.21
+ $X2=5.19 $Y2=0.965
r183 52 76 5.29321 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=5.19 $Y=0.6
+ $X2=5.19 $Y2=0.427
r184 52 55 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.19 $Y=0.6
+ $X2=5.19 $Y2=0.965
r185 51 74 7.02821 $w=1.7e-07 $l=1.45774e-07 $layer=LI1_cond $X=4.415 $Y=1.295
+ $X2=4.29 $Y2=1.34
r186 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.105 $Y=1.295
+ $X2=5.19 $Y2=1.21
r187 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.105 $Y=1.295
+ $X2=4.415 $Y2=1.295
r188 46 74 0.00168595 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=4.29 $Y=1.21
+ $X2=4.29 $Y2=1.34
r189 46 48 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=4.29 $Y=1.21
+ $X2=4.29 $Y2=0.515
r190 45 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.485 $Y=1.385
+ $X2=3.36 $Y2=1.385
r191 44 74 7.02821 $w=1.7e-07 $l=1.45774e-07 $layer=LI1_cond $X=4.165 $Y=1.385
+ $X2=4.29 $Y2=1.34
r192 44 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.165 $Y=1.385
+ $X2=3.485 $Y2=1.385
r193 40 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=1.3
+ $X2=3.36 $Y2=1.385
r194 40 42 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=3.36 $Y=1.3
+ $X2=3.36 $Y2=0.515
r195 39 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.555 $Y=1.385
+ $X2=2.43 $Y2=1.385
r196 38 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.235 $Y=1.385
+ $X2=3.36 $Y2=1.385
r197 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.235 $Y=1.385
+ $X2=2.555 $Y2=1.385
r198 34 72 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=1.3
+ $X2=2.43 $Y2=1.385
r199 34 36 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=2.43 $Y=1.3
+ $X2=2.43 $Y2=0.515
r200 32 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.305 $Y=1.385
+ $X2=2.43 $Y2=1.385
r201 32 33 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.305 $Y=1.385
+ $X2=1.695 $Y2=1.385
r202 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.61 $Y=1.3
+ $X2=1.695 $Y2=1.385
r203 28 30 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.61 $Y=1.3
+ $X2=1.61 $Y2=0.515
r204 9 70 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.37 $X2=8.84 $Y2=0.515
r205 8 64 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=7.7
+ $Y=0.37 $X2=7.84 $Y2=0.66
r206 7 81 182 $w=1.7e-07 $l=3.80789e-07 $layer=licon1_NDIFF $count=1 $X=6.77
+ $Y=0.37 $X2=6.98 $Y2=0.66
r207 6 59 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.91
+ $Y=0.37 $X2=6.05 $Y2=0.515
r208 5 76 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.05
+ $Y=0.37 $X2=5.19 $Y2=0.515
r209 5 55 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.05
+ $Y=0.37 $X2=5.19 $Y2=0.965
r210 4 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.19
+ $Y=0.37 $X2=4.33 $Y2=0.515
r211 3 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.26
+ $Y=0.37 $X2=3.4 $Y2=0.515
r212 2 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.33
+ $Y=0.37 $X2=2.47 $Y2=0.515
r213 1 30 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.465
+ $Y=0.37 $X2=1.61 $Y2=0.515
.ends

