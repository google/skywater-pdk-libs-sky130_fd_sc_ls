* File: sky130_fd_sc_ls__dfxtp_2.spice
* Created: Fri Aug 28 13:16:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dfxtp_2.pex.spice"
.subckt sky130_fd_sc_ls__dfxtp_2  VNB VPB CLK D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1022 N_VGND_M1022_d N_CLK_M1022_g N_A_27_74#_M1022_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1628 AS=0.2109 PD=1.18 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1023 N_A_206_368#_M1023_d N_A_27_74#_M1023_g N_VGND_M1022_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2775 AS=0.1628 PD=2.23 PS=1.18 NRD=14.592 NRS=25.944 M=1 R=4.93333
+ SA=75000.8 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1009 N_A_431_508#_M1009_d N_D_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.318675 PD=0.7 PS=2.49 NRD=0 NRS=201.06 M=1 R=2.8 SA=75000.5
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1012 N_A_538_429#_M1012_d N_A_27_74#_M1012_g N_A_431_508#_M1009_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.076125 AS=0.0588 PD=0.835 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1010 A_708_101# N_A_206_368#_M1010_g N_A_538_429#_M1012_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.076125 PD=0.66 PS=0.835 NRD=18.564 NRS=7.14 M=1 R=2.8
+ SA=75001.1 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_A_695_459#_M1025_g A_708_101# VNB NSHORT L=0.15 W=0.42
+ AD=0.180816 AS=0.0504 PD=1.2167 PS=0.66 NRD=107.28 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_695_459#_M1002_d N_A_538_429#_M1002_g N_VGND_M1025_d VNB NSHORT
+ L=0.15 W=0.55 AD=0.077 AS=0.236784 PD=0.83 PS=1.5933 NRD=0 NRS=73.08 M=1
+ R=3.66667 SA=75001.9 SB=75001.2 A=0.0825 P=1.4 MULT=1
MM1005 N_A_1019_424#_M1005_d N_A_206_368#_M1005_g N_A_695_459#_M1002_d VNB
+ NSHORT L=0.15 W=0.55 AD=0.139229 AS=0.077 PD=1.33247 PS=0.83 NRD=32.724 NRS=0
+ M=1 R=3.66667 SA=75002.4 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1013 A_1172_124# N_A_27_74#_M1013_g N_A_1019_424#_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.106321 PD=0.66 PS=1.01753 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75002.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_1217_314#_M1001_g A_1172_124# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75003.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_1019_424#_M1014_g N_A_1217_314#_M1014_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.11405 AS=0.15675 PD=0.972093 PS=1.67 NRD=5.448 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75001.2 A=0.0825 P=1.4 MULT=1
MM1004 N_Q_M1004_d N_A_1217_314#_M1004_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.15345 PD=1.02 PS=1.30791 NRD=0 NRS=15.396 M=1 R=4.93333
+ SA=75000.6 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1015 N_Q_M1004_d N_A_1217_314#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_VPWR_M1016_d N_CLK_M1016_g N_A_27_74#_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1017 N_A_206_368#_M1017_d N_A_27_74#_M1017_g N_VPWR_M1016_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1020 N_A_431_508#_M1020_d N_D_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.115412 AS=0.2474 PD=1.2 PS=2.13 NRD=103.09 NRS=250.486 M=1 R=2.8
+ SA=75000.3 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1006 N_A_538_429#_M1006_d N_A_206_368#_M1006_g N_A_431_508#_M1020_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.112612 AS=0.115412 PD=1.175 PS=1.2 NRD=4.6886
+ NRS=4.6886 M=1 R=2.8 SA=75000.3 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1003 A_644_504# N_A_27_74#_M1003_g N_A_538_429#_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.112612 PD=0.69 PS=1.175 NRD=37.5088 NRS=99.9578 M=1
+ R=2.8 SA=75000.3 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1018 N_VPWR_M1018_d N_A_695_459#_M1018_g A_644_504# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.139883 AS=0.0567 PD=1.07 PS=0.69 NRD=130.414 NRS=37.5088 M=1 R=2.8
+ SA=75000.7 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1011 N_A_695_459#_M1011_d N_A_538_429#_M1011_g N_VPWR_M1018_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2625 AS=0.279767 PD=1.465 PS=2.14 NRD=3.5066 NRS=65.207 M=1
+ R=5.6 SA=75000.8 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1024 N_A_1019_424#_M1024_d N_A_27_74#_M1024_g N_A_695_459#_M1011_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1876 AS=0.2625 PD=1.62667 PS=1.465 NRD=2.3443 NRS=77.3816
+ M=1 R=5.6 SA=75001.6 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1007 A_1125_508# N_A_206_368#_M1007_g N_A_1019_424#_M1024_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.09975 AS=0.0938 PD=0.895 PS=0.813333 NRD=85.5965 NRS=44.5417 M=1
+ R=2.8 SA=75002.6 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_1217_314#_M1008_g A_1125_508# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1218 AS=0.09975 PD=1.42 PS=0.895 NRD=4.6886 NRS=85.5965 M=1 R=2.8
+ SA=75003.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_VPWR_M1019_d N_A_1019_424#_M1019_g N_A_1217_314#_M1019_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.182453 AS=0.295 PD=1.39151 PS=2.59 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1019_d N_A_1217_314#_M1000_g N_Q_M1000_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.204347 AS=0.168 PD=1.55849 PS=1.42 NRD=11.426 NRS=1.7533 M=1
+ R=7.46667 SA=75000.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1021 N_VPWR_M1021_d N_A_1217_314#_M1021_g N_Q_M1000_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX26_noxref VNB VPB NWDIODE A=16.7772 P=21.76
c_1509 A_708_101# 0 4.2343e-20 $X=3.54 $Y=0.505
*
.include "sky130_fd_sc_ls__dfxtp_2.pxi.spice"
*
.ends
*
*
