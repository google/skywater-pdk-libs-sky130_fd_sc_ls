* NGSPICE file created from sky130_fd_sc_ls__buf_16.ext - technology: sky130A

.subckt sky130_fd_sc_ls__buf_16 A VGND VNB VPB VPWR X
M1000 X a_83_260# VGND VNB nshort w=740000u l=150000u
+  ad=1.6576e+12p pd=1.632e+07u as=2.8305e+12p ps=2.541e+07u
M1001 VPWR a_83_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=4.1328e+12p pd=3.426e+07u as=2.688e+12p ps=2.272e+07u
M1002 VPWR A a_83_260# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=1.008e+12p ps=8.52e+06u
M1003 VPWR A a_83_260# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_83_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A a_83_260# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=6.734e+11p ps=6.26e+06u
M1006 X a_83_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_83_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_83_260# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_83_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_83_260# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_83_260# A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_83_260# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_83_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_83_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_83_260# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A a_83_260# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A a_83_260# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_83_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_83_260# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_83_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_83_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_83_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_83_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_83_260# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 X a_83_260# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_83_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_83_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_83_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR A a_83_260# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 X a_83_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_83_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 X a_83_260# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND a_83_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 X a_83_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_83_260# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND a_83_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_83_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 X a_83_260# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND a_83_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_83_260# A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR a_83_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 X a_83_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_83_260# A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

