* File: sky130_fd_sc_ls__or4bb_2.pex.spice
* Created: Wed Sep  2 11:26:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__OR4BB_2%D_N 1 2 3 5 6 8 9 13
c32 6 0 1.19082e-19 $X=0.5 $Y=1.35
r33 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.515 $X2=0.385 $Y2=1.515
r34 9 13 4.06745 $w=4.23e-07 $l=1.5e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.515
r35 6 12 38.5406 $w=3.17e-07 $l=2.08315e-07 $layer=POLY_cond $X=0.5 $Y=1.35
+ $X2=0.402 $Y2=1.515
r36 6 8 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.5 $Y=1.35 $X2=0.5
+ $Y2=0.965
r37 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=2.045
+ $X2=0.495 $Y2=2.54
r38 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.495 $Y=1.955 $X2=0.495
+ $Y2=2.045
r39 1 12 47.701 $w=3.17e-07 $l=2.97893e-07 $layer=POLY_cond $X=0.495 $Y=1.77
+ $X2=0.402 $Y2=1.515
r40 1 2 71.9113 $w=1.8e-07 $l=1.85e-07 $layer=POLY_cond $X=0.495 $Y=1.77
+ $X2=0.495 $Y2=1.955
.ends

.subckt PM_SKY130_FD_SC_LS__OR4BB_2%A_182_270# 1 2 3 10 12 15 16 17 18 20 21 23
+ 25 26 30 35 36 38 43 45 47
c119 36 0 2.10213e-20 $X=3.405 $Y=1.215
r120 47 49 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=3.57 $Y=1.07
+ $X2=3.57 $Y2=1.215
r121 41 51 6.98973 $w=3.31e-07 $l=4.8e-08 $layer=POLY_cond $X=1.545 $Y=1.515
+ $X2=1.545 $Y2=1.467
r122 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=1.515 $X2=1.565 $Y2=1.515
r123 38 40 13.7594 $w=2.66e-07 $l=3e-07 $layer=LI1_cond $X=1.565 $Y=1.215
+ $X2=1.565 $Y2=1.515
r124 37 45 4.30018 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=1.215
+ $X2=2.475 $Y2=1.215
r125 36 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=1.215
+ $X2=3.57 $Y2=1.215
r126 36 37 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=3.405 $Y=1.215
+ $X2=2.64 $Y2=1.215
r127 35 43 12.9201 $w=2.88e-07 $l=3.86588e-07 $layer=LI1_cond $X=2.52 $Y=2.61
+ $X2=2.215 $Y2=2.795
r128 34 45 1.96316 $w=1.7e-07 $l=1.05119e-07 $layer=LI1_cond $X=2.52 $Y=1.3
+ $X2=2.475 $Y2=1.215
r129 34 35 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=2.52 $Y=1.3
+ $X2=2.52 $Y2=2.61
r130 30 33 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=2.475 $Y=0.745
+ $X2=2.475 $Y2=1.095
r131 28 45 1.96316 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=1.13
+ $X2=2.475 $Y2=1.215
r132 28 33 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.475 $Y=1.13
+ $X2=2.475 $Y2=1.095
r133 27 38 3.35683 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.73 $Y=1.215
+ $X2=1.565 $Y2=1.215
r134 26 45 4.30018 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=1.215
+ $X2=2.475 $Y2=1.215
r135 26 27 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.31 $Y=1.215
+ $X2=1.73 $Y2=1.215
r136 21 41 50.9845 $w=3.31e-07 $l=2.93684e-07 $layer=POLY_cond $X=1.45 $Y=1.765
+ $X2=1.545 $Y2=1.515
r137 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.45 $Y=1.765
+ $X2=1.45 $Y2=2.4
r138 18 51 31.6172 $w=3.31e-07 $l=1.59339e-07 $layer=POLY_cond $X=1.445 $Y=1.35
+ $X2=1.545 $Y2=1.467
r139 18 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.445 $Y=1.35
+ $X2=1.445 $Y2=0.87
r140 17 25 47.6288 $w=1.8e-07 $l=1.17e-07 $layer=POLY_cond $X=1 $Y=1.467 $X2=1
+ $Y2=1.35
r141 16 51 10.9133 $w=2.35e-07 $l=1.85e-07 $layer=POLY_cond $X=1.36 $Y=1.467
+ $X2=1.545 $Y2=1.467
r142 16 17 71.3643 $w=2.35e-07 $l=2.7e-07 $layer=POLY_cond $X=1.36 $Y=1.467
+ $X2=1.09 $Y2=1.467
r143 15 25 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.015 $Y=0.87
+ $X2=1.015 $Y2=1.35
r144 10 17 117.985 $w=1.8e-07 $l=2.98e-07 $layer=POLY_cond $X=1 $Y=1.765 $X2=1
+ $Y2=1.467
r145 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1 $Y=1.765 $X2=1
+ $Y2=2.4
r146 3 43 600 $w=1.7e-07 $l=8.99972e-07 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.96 $X2=2.215 $Y2=2.795
r147 2 47 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=3.43
+ $Y=0.68 $X2=3.57 $Y2=1.07
r148 1 33 182 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_NDIFF $count=1 $X=2.255
+ $Y=0.6 $X2=2.475 $Y2=1.095
r149 1 30 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=2.255
+ $Y=0.6 $X2=2.475 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LS__OR4BB_2%A_27_424# 1 2 9 11 13 18 20 21 23 24 28 32
+ 35 37
r88 37 38 35.1036 $w=3.57e-07 $l=2.6e-07 $layer=POLY_cond $X=2.18 $Y=1.677
+ $X2=2.44 $Y2=1.677
r89 34 35 5.76029 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=2.27
+ $X2=0.89 $Y2=2.27
r90 32 34 18.134 $w=3.38e-07 $l=5.35e-07 $layer=LI1_cond $X=0.27 $Y=2.27
+ $X2=0.805 $Y2=2.27
r91 29 37 6.07563 $w=3.57e-07 $l=4.5e-08 $layer=POLY_cond $X=2.135 $Y=1.677
+ $X2=2.18 $Y2=1.677
r92 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.135
+ $Y=1.635 $X2=2.135 $Y2=1.635
r93 26 28 24.8068 $w=2.93e-07 $l=6.35e-07 $layer=LI1_cond $X=2.117 $Y=2.27
+ $X2=2.117 $Y2=1.635
r94 24 26 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=1.97 $Y=2.355
+ $X2=2.117 $Y2=2.27
r95 24 35 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=1.97 $Y=2.355
+ $X2=0.89 $Y2=2.355
r96 23 34 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.805 $Y=2.1
+ $X2=0.805 $Y2=2.27
r97 22 23 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.805 $Y=1.18
+ $X2=0.805 $Y2=2.1
r98 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.72 $Y=1.095
+ $X2=0.805 $Y2=1.18
r99 20 21 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.72 $Y=1.095
+ $X2=0.45 $Y2=1.095
r100 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.285 $Y=1.01
+ $X2=0.45 $Y2=1.095
r101 16 18 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=1.01
+ $X2=0.285 $Y2=0.925
r102 11 38 23.1043 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.44 $Y=1.885
+ $X2=2.44 $Y2=1.677
r103 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.44 $Y=1.885
+ $X2=2.44 $Y2=2.46
r104 7 37 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.18 $Y=1.47
+ $X2=2.18 $Y2=1.677
r105 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.18 $Y=1.47 $X2=2.18
+ $Y2=0.92
r106 2 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.27 $Y2=2.265
r107 1 18 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.69 $X2=0.285 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LS__OR4BB_2%A_548_110# 1 2 9 11 13 16 20 22 25 27 34 36
c76 16 0 1.16141e-19 $X=2.905 $Y=1.635
c77 9 0 2.06399e-20 $X=2.815 $Y=1
r78 33 36 20.1388 $w=1.88e-07 $l=3.45e-07 $layer=LI1_cond $X=4.18 $Y=2.045
+ $X2=4.525 $Y2=2.045
r79 33 34 5.10991 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=4.18 $Y=2.045
+ $X2=4.095 $Y2=2.045
r80 25 29 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.56 $Y=1.045
+ $X2=4.18 $Y2=1.045
r81 25 27 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=4.56 $Y=0.96
+ $X2=4.56 $Y2=0.73
r82 22 33 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.18 $Y=1.95 $X2=4.18
+ $Y2=2.045
r83 21 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.18 $Y=1.13
+ $X2=4.18 $Y2=1.045
r84 21 22 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=4.18 $Y=1.13
+ $X2=4.18 $Y2=1.95
r85 20 34 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=3.07 $Y=2.055
+ $X2=4.095 $Y2=2.055
r86 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.905
+ $Y=1.635 $X2=2.905 $Y2=1.635
r87 14 20 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=2.922 $Y=1.97
+ $X2=3.07 $Y2=2.055
r88 14 16 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=2.922 $Y=1.97
+ $X2=2.922 $Y2=1.635
r89 11 17 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.86 $Y=1.885
+ $X2=2.905 $Y2=1.635
r90 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.86 $Y=1.885
+ $X2=2.86 $Y2=2.46
r91 7 17 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.815 $Y=1.47
+ $X2=2.905 $Y2=1.635
r92 7 9 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.815 $Y=1.47 $X2=2.815
+ $Y2=1
r93 2 36 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=4.375
+ $Y=1.96 $X2=4.525 $Y2=2.115
r94 1 27 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.38
+ $Y=0.455 $X2=4.52 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_LS__OR4BB_2%B 4 5 6 7 9 14 16 22
c45 22 0 2.06399e-20 $X=3.485 $Y=0.462
r46 16 22 3.89033 $w=4.13e-07 $l=1.15e-07 $layer=LI1_cond $X=3.6 $Y=0.462
+ $X2=3.485 $Y2=0.462
r47 14 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.315 $Y=0.405
+ $X2=3.315 $Y2=0.57
r48 13 22 6.21953 $w=3.13e-07 $l=1.7e-07 $layer=LI1_cond $X=3.315 $Y=0.412
+ $X2=3.485 $Y2=0.412
r49 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.315
+ $Y=0.405 $X2=3.315 $Y2=0.405
r50 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.37 $Y=1.885
+ $X2=3.37 $Y2=2.46
r51 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.37 $Y=1.795 $X2=3.37
+ $Y2=1.885
r52 5 10 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.37 $Y=1.485 $X2=3.37
+ $Y2=1.395
r53 5 6 120.5 $w=1.8e-07 $l=3.1e-07 $layer=POLY_cond $X=3.37 $Y=1.485 $X2=3.37
+ $Y2=1.795
r54 4 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.355 $Y=1 $X2=3.355
+ $Y2=1.395
r55 4 20 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.355 $Y=1 $X2=3.355
+ $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LS__OR4BB_2%A 1 3 6 8 12
c34 6 0 2.10213e-20 $X=3.795 $Y=1
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.835
+ $Y=1.635 $X2=3.835 $Y2=1.635
r36 8 12 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=3.6 $Y=1.635
+ $X2=3.835 $Y2=1.635
r37 4 11 38.5562 $w=2.99e-07 $l=1.83916e-07 $layer=POLY_cond $X=3.795 $Y=1.47
+ $X2=3.835 $Y2=1.635
r38 4 6 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.795 $Y=1.47 $X2=3.795
+ $Y2=1
r39 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=3.76 $Y=1.885
+ $X2=3.835 $Y2=1.635
r40 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.76 $Y=1.885
+ $X2=3.76 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__OR4BB_2%C_N 2 3 5 8 10 16 17
r32 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.53
+ $Y=1.465 $X2=4.53 $Y2=1.465
r33 14 16 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=4.305 $Y=1.465
+ $X2=4.53 $Y2=1.465
r34 12 14 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=4.3 $Y=1.465
+ $X2=4.305 $Y2=1.465
r35 10 17 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=4.565 $Y=1.665
+ $X2=4.565 $Y2=1.465
r36 6 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.3
+ $X2=4.305 $Y2=1.465
r37 6 8 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=4.305 $Y=1.3 $X2=4.305
+ $Y2=0.73
r38 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.3 $Y=1.885 $X2=4.3
+ $Y2=2.38
r39 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.3 $Y=1.795 $X2=4.3
+ $Y2=1.885
r40 1 12 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.3 $Y=1.63 $X2=4.3
+ $Y2=1.465
r41 1 2 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.3 $Y=1.63 $X2=4.3
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__OR4BB_2%VPWR 1 2 3 12 16 20 25 26 27 29 34 47 48 51
+ 54
r54 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r57 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r58 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r59 42 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 41 44 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r61 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r62 39 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.84 $Y=3.33
+ $X2=1.675 $Y2=3.33
r63 39 41 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.84 $Y=3.33 $X2=2.16
+ $Y2=3.33
r64 38 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r67 35 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=0.77 $Y2=3.33
r68 35 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=1.2 $Y2=3.33
r69 34 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.51 $Y=3.33
+ $X2=1.675 $Y2=3.33
r70 34 37 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.51 $Y=3.33 $X2=1.2
+ $Y2=3.33
r71 32 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r73 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.77 $Y2=3.33
r74 29 31 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.24 $Y2=3.33
r75 27 45 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r76 27 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r77 25 44 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.82 $Y=3.33 $X2=3.6
+ $Y2=3.33
r78 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.82 $Y=3.33
+ $X2=3.985 $Y2=3.33
r79 24 47 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=4.15 $Y=3.33
+ $X2=4.56 $Y2=3.33
r80 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.15 $Y=3.33
+ $X2=3.985 $Y2=3.33
r81 20 23 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.985 $Y=2.395
+ $X2=3.985 $Y2=2.795
r82 18 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.985 $Y=3.245
+ $X2=3.985 $Y2=3.33
r83 18 23 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.985 $Y=3.245
+ $X2=3.985 $Y2=2.795
r84 14 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.675 $Y=3.245
+ $X2=1.675 $Y2=3.33
r85 14 16 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.675 $Y=3.245
+ $X2=1.675 $Y2=2.795
r86 10 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=3.245
+ $X2=0.77 $Y2=3.33
r87 10 12 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.77 $Y=3.245
+ $X2=0.77 $Y2=2.795
r88 3 23 600 $w=1.7e-07 $l=9.06904e-07 $layer=licon1_PDIFF $count=1 $X=3.835
+ $Y=1.96 $X2=3.985 $Y2=2.795
r89 3 20 600 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_PDIFF $count=1 $X=3.835
+ $Y=1.96 $X2=3.985 $Y2=2.395
r90 2 16 600 $w=1.7e-07 $l=1.02727e-06 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.84 $X2=1.675 $Y2=2.795
r91 1 12 600 $w=1.7e-07 $l=7.68521e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=2.12 $X2=0.77 $Y2=2.795
.ends

.subckt PM_SKY130_FD_SC_LS__OR4BB_2%X 1 2 10 12 13 15 16
c27 10 0 1.19082e-19 $X=1.187 $Y=1.18
r28 16 23 12.6543 $w=2.53e-07 $l=2.8e-07 $layer=LI1_cond $X=1.187 $Y=0.925
+ $X2=1.187 $Y2=0.645
r29 15 23 4.06745 $w=2.53e-07 $l=9e-08 $layer=LI1_cond $X=1.187 $Y=0.555
+ $X2=1.187 $Y2=0.645
r30 12 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=2.015
+ $X2=1.225 $Y2=1.85
r31 10 13 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.145 $Y=1.18
+ $X2=1.145 $Y2=1.85
r32 9 16 5.78481 $w=2.53e-07 $l=1.28e-07 $layer=LI1_cond $X=1.187 $Y=1.053
+ $X2=1.187 $Y2=0.925
r33 9 10 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=1.187 $Y=1.053
+ $X2=1.187 $Y2=1.18
r34 2 12 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.84 $X2=1.225 $Y2=2.015
r35 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.09
+ $Y=0.5 $X2=1.23 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__OR4BB_2%VGND 1 2 3 4 15 19 22 25 28 29 33 35 37 42
+ 51 57 58 61 64 67
r81 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r82 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r83 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r84 58 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r85 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r86 55 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.255 $Y=0 $X2=4.09
+ $Y2=0
r87 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.255 $Y=0 $X2=4.56
+ $Y2=0
r88 54 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r89 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r90 51 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=4.09
+ $Y2=0
r91 51 53 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=3.6
+ $Y2=0
r92 50 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r93 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r94 47 64 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=1.805
+ $Y2=0
r95 47 49 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=2.64
+ $Y2=0
r96 46 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r97 46 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r98 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r99 43 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.755
+ $Y2=0
r100 43 45 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.2
+ $Y2=0
r101 42 64 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=1.805
+ $Y2=0
r102 42 45 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=1.2
+ $Y2=0
r103 40 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r104 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r105 37 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.755
+ $Y2=0
r106 37 39 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.24
+ $Y2=0
r107 35 50 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r108 35 65 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r109 30 33 7.07181 $w=2.18e-07 $l=1.35e-07 $layer=LI1_cond $X=2.895 $Y=0.85
+ $X2=3.03 $Y2=0.85
r110 28 49 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.64
+ $Y2=0
r111 28 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.895
+ $Y2=0
r112 27 53 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.98 $Y=0 $X2=3.6
+ $Y2=0
r113 27 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=0 $X2=2.895
+ $Y2=0
r114 23 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=0.085
+ $X2=4.09 $Y2=0
r115 23 25 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=4.09 $Y=0.085
+ $X2=4.09 $Y2=0.61
r116 22 30 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.895 $Y=0.74
+ $X2=2.895 $Y2=0.85
r117 21 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=0.085
+ $X2=2.895 $Y2=0
r118 21 22 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.895 $Y=0.085
+ $X2=2.895 $Y2=0.74
r119 17 64 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=0.085
+ $X2=1.805 $Y2=0
r120 17 19 18.3312 $w=4.58e-07 $l=7.05e-07 $layer=LI1_cond $X=1.805 $Y=0.085
+ $X2=1.805 $Y2=0.79
r121 13 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0
r122 13 15 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0.66
r123 4 25 182 $w=1.7e-07 $l=2.52587e-07 $layer=licon1_NDIFF $count=1 $X=3.87
+ $Y=0.68 $X2=4.09 $Y2=0.61
r124 3 33 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=2.89
+ $Y=0.68 $X2=3.03 $Y2=0.85
r125 2 19 182 $w=1.7e-07 $l=4.20714e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.5 $X2=1.82 $Y2=0.79
r126 1 15 182 $w=1.7e-07 $l=2.34521e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.69 $X2=0.795 $Y2=0.66
.ends

