* File: sky130_fd_sc_ls__decaphe_2.pex.spice
* Created: Wed Sep  2 10:59:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DECAPHE_2%VGND 3 5 7 10 14 18 19
r11 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r12 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r13 16 22 5.34931 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.235
+ $Y2=0
r14 16 18 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.72
+ $Y2=0
r15 10 19 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=0 $X2=0.72
+ $Y2=0
r16 10 23 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=0 $X2=0.24
+ $Y2=0
r17 8 14 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.48 $Y2=1.465
r18 7 8 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r19 5 22 2.89091 $w=3.85e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.277 $Y=0.085
+ $X2=0.235 $Y2=0
r20 5 7 41.3083 $w=3.83e-07 $l=1.38e-06 $layer=LI1_cond $X=0.277 $Y=0.085
+ $X2=0.277 $Y2=1.465
r21 1 14 18.2676 $w=1.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.63
+ $X2=0.48 $Y2=1.465
r22 1 3 353.889 $w=1.7e-07 $l=8.37e-07 $layer=POLY_cond $X=0.48 $Y=1.63 $X2=0.48
+ $Y2=2.467
.ends

.subckt PM_SKY130_FD_SC_LS__DECAPHE_2%VPWR 1 9 15 18 24
r7 19 24 0.0166838 $w=9.6e-07 $l=1.22e-07 $layer=MET1_cond $X=0.48 $Y=3.33
+ $X2=0.48 $Y2=3.208
r8 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r9 15 24 0.000136752 $w=9.6e-07 $l=1e-09 $layer=MET1_cond $X=0.48 $Y=3.207
+ $X2=0.48 $Y2=3.208
r10 9 13 14.6103 $w=7.88e-07 $l=9.65e-07 $layer=LI1_cond $X=0.48 $Y=1.985
+ $X2=0.48 $Y2=2.95
r11 7 18 1.49888 $w=9.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.48 $Y=3.245
+ $X2=0.48 $Y2=3.33
r12 7 13 4.46637 $w=7.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.48 $Y=3.245
+ $X2=0.48 $Y2=2.95
r13 1 13 400 $w=1.7e-07 $l=1.17556e-06 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.84 $X2=0.7 $Y2=2.95
r14 1 13 400 $w=1.7e-07 $l=1.17083e-06 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.84 $X2=0.26 $Y2=2.95
r15 1 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.84 $X2=0.7 $Y2=1.985
r16 1 9 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.84 $X2=0.26 $Y2=1.985
.ends

