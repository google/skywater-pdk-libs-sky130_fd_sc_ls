* File: sky130_fd_sc_ls__clkbuf_1.spice
* Created: Wed Sep  2 10:57:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__clkbuf_1.pex.spice"
.subckt sky130_fd_sc_ls__clkbuf_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_27_74#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1638 AS=0.1197 PD=1.2 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_27_74#_M1002_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.119 AS=0.1638 PD=1.41 PS=1.2 NRD=0 NRS=19.992 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_27_74#_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.3304 PD=1.52 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1001 N_X_M1001_d N_A_27_74#_M1001_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.224 PD=2.83 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.8 SB=75000.2 A=0.168 P=2.54 MULT=1
DX4_noxref VNB VPB NWDIODE A=4.278 P=8.32
*
.include "sky130_fd_sc_ls__clkbuf_1.pxi.spice"
*
.ends
*
*
