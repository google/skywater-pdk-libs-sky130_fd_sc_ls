* File: sky130_fd_sc_ls__dlxbn_2.spice
* Created: Fri Aug 28 13:19:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dlxbn_2.pex.spice"
.subckt sky130_fd_sc_ls__dlxbn_2  VNB VPB D GATE_N VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_D_M1021_g N_A_27_136#_M1021_s VNB NSHORT L=0.15 W=0.55
+ AD=0.171076 AS=0.15675 PD=1.27054 PS=1.67 NRD=55.86 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1001 N_A_232_98#_M1001_d N_GATE_N_M1001_g N_VGND_M1021_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.230174 PD=2.05 PS=1.70946 NRD=0 NRS=41.52 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A_232_98#_M1005_g N_A_343_74#_M1005_s VNB NSHORT L=0.15
+ W=0.74 AD=0.206959 AS=0.2817 PD=1.49609 PS=2.29 NRD=36.432 NRS=2.016 M=1
+ R=4.93333 SA=75000.3 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1012 A_569_79# N_A_27_136#_M1012_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.178991 PD=0.88 PS=1.29391 NRD=12.18 NRS=18.744 M=1 R=4.26667
+ SA=75000.9 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1013 N_A_647_79#_M1013_d N_A_232_98#_M1013_g A_569_79# VNB NSHORT L=0.15
+ W=0.64 AD=0.238611 AS=0.0768 PD=1.75094 PS=0.88 NRD=27.18 NRS=12.18 M=1
+ R=4.26667 SA=75001.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1025 A_839_123# N_A_343_74#_M1025_g N_A_647_79#_M1013_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0651 AS=0.156589 PD=0.73 PS=1.14906 NRD=28.56 NRS=0 M=1 R=2.8
+ SA=75002.3 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_A_887_270#_M1023_g A_839_123# VNB NSHORT L=0.15 W=0.42
+ AD=0.0905534 AS=0.0651 PD=0.829138 PS=0.73 NRD=7.14 NRS=28.56 M=1 R=2.8
+ SA=75002.7 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1016 N_A_887_270#_M1016_d N_A_647_79#_M1016_g N_VGND_M1023_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.159547 PD=2.05 PS=1.46086 NRD=0 NRS=16.212 M=1 R=4.93333
+ SA=75001.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_Q_M1002_d N_A_887_270#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1009 N_Q_M1002_d N_A_887_270#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.166607 PD=1.02 PS=1.25478 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1017 N_A_1442_94#_M1017_d N_A_887_270#_M1017_g N_VGND_M1009_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.144093 PD=1.85 PS=1.08522 NRD=0 NRS=15.468 M=1
+ R=4.26667 SA=75001.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_Q_N_M1007_d N_A_1442_94#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.3 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1015 N_Q_N_M1007_d N_A_1442_94#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_D_M1000_g N_A_27_136#_M1000_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.147 AS=0.3192 PD=1.19 PS=2.44 NRD=2.3443 NRS=22.261 M=1 R=5.6 SA=75000.3
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1006 N_A_232_98#_M1006_d N_GATE_N_M1006_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.147 PD=2.27 PS=1.19 NRD=2.3443 NRS=14.0658 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_VPWR_M1008_d N_A_232_98#_M1008_g N_A_343_74#_M1008_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.169187 AS=0.2478 PD=1.26457 PS=2.27 NRD=23.443 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75002.2 A=0.126 P=1.98 MULT=1
MM1022 A_565_392# N_A_27_136#_M1022_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.201413 PD=1.27 PS=1.50543 NRD=15.7403 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1014 N_A_647_79#_M1014_d N_A_343_74#_M1014_g A_565_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.307887 AS=0.135 PD=2.35915 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75001.1 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1004 A_814_392# N_A_232_98#_M1004_g N_A_647_79#_M1014_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0798 AS=0.129313 PD=0.8 PS=0.990845 NRD=63.3158 NRS=4.6886 M=1
+ R=2.8 SA=75002 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1018 N_VPWR_M1018_d N_A_887_270#_M1018_g A_814_392# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.134891 AS=0.0798 PD=0.891818 PS=0.8 NRD=63.3158 NRS=63.3158 M=1 R=2.8
+ SA=75002.5 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1019 N_A_887_270#_M1019_d N_A_647_79#_M1019_g N_VPWR_M1018_d VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.3304 AS=0.359709 PD=2.83 PS=2.37818 NRD=1.7533 NRS=17.5724
+ M=1 R=7.46667 SA=75001.4 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1003_d N_A_887_270#_M1003_g N_Q_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1024 N_VPWR_M1024_d N_A_887_270#_M1024_g N_Q_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.204347 AS=0.168 PD=1.55849 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1010 N_A_1442_94#_M1010_d N_A_887_270#_M1010_g N_VPWR_M1024_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.182453 PD=2.59 PS=1.39151 NRD=1.9503 NRS=12.7853 M=1
+ R=6.66667 SA=75001.2 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1011 N_Q_N_M1011_d N_A_1442_94#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1020 N_Q_N_M1011_d N_A_1442_94#_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX26_noxref VNB VPB NWDIODE A=17.67 P=22.72
c_89 VNB 0 1.28661e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__dlxbn_2.pxi.spice"
*
.ends
*
*
