* File: sky130_fd_sc_ls__and2_2.pxi.spice
* Created: Fri Aug 28 13:02:45 2020
* 
x_PM_SKY130_FD_SC_LS__AND2_2%A N_A_c_52_n N_A_c_57_n N_A_M1005_g N_A_M1003_g A
+ N_A_c_54_n N_A_c_55_n PM_SKY130_FD_SC_LS__AND2_2%A
x_PM_SKY130_FD_SC_LS__AND2_2%B N_B_M1001_g N_B_c_82_n N_B_c_86_n N_B_M1006_g B
+ N_B_c_83_n N_B_c_84_n PM_SKY130_FD_SC_LS__AND2_2%B
x_PM_SKY130_FD_SC_LS__AND2_2%A_31_74# N_A_31_74#_M1003_s N_A_31_74#_M1005_d
+ N_A_31_74#_c_126_n N_A_31_74#_M1002_g N_A_31_74#_c_134_n N_A_31_74#_M1000_g
+ N_A_31_74#_c_127_n N_A_31_74#_M1007_g N_A_31_74#_c_135_n N_A_31_74#_M1004_g
+ N_A_31_74#_c_128_n N_A_31_74#_c_129_n N_A_31_74#_c_130_n N_A_31_74#_c_136_n
+ N_A_31_74#_c_137_n N_A_31_74#_c_138_n N_A_31_74#_c_131_n N_A_31_74#_c_132_n
+ N_A_31_74#_c_133_n PM_SKY130_FD_SC_LS__AND2_2%A_31_74#
x_PM_SKY130_FD_SC_LS__AND2_2%VPWR N_VPWR_M1005_s N_VPWR_M1006_d N_VPWR_M1004_d
+ N_VPWR_c_220_n N_VPWR_c_221_n N_VPWR_c_222_n N_VPWR_c_223_n N_VPWR_c_224_n
+ VPWR N_VPWR_c_225_n N_VPWR_c_226_n N_VPWR_c_227_n N_VPWR_c_219_n
+ PM_SKY130_FD_SC_LS__AND2_2%VPWR
x_PM_SKY130_FD_SC_LS__AND2_2%X N_X_M1002_d N_X_M1000_s N_X_c_257_n N_X_c_258_n
+ N_X_c_260_n X X X PM_SKY130_FD_SC_LS__AND2_2%X
x_PM_SKY130_FD_SC_LS__AND2_2%VGND N_VGND_M1001_d N_VGND_M1007_s N_VGND_c_291_n
+ N_VGND_c_292_n N_VGND_c_293_n VGND N_VGND_c_294_n N_VGND_c_295_n
+ N_VGND_c_296_n N_VGND_c_297_n PM_SKY130_FD_SC_LS__AND2_2%VGND
cc_1 VNB N_A_c_52_n 0.00192204f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.795
cc_2 VNB N_A_M1003_g 0.0297549f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_3 VNB N_A_c_54_n 0.0050357f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_A_c_55_n 0.0582211f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.465
cc_5 VNB N_B_M1001_g 0.0215375f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.885
cc_6 VNB N_B_c_82_n 0.00136699f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.3
cc_7 VNB N_B_c_83_n 0.0291159f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_8 VNB N_B_c_84_n 0.00419749f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_9 VNB N_A_31_74#_c_126_n 0.0174733f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_10 VNB N_A_31_74#_c_127_n 0.0188592f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_11 VNB N_A_31_74#_c_128_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_12 VNB N_A_31_74#_c_129_n 0.00780948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_31_74#_c_130_n 0.00898165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_31_74#_c_131_n 0.00473431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_31_74#_c_132_n 6.4908e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_31_74#_c_133_n 0.056599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_219_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_X_c_257_n 0.00239236f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_19 VNB N_X_c_258_n 0.0188945f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_20 VNB N_VGND_c_291_n 0.006479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_292_n 0.0118321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_293_n 0.0255459f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_23 VNB N_VGND_c_294_n 0.029813f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.465
cc_24 VNB N_VGND_c_295_n 0.0193156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_296_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_297_n 0.166974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VPB N_A_c_52_n 0.00915684f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.795
cc_28 VPB N_A_c_57_n 0.028153f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.885
cc_29 VPB N_A_c_54_n 0.00745299f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_30 VPB N_B_c_82_n 0.00650397f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.3
cc_31 VPB N_B_c_86_n 0.0223997f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=0.74
cc_32 VPB N_B_c_84_n 0.00533089f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_33 VPB N_A_31_74#_c_134_n 0.015159f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_34 VPB N_A_31_74#_c_135_n 0.0165392f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.465
cc_35 VPB N_A_31_74#_c_136_n 0.0020678f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_A_31_74#_c_137_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_A_31_74#_c_138_n 7.05414e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_A_31_74#_c_132_n 0.00133441f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_31_74#_c_133_n 0.0140421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_220_n 0.0117486f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_41 VPB N_VPWR_c_221_n 0.0501311f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_42 VPB N_VPWR_c_222_n 0.0052096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_223_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_224_n 0.0461938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_225_n 0.0175706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_226_n 0.0186844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_227_n 0.00614589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_219_n 0.0571235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_X_c_258_n 0.00210119f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=0.74
cc_50 VPB N_X_c_260_n 0.00958413f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_51 VPB X 0.00217096f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.465
cc_52 N_A_M1003_g N_B_M1001_g 0.0550561f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_53 N_A_c_52_n N_B_c_82_n 0.00581924f $X=0.5 $Y=1.795 $X2=0 $Y2=0
cc_54 N_A_c_57_n N_B_c_86_n 0.0139779f $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_55 N_A_c_54_n N_B_c_83_n 2.28826e-19 $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_56 N_A_c_55_n N_B_c_83_n 0.0209293f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_57 N_A_c_54_n N_B_c_84_n 0.0391299f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_58 N_A_c_55_n N_B_c_84_n 0.00404395f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_59 N_A_M1003_g N_A_31_74#_c_128_n 0.012125f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_60 N_A_M1003_g N_A_31_74#_c_129_n 0.0146407f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_61 N_A_M1003_g N_A_31_74#_c_130_n 0.00206782f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_62 N_A_c_54_n N_A_31_74#_c_130_n 0.0260039f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_63 N_A_c_55_n N_A_31_74#_c_130_n 0.00265493f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_64 N_A_c_57_n N_A_31_74#_c_136_n 7.89448e-19 $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_65 N_A_c_57_n N_A_31_74#_c_137_n 0.00304898f $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_66 N_A_c_57_n N_VPWR_c_221_n 0.016367f $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_67 N_A_c_54_n N_VPWR_c_221_n 0.0293457f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_68 N_A_c_55_n N_VPWR_c_221_n 0.00165041f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_69 N_A_c_57_n N_VPWR_c_225_n 0.00413917f $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_70 N_A_c_57_n N_VPWR_c_219_n 0.0081781f $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_71 N_A_M1003_g N_VGND_c_291_n 0.00180653f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_72 N_A_M1003_g N_VGND_c_294_n 0.00434272f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_73 N_A_M1003_g N_VGND_c_297_n 0.00824704f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_74 N_B_M1001_g N_A_31_74#_c_126_n 0.0259185f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_75 N_B_c_82_n N_A_31_74#_c_134_n 0.00382859f $X=0.95 $Y=1.795 $X2=0 $Y2=0
cc_76 N_B_c_86_n N_A_31_74#_c_134_n 0.0243716f $X=0.95 $Y=1.885 $X2=0 $Y2=0
cc_77 N_B_M1001_g N_A_31_74#_c_128_n 0.00208517f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_78 N_B_M1001_g N_A_31_74#_c_129_n 0.0144246f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_79 N_B_c_83_n N_A_31_74#_c_129_n 0.00493688f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_80 N_B_c_84_n N_A_31_74#_c_129_n 0.0374224f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_81 N_B_c_86_n N_A_31_74#_c_136_n 9.93639e-19 $X=0.95 $Y=1.885 $X2=0 $Y2=0
cc_82 N_B_c_83_n N_A_31_74#_c_136_n 3.30055e-19 $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_83 N_B_c_84_n N_A_31_74#_c_136_n 0.0225259f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_84 N_B_c_86_n N_A_31_74#_c_137_n 0.00996212f $X=0.95 $Y=1.885 $X2=0 $Y2=0
cc_85 N_B_c_86_n N_A_31_74#_c_138_n 0.0126729f $X=0.95 $Y=1.885 $X2=0 $Y2=0
cc_86 N_B_c_83_n N_A_31_74#_c_138_n 0.00166044f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_87 N_B_c_84_n N_A_31_74#_c_138_n 0.0147428f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_88 N_B_M1001_g N_A_31_74#_c_131_n 0.00350413f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_89 N_B_c_83_n N_A_31_74#_c_131_n 0.00159524f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_90 N_B_c_84_n N_A_31_74#_c_131_n 0.0208197f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_91 N_B_c_82_n N_A_31_74#_c_132_n 0.00258519f $X=0.95 $Y=1.795 $X2=0 $Y2=0
cc_92 N_B_c_86_n N_A_31_74#_c_132_n 0.00127545f $X=0.95 $Y=1.885 $X2=0 $Y2=0
cc_93 N_B_c_83_n N_A_31_74#_c_132_n 4.8742e-19 $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_94 N_B_c_84_n N_A_31_74#_c_132_n 0.0184082f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_95 N_B_c_82_n N_A_31_74#_c_133_n 0.00499917f $X=0.95 $Y=1.795 $X2=0 $Y2=0
cc_96 N_B_c_83_n N_A_31_74#_c_133_n 0.0198726f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_97 N_B_c_84_n N_A_31_74#_c_133_n 7.22997e-19 $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_98 N_B_c_86_n N_VPWR_c_221_n 6.58931e-19 $X=0.95 $Y=1.885 $X2=0 $Y2=0
cc_99 N_B_c_86_n N_VPWR_c_222_n 0.00546864f $X=0.95 $Y=1.885 $X2=0 $Y2=0
cc_100 N_B_c_86_n N_VPWR_c_225_n 0.00445602f $X=0.95 $Y=1.885 $X2=0 $Y2=0
cc_101 N_B_c_86_n N_VPWR_c_219_n 0.00857556f $X=0.95 $Y=1.885 $X2=0 $Y2=0
cc_102 N_B_M1001_g N_VGND_c_291_n 0.0120683f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_103 N_B_M1001_g N_VGND_c_294_n 0.00383152f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_104 N_B_M1001_g N_VGND_c_297_n 0.0075725f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_31_74#_c_138_n N_VPWR_M1006_d 0.00749749f $X=1.255 $Y=2.035 $X2=0
+ $Y2=0
cc_106 N_A_31_74#_c_132_n N_VPWR_M1006_d 0.00131481f $X=1.34 $Y=1.95 $X2=0 $Y2=0
cc_107 N_A_31_74#_c_136_n N_VPWR_c_221_n 0.0123997f $X=0.765 $Y=2.12 $X2=0 $Y2=0
cc_108 N_A_31_74#_c_137_n N_VPWR_c_221_n 0.0576594f $X=0.725 $Y=2.815 $X2=0
+ $Y2=0
cc_109 N_A_31_74#_c_134_n N_VPWR_c_222_n 0.0107533f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_110 N_A_31_74#_c_135_n N_VPWR_c_222_n 5.65429e-19 $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_111 N_A_31_74#_c_137_n N_VPWR_c_222_n 0.0256025f $X=0.725 $Y=2.815 $X2=0
+ $Y2=0
cc_112 N_A_31_74#_c_138_n N_VPWR_c_222_n 0.020844f $X=1.255 $Y=2.035 $X2=0 $Y2=0
cc_113 N_A_31_74#_c_135_n N_VPWR_c_224_n 0.0104242f $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_114 N_A_31_74#_c_137_n N_VPWR_c_225_n 0.0110241f $X=0.725 $Y=2.815 $X2=0
+ $Y2=0
cc_115 N_A_31_74#_c_134_n N_VPWR_c_226_n 0.00429299f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_116 N_A_31_74#_c_135_n N_VPWR_c_226_n 0.00445602f $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_117 N_A_31_74#_c_134_n N_VPWR_c_219_n 0.00847721f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_118 N_A_31_74#_c_135_n N_VPWR_c_219_n 0.0086105f $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_119 N_A_31_74#_c_137_n N_VPWR_c_219_n 0.00909194f $X=0.725 $Y=2.815 $X2=0
+ $Y2=0
cc_120 N_A_31_74#_c_126_n N_X_c_257_n 0.0105697f $X=1.415 $Y=1.22 $X2=0 $Y2=0
cc_121 N_A_31_74#_c_127_n N_X_c_257_n 0.0249871f $X=1.845 $Y=1.22 $X2=0 $Y2=0
cc_122 N_A_31_74#_c_131_n N_X_c_257_n 0.0126837f $X=1.34 $Y=1.55 $X2=0 $Y2=0
cc_123 N_A_31_74#_c_133_n N_X_c_257_n 0.0010614f $X=1.845 $Y=1.492 $X2=0 $Y2=0
cc_124 N_A_31_74#_c_126_n N_X_c_258_n 6.22718e-19 $X=1.415 $Y=1.22 $X2=0 $Y2=0
cc_125 N_A_31_74#_c_127_n N_X_c_258_n 0.00695403f $X=1.845 $Y=1.22 $X2=0 $Y2=0
cc_126 N_A_31_74#_c_131_n N_X_c_258_n 0.0311249f $X=1.34 $Y=1.55 $X2=0 $Y2=0
cc_127 N_A_31_74#_c_132_n N_X_c_258_n 0.00559f $X=1.34 $Y=1.95 $X2=0 $Y2=0
cc_128 N_A_31_74#_c_133_n N_X_c_258_n 0.0231474f $X=1.845 $Y=1.492 $X2=0 $Y2=0
cc_129 N_A_31_74#_c_134_n N_X_c_260_n 7.38062e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A_31_74#_c_135_n N_X_c_260_n 0.0102846f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A_31_74#_c_131_n N_X_c_260_n 0.00566518f $X=1.34 $Y=1.55 $X2=0 $Y2=0
cc_132 N_A_31_74#_c_132_n N_X_c_260_n 0.0128811f $X=1.34 $Y=1.95 $X2=0 $Y2=0
cc_133 N_A_31_74#_c_133_n N_X_c_260_n 0.00672165f $X=1.845 $Y=1.492 $X2=0 $Y2=0
cc_134 N_A_31_74#_c_134_n X 0.00703236f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A_31_74#_c_135_n X 0.0177445f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A_31_74#_c_138_n X 0.0137304f $X=1.255 $Y=2.035 $X2=0 $Y2=0
cc_137 N_A_31_74#_c_132_n X 0.00430791f $X=1.34 $Y=1.95 $X2=0 $Y2=0
cc_138 N_A_31_74#_c_129_n A_118_74# 0.0048076f $X=1.255 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_139 N_A_31_74#_c_129_n N_VGND_M1001_d 0.00230675f $X=1.255 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_140 N_A_31_74#_c_131_n N_VGND_M1001_d 3.09855e-19 $X=1.34 $Y=1.55 $X2=-0.19
+ $Y2=-0.245
cc_141 N_A_31_74#_c_126_n N_VGND_c_291_n 0.00543307f $X=1.415 $Y=1.22 $X2=0
+ $Y2=0
cc_142 N_A_31_74#_c_128_n N_VGND_c_291_n 0.0139395f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_143 N_A_31_74#_c_129_n N_VGND_c_291_n 0.0195279f $X=1.255 $Y=1.045 $X2=0
+ $Y2=0
cc_144 N_A_31_74#_c_131_n N_VGND_c_291_n 0.00252453f $X=1.34 $Y=1.55 $X2=0 $Y2=0
cc_145 N_A_31_74#_c_127_n N_VGND_c_293_n 0.00500034f $X=1.845 $Y=1.22 $X2=0
+ $Y2=0
cc_146 N_A_31_74#_c_128_n N_VGND_c_294_n 0.0145639f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_147 N_A_31_74#_c_126_n N_VGND_c_295_n 0.00433139f $X=1.415 $Y=1.22 $X2=0
+ $Y2=0
cc_148 N_A_31_74#_c_127_n N_VGND_c_295_n 0.00433139f $X=1.845 $Y=1.22 $X2=0
+ $Y2=0
cc_149 N_A_31_74#_c_126_n N_VGND_c_297_n 0.00817409f $X=1.415 $Y=1.22 $X2=0
+ $Y2=0
cc_150 N_A_31_74#_c_127_n N_VGND_c_297_n 0.00451721f $X=1.845 $Y=1.22 $X2=0
+ $Y2=0
cc_151 N_A_31_74#_c_128_n N_VGND_c_297_n 0.0119984f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_152 N_VPWR_c_222_n X 0.0454264f $X=1.225 $Y=2.455 $X2=0 $Y2=0
cc_153 N_VPWR_c_224_n X 0.0604541f $X=2.13 $Y=2.225 $X2=0 $Y2=0
cc_154 N_VPWR_c_226_n X 0.0110241f $X=2.045 $Y=3.33 $X2=0 $Y2=0
cc_155 N_VPWR_c_219_n X 0.00909194f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_156 N_X_c_257_n N_VGND_M1007_s 0.00752423f $X=1.925 $Y=1.02 $X2=0 $Y2=0
cc_157 N_X_c_258_n N_VGND_M1007_s 0.00339584f $X=1.925 $Y=1.72 $X2=0 $Y2=0
cc_158 N_X_c_257_n N_VGND_c_291_n 0.0166176f $X=1.925 $Y=1.02 $X2=0 $Y2=0
cc_159 N_X_c_257_n N_VGND_c_293_n 0.0155529f $X=1.925 $Y=1.02 $X2=0 $Y2=0
cc_160 N_X_c_257_n N_VGND_c_295_n 0.0143518f $X=1.925 $Y=1.02 $X2=0 $Y2=0
cc_161 N_X_c_257_n N_VGND_c_297_n 0.0179048f $X=1.925 $Y=1.02 $X2=0 $Y2=0
