* File: sky130_fd_sc_ls__a41oi_2.spice
* Created: Fri Aug 28 13:02:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a41oi_2.pex.spice"
.subckt sky130_fd_sc_ls__a41oi_2  VNB VPB B1 A1 A2 A3 A4 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1007 N_Y_M1007_d N_B1_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1004_d N_A1_M1004_g N_A_239_74#_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1016 N_Y_M1004_d N_A1_M1016_g N_A_239_74#_M1016_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1003 N_A_239_74#_M1016_s N_A2_M1003_g N_A_512_74#_M1003_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1011 N_A_239_74#_M1011_d N_A2_M1011_g N_A_512_74#_M1003_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_709_74#_M1000_d N_A3_M1000_g N_A_512_74#_M1000_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1012 N_A_709_74#_M1012_d N_A3_M1012_g N_A_512_74#_M1000_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1008 N_A_709_74#_M1012_d N_A4_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1221 PD=1.02 PS=1.07 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1010 N_A_709_74#_M1010_d N_A4_M1010_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2257 AS=0.1221 PD=2.09 PS=1.07 NRD=3.24 NRS=8.1 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_27_368#_M1006_d N_B1_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.2 SB=75005 A=0.168 P=2.54 MULT=1
MM1009 N_A_27_368#_M1009_d N_B1_M1009_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75004.5 A=0.168 P=2.54 MULT=1
MM1005 N_A_27_368#_M1009_d N_A1_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.3304 PD=1.47 PS=1.71 NRD=1.7533 NRS=27.2451 M=1 R=7.46667
+ SA=75001.2 SB=75004 A=0.168 P=2.54 MULT=1
MM1015 N_A_27_368#_M1015_d N_A1_M1015_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=1.71 NRD=1.7533 NRS=27.2451 M=1 R=7.46667
+ SA=75002 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1013_d N_A2_M1013_g N_A_27_368#_M1015_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.4 SB=75002.8 A=0.168 P=2.54 MULT=1
MM1018 N_VPWR_M1013_d N_A2_M1018_g N_A_27_368#_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1001 N_VPWR_M1001_d N_A3_M1001_g N_A_27_368#_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.4 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1001_d N_A3_M1002_g N_A_27_368#_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.2156 PD=1.52 PS=1.505 NRD=10.5395 NRS=4.3931 M=1 R=7.46667
+ SA=75004 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1014_d N_A4_M1014_g N_A_27_368#_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.2156 PD=1.42 PS=1.505 NRD=1.7533 NRS=14.0658 M=1 R=7.46667
+ SA=75004.5 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1017 N_VPWR_M1014_d N_A4_M1017_g N_A_27_368#_M1017_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3584 PD=1.42 PS=2.88 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75004.9 SB=75000.2 A=0.168 P=2.54 MULT=1
DX19_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ls__a41oi_2.pxi.spice"
*
.ends
*
*
