* File: sky130_fd_sc_ls__a31oi_4.spice
* Created: Wed Sep  2 10:52:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a31oi_4.pex.spice"
.subckt sky130_fd_sc_ls__a31oi_4  VNB VPB A3 A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1009 N_A_30_74#_M1009_d N_A3_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1011 N_A_30_74#_M1011_d N_A3_M1011_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1026 N_A_30_74#_M1011_d N_A3_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1027 N_A_30_74#_M1027_d N_A3_M1027_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.6
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1004 N_A_475_74#_M1004_d N_A2_M1004_g N_A_30_74#_M1027_d VNB NSHORT L=0.15
+ W=0.74 AD=0.1073 AS=0.1036 PD=1.03 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75002 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1008 N_A_475_74#_M1004_d N_A2_M1008_g N_A_30_74#_M1008_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1073 AS=0.1036 PD=1.03 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1012 N_A_475_74#_M1012_d N_A2_M1012_g N_A_30_74#_M1008_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1020 N_A_475_74#_M1012_d N_A2_M1020_g N_A_30_74#_M1020_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1554 AS=0.202325 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75003.4 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_475_74#_M1005_d N_A1_M1005_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.19805 PD=1.31 PS=2.07 NRD=23.508 NRS=0.804 M=1 R=4.93333
+ SA=75000.2 SB=75003.6 A=0.111 P=1.78 MULT=1
MM1017 N_A_475_74#_M1005_d N_A1_M1017_g N_Y_M1017_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=1.31 PS=1.09 NRD=23.508 NRS=0 M=1 R=4.93333 SA=75000.9
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1018 N_A_475_74#_M1018_d N_A1_M1018_g N_Y_M1017_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.4
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1029 N_A_475_74#_M1018_d N_A1_M1029_g N_Y_M1029_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.8
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1029_s N_B1_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.40885 PD=1.09 PS=1.845 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1024 N_Y_M1024_d N_B1_M1024_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.40885 PD=2.05 PS=1.845 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_A_27_368#_M1001_d N_A3_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75007.8 A=0.168 P=2.54 MULT=1
MM1015 N_A_27_368#_M1015_d N_A3_M1015_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75007.4 A=0.168 P=2.54 MULT=1
MM1016 N_A_27_368#_M1015_d N_A3_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75006.9 A=0.168 P=2.54 MULT=1
MM1022 N_A_27_368#_M1022_d N_A3_M1022_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75006.5 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A2_M1006_g N_A_27_368#_M1022_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75006 A=0.168 P=2.54 MULT=1
MM1010 N_VPWR_M1006_d N_A2_M1010_g N_A_27_368#_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75005.5 A=0.168 P=2.54 MULT=1
MM1019 N_VPWR_M1019_d N_A2_M1019_g N_A_27_368#_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003 SB=75005.1 A=0.168 P=2.54 MULT=1
MM1025 N_VPWR_M1019_d N_A2_M1025_g N_A_27_368#_M1025_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.5 SB=75004.6 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_27_368#_M1025_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75004 SB=75004.1 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1002_d N_A1_M1003_g N_A_27_368#_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.4648 PD=1.47 PS=1.95 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75004.5 SB=75003.6 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_27_368#_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.4648 PD=1.52 PS=1.95 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75005.4 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1028 N_VPWR_M1007_d N_A1_M1028_g N_A_27_368#_M1028_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.224 AS=0.1848 PD=1.52 PS=1.45 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75006 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1000 N_A_27_368#_M1028_s N_B1_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1848 AS=0.1792 PD=1.45 PS=1.44 NRD=7.0329 NRS=5.2599 M=1 R=7.46667
+ SA=75006.5 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1014 N_A_27_368#_M1014_d N_B1_M1014_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.1792 PD=1.42 PS=1.44 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.9 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1021 N_A_27_368#_M1014_d N_B1_M1021_g N_Y_M1021_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.4 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1023 N_A_27_368#_M1023_d N_B1_M1023_g N_Y_M1021_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.8 SB=75000.2 A=0.168 P=2.54 MULT=1
DX30_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_ls__a31oi_4.pxi.spice"
*
.ends
*
*
