* File: sky130_fd_sc_ls__and4b_4.spice
* Created: Wed Sep  2 10:55:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__and4b_4.pex.spice"
.subckt sky130_fd_sc_ls__and4b_4  VNB VPB A_N D C B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* C	C
* D	D
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_A_N_M1014_g N_A_27_368#_M1014_s VNB NSHORT L=0.15 W=0.64
+ AD=0.131803 AS=0.1824 PD=1.06203 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.3 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1014_d N_A_199_294#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.152397 AS=0.1036 PD=1.22797 PS=1.02 NRD=20.268 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_199_294#_M1013_g N_X_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1813 AS=0.1036 PD=1.23 PS=1.02 NRD=16.212 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1013_d N_A_199_294#_M1021_g N_X_M1021_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1813 AS=0.1036 PD=1.23 PS=1.02 NRD=17.832 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1025 N_VGND_M1025_d N_A_199_294#_M1025_g N_X_M1021_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1000 N_A_664_125#_M1000_d N_C_M1000_g N_A_751_125#_M1000_s VNB NSHORT L=0.15
+ W=0.64 AD=0.178725 AS=0.104 PD=1.85 PS=0.965 NRD=0 NRS=3.744 M=1 R=4.26667
+ SA=75000.2 SB=75003.6 A=0.096 P=1.58 MULT=1
MM1012 N_VGND_M1012_d N_D_M1012_g N_A_751_125#_M1000_s VNB NSHORT L=0.15 W=0.64
+ AD=0.174875 AS=0.104 PD=1.315 PS=0.965 NRD=40.92 NRS=4.68 M=1 R=4.26667
+ SA=75000.7 SB=75003.2 A=0.096 P=1.58 MULT=1
MM1020 N_VGND_M1012_d N_D_M1020_g N_A_751_125#_M1020_s VNB NSHORT L=0.15 W=0.64
+ AD=0.174875 AS=0.0896 PD=1.315 PS=0.92 NRD=40.92 NRS=0 M=1 R=4.26667
+ SA=75001.3 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1017 N_A_664_125#_M1017_d N_C_M1017_g N_A_751_125#_M1020_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.7 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1005 N_A_664_125#_M1017_d N_B_M1005_g N_A_1136_125#_M1005_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.1 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1015 N_A_1136_125#_M1005_s N_A_27_368#_M1015_g N_A_199_294#_M1015_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.6 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1023 N_A_1136_125#_M1023_d N_A_27_368#_M1023_g N_A_199_294#_M1015_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.16 AS=0.0896 PD=1.14 PS=0.92 NRD=20.616 NRS=0 M=1 R=4.26667
+ SA=75003 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1019 N_A_664_125#_M1019_d N_B_M1019_g N_A_1136_125#_M1023_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1792 AS=0.16 PD=1.84 PS=1.14 NRD=0 NRS=20.616 M=1 R=4.26667
+ SA=75003.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_A_N_M1016_g N_A_27_368#_M1016_s VPB PHIGHVT L=0.15 W=1
+ AD=0.222075 AS=0.295 PD=1.46226 PS=2.59 NRD=23.6203 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75006.3 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1016_d N_A_199_294#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.248725 AS=0.168 PD=1.63774 PS=1.42 NRD=6.1464 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75005.8 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1004_d N_A_199_294#_M1004_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1848 AS=0.168 PD=1.45 PS=1.42 NRD=4.3931 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75005.4 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1004_d N_A_199_294#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1848 AS=0.2296 PD=1.45 PS=1.53 NRD=4.3931 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75004.9 A=0.168 P=2.54 MULT=1
MM1022 N_VPWR_M1022_d N_A_199_294#_M1022_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.228121 AS=0.2296 PD=1.60604 PS=1.53 NRD=2.6201 NRS=21.0987 M=1 R=7.46667
+ SA=75002.2 SB=75004.3 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1022_d N_C_M1009_g N_A_199_294#_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.203679 AS=0.15 PD=1.43396 PS=1.3 NRD=20.685 NRS=1.9503 M=1 R=6.66667
+ SA=75002.8 SB=75004.3 A=0.15 P=2.3 MULT=1
MM1006 N_A_199_294#_M1009_s N_D_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.1925 PD=1.3 PS=1.385 NRD=1.9503 NRS=18.715 M=1 R=6.66667
+ SA=75003.2 SB=75003.8 A=0.15 P=2.3 MULT=1
MM1018 N_A_199_294#_M1018_d N_D_M1018_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.43 AS=0.1925 PD=1.86 PS=1.385 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75003.8 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_C_M1011_g N_A_199_294#_M1018_d VPB PHIGHVT L=0.15 W=1
+ AD=0.16 AS=0.43 PD=1.32 PS=1.86 NRD=3.9203 NRS=1.9503 M=1 R=6.66667 SA=75004.8
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1001 N_A_199_294#_M1001_d N_B_M1001_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.16 PD=1.3 PS=1.32 NRD=1.9503 NRS=3.9203 M=1 R=6.66667 SA=75005.2
+ SB=75001.8 A=0.15 P=2.3 MULT=1
MM1002 N_A_199_294#_M1001_d N_A_27_368#_M1002_g N_VPWR_M1002_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75005.7 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1024 N_A_199_294#_M1024_d N_A_27_368#_M1024_g N_VPWR_M1002_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75006.1 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1010 N_A_199_294#_M1024_d N_B_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.53 PD=1.3 PS=3.06 NRD=1.9503 NRS=24.6053 M=1 R=6.66667 SA=75006.6
+ SB=75000.5 A=0.15 P=2.3 MULT=1
DX26_noxref VNB VPB NWDIODE A=14.9916 P=19.84
c_80 VNB 0 5.40706e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__and4b_4.pxi.spice"
*
.ends
*
*
