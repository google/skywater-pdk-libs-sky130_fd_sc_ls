* File: sky130_fd_sc_ls__dlrtn_1.pex.spice
* Created: Fri Aug 28 13:18:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DLRTN_1%D 3 5 7 8
c26 5 0 1.54286e-19 $X=0.51 $Y=1.895
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.615 $X2=0.6 $Y2=1.615
r28 8 12 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.72 $Y=1.615 $X2=0.6
+ $Y2=1.615
r29 5 11 56.8989 $w=3.02e-07 $l=3.18371e-07 $layer=POLY_cond $X=0.51 $Y=1.895
+ $X2=0.592 $Y2=1.615
r30 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.51 $Y=1.895 $X2=0.51
+ $Y2=2.39
r31 1 11 38.5446 $w=3.02e-07 $l=2.07918e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.592 $Y2=1.615
r32 1 3 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_1%GATE_N 3 5 7 8
r34 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r35 5 11 57.6553 $w=2.91e-07 $l=2.99333e-07 $layer=POLY_cond $X=1.13 $Y=1.895
+ $X2=1.17 $Y2=1.615
r36 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.13 $Y=1.895 $X2=1.13
+ $Y2=2.39
r37 1 11 38.6072 $w=2.91e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.085 $Y=1.45
+ $X2=1.17 $Y2=1.615
r38 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.085 $Y=1.45
+ $X2=1.085 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_1%A_232_98# 1 2 7 9 12 16 19 20 22 24 27 29 34
+ 35 37 38 41 45 46
c123 27 0 1.46239e-19 $X=3.875 $Y=1.805
r124 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.505 $X2=1.74 $Y2=1.505
r125 45 46 9.42615 $w=4.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.432 $Y=2.115
+ $X2=1.432 $Y2=1.95
r126 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.08
+ $Y=2.195 $X2=4.08 $Y2=2.195
r127 39 41 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.08 $Y=2.52
+ $X2=4.08 $Y2=2.195
r128 37 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.915 $Y=2.605
+ $X2=4.08 $Y2=2.52
r129 37 38 146.139 $w=1.68e-07 $l=2.24e-06 $layer=LI1_cond $X=3.915 $Y=2.605
+ $X2=1.675 $Y2=2.605
r130 35 49 9.11389 $w=2.71e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.59 $Y=1.67
+ $X2=1.675 $Y2=1.505
r131 35 46 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.59 $Y=1.67
+ $X2=1.59 $Y2=1.95
r132 34 38 9.10402 $w=1.7e-07 $l=2.82319e-07 $layer=LI1_cond $X=1.432 $Y=2.52
+ $X2=1.675 $Y2=2.605
r133 33 45 1.89893 $w=4.83e-07 $l=7.7e-08 $layer=LI1_cond $X=1.432 $Y=2.192
+ $X2=1.432 $Y2=2.115
r134 33 34 8.08894 $w=4.83e-07 $l=3.28e-07 $layer=LI1_cond $X=1.432 $Y=2.192
+ $X2=1.432 $Y2=2.52
r135 29 49 18.9077 $w=2.71e-07 $l=4.2e-07 $layer=LI1_cond $X=1.675 $Y=1.085
+ $X2=1.675 $Y2=1.505
r136 29 31 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.505 $Y=1.085
+ $X2=1.3 $Y2=1.085
r137 25 27 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=3.72 $Y=1.805
+ $X2=3.875 $Y2=1.805
r138 24 50 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=2.065 $Y=1.505
+ $X2=1.74 $Y2=1.505
r139 20 42 52.5187 $w=3.81e-07 $l=3.29454e-07 $layer=POLY_cond $X=3.89 $Y=2.465
+ $X2=4.022 $Y2=2.195
r140 20 22 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.89 $Y=2.465
+ $X2=3.89 $Y2=2.75
r141 19 42 39.2352 $w=3.81e-07 $l=2.26892e-07 $layer=POLY_cond $X=3.875 $Y=2.03
+ $X2=4.022 $Y2=2.195
r142 18 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.875 $Y=1.88
+ $X2=3.875 $Y2=1.805
r143 18 19 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.875 $Y=1.88
+ $X2=3.875 $Y2=2.03
r144 14 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.72 $Y=1.73
+ $X2=3.72 $Y2=1.805
r145 14 16 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=3.72 $Y=1.73
+ $X2=3.72 $Y2=0.69
r146 10 24 43.4747 $w=1.95e-07 $l=1.85257e-07 $layer=POLY_cond $X=2.225 $Y=1.34
+ $X2=2.182 $Y2=1.505
r147 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.225 $Y=1.34
+ $X2=2.225 $Y2=0.78
r148 7 24 96.6183 $w=1.95e-07 $l=3.93268e-07 $layer=POLY_cond $X=2.155 $Y=1.885
+ $X2=2.182 $Y2=1.505
r149 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.155 $Y=1.885
+ $X2=2.155 $Y2=2.38
r150 2 45 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.205
+ $Y=1.97 $X2=1.355 $Y2=2.115
r151 1 31 182 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.49 $X2=1.3 $Y2=1.035
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_1%A_27_136# 1 2 7 8 9 11 12 14 16 20 25 26 29
+ 32 34 35
c81 35 0 1.54286e-19 $X=0.272 $Y=1.95
c82 7 0 7.69973e-20 $X=2.775 $Y=1.59
r83 34 35 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.272 $Y=2.115
+ $X2=0.272 $Y2=1.95
r84 32 35 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.18 $Y=1.25 $X2=0.18
+ $Y2=1.95
r85 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.7
+ $Y=1.425 $X2=2.7 $Y2=1.425
r86 27 29 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.7 $Y=0.75 $X2=2.7
+ $Y2=1.425
r87 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.535 $Y=0.665
+ $X2=2.7 $Y2=0.75
r88 25 26 136.353 $w=1.68e-07 $l=2.09e-06 $layer=LI1_cond $X=2.535 $Y=0.665
+ $X2=0.445 $Y2=0.665
r89 18 32 8.81775 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=0.27 $Y=1.075
+ $X2=0.27 $Y2=1.25
r90 18 20 3.95123 $w=3.48e-07 $l=1.2e-07 $layer=LI1_cond $X=0.27 $Y=1.075
+ $X2=0.27 $Y2=0.955
r91 17 26 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=0.27 $Y=0.75
+ $X2=0.445 $Y2=0.665
r92 17 20 6.75002 $w=3.48e-07 $l=2.05e-07 $layer=LI1_cond $X=0.27 $Y=0.75
+ $X2=0.27 $Y2=0.955
r93 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.33 $Y=1.085
+ $X2=3.33 $Y2=0.69
r94 13 30 47.839 $w=2.67e-07 $l=3.37565e-07 $layer=POLY_cond $X=2.865 $Y=1.16
+ $X2=2.7 $Y2=1.425
r95 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.255 $Y=1.16
+ $X2=3.33 $Y2=1.085
r96 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.255 $Y=1.16
+ $X2=2.865 $Y2=1.16
r97 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.775 $Y=1.885
+ $X2=2.775 $Y2=2.46
r98 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.775 $Y=1.795 $X2=2.775
+ $Y2=1.885
r99 7 30 34.9261 $w=2.67e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.775 $Y=1.59
+ $X2=2.7 $Y2=1.425
r100 7 8 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=2.775 $Y=1.59
+ $X2=2.775 $Y2=1.795
r101 2 34 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=1.97 $X2=0.285 $Y2=2.115
r102 1 20 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.68 $X2=0.28 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_1%A_357_392# 1 2 7 9 12 15 16 21 23 25 26 31
+ 37
c94 31 0 7.69973e-20 $X=2.16 $Y=1.045
c95 25 0 1.0947e-19 $X=4.17 $Y=1.355
c96 16 0 1.46239e-19 $X=3.075 $Y=1.925
r97 36 37 7.70264 $w=5.08e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=2.095
+ $X2=2.245 $Y2=2.095
r98 34 36 5.39408 $w=5.08e-07 $l=2.3e-07 $layer=LI1_cond $X=1.93 $Y=2.095
+ $X2=2.16 $Y2=2.095
r99 29 31 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.01 $Y=1.045
+ $X2=2.16 $Y2=1.045
r100 26 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.17 $Y=1.355
+ $X2=4.17 $Y2=1.19
r101 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.17
+ $Y=1.355 $X2=4.17 $Y2=1.355
r102 23 25 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=3.405 $Y=1.355
+ $X2=4.17 $Y2=1.355
r103 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.24
+ $Y=1.61 $X2=3.24 $Y2=1.61
r104 19 21 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.24 $Y=1.84
+ $X2=3.24 $Y2=1.61
r105 18 23 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=3.24 $Y=1.52
+ $X2=3.405 $Y2=1.355
r106 18 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.24 $Y=1.52 $X2=3.24
+ $Y2=1.61
r107 16 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.075 $Y=1.925
+ $X2=3.24 $Y2=1.84
r108 16 37 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.075 $Y=1.925
+ $X2=2.245 $Y2=1.925
r109 15 36 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.16 $Y=1.84
+ $X2=2.16 $Y2=2.095
r110 14 31 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.16 $Y=1.17
+ $X2=2.16 $Y2=1.045
r111 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.16 $Y=1.17
+ $X2=2.16 $Y2=1.84
r112 12 40 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.195 $Y=0.58
+ $X2=4.195 $Y2=1.19
r113 7 22 56.7567 $w=2.92e-07 $l=2.96648e-07 $layer=POLY_cond $X=3.195 $Y=1.885
+ $X2=3.24 $Y2=1.61
r114 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.195 $Y=1.885
+ $X2=3.195 $Y2=2.46
r115 2 34 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=1.785
+ $Y=1.96 $X2=1.93 $Y2=2.145
r116 1 29 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.41 $X2=2.01 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_1%A_897_406# 1 2 7 9 12 15 18 20 22 24 25 32
+ 38 40 41 42 47 50
c112 42 0 4.25141e-20 $X=5.715 $Y=1.72
c113 38 0 1.23233e-19 $X=6.415 $Y=1.805
c114 25 0 1.40957e-19 $X=5.465 $Y=2.195
c115 20 0 1.72324e-19 $X=6.695 $Y=1.765
c116 15 0 1.0947e-19 $X=4.65 $Y=2.03
r117 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.61
+ $Y=1.485 $X2=6.61 $Y2=1.485
r118 45 47 3.46863 $w=4.98e-07 $l=1.45e-07 $layer=LI1_cond $X=5.715 $Y=2.195
+ $X2=5.715 $Y2=2.34
r119 44 45 5.02353 $w=4.98e-07 $l=2.1e-07 $layer=LI1_cond $X=5.715 $Y=1.985
+ $X2=5.715 $Y2=2.195
r120 41 44 4.30588 $w=4.98e-07 $l=1.8e-07 $layer=LI1_cond $X=5.715 $Y=1.805
+ $X2=5.715 $Y2=1.985
r121 41 42 7.60339 $w=4.98e-07 $l=8.5e-08 $layer=LI1_cond $X=5.715 $Y=1.805
+ $X2=5.715 $Y2=1.72
r122 40 42 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.55 $Y=1.13
+ $X2=5.55 $Y2=1.72
r123 39 41 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=5.965 $Y=1.805
+ $X2=5.715 $Y2=1.805
r124 38 50 13.9429 $w=2.8e-07 $l=4e-07 $layer=LI1_cond $X=6.415 $Y=1.805
+ $X2=6.595 $Y2=1.485
r125 38 39 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.415 $Y=1.805
+ $X2=5.965 $Y2=1.805
r126 30 40 9.56083 $w=3.93e-07 $l=1.97e-07 $layer=LI1_cond $X=5.437 $Y=0.933
+ $X2=5.437 $Y2=1.13
r127 30 32 12.1955 $w=3.93e-07 $l=4.18e-07 $layer=LI1_cond $X=5.437 $Y=0.933
+ $X2=5.437 $Y2=0.515
r128 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.65
+ $Y=2.195 $X2=4.65 $Y2=2.195
r129 25 45 3.16914 $w=3.3e-07 $l=2.5e-07 $layer=LI1_cond $X=5.465 $Y=2.195
+ $X2=5.715 $Y2=2.195
r130 25 27 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=5.465 $Y=2.195
+ $X2=4.65 $Y2=2.195
r131 23 24 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=4.635 $Y=1.34
+ $X2=4.635 $Y2=1.49
r132 20 51 57.1617 $w=2.98e-07 $l=3.1749e-07 $layer=POLY_cond $X=6.695 $Y=1.765
+ $X2=6.615 $Y2=1.485
r133 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.695 $Y=1.765
+ $X2=6.695 $Y2=2.4
r134 16 51 38.561 $w=2.98e-07 $l=1.72337e-07 $layer=POLY_cond $X=6.6 $Y=1.32
+ $X2=6.615 $Y2=1.485
r135 16 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.6 $Y=1.32 $X2=6.6
+ $Y2=0.74
r136 15 28 38.5916 $w=2.93e-07 $l=1.65e-07 $layer=POLY_cond $X=4.65 $Y=2.03
+ $X2=4.65 $Y2=2.195
r137 15 24 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=4.65 $Y=2.03
+ $X2=4.65 $Y2=1.49
r138 12 23 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.62 $Y=0.58
+ $X2=4.62 $Y2=1.34
r139 7 28 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=4.575 $Y=2.465
+ $X2=4.65 $Y2=2.195
r140 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.575 $Y=2.465
+ $X2=4.575 $Y2=2.75
r141 2 47 300 $w=1.7e-07 $l=6.06218e-07 $layer=licon1_PDIFF $count=2 $X=5.565
+ $Y=1.84 $X2=5.8 $Y2=2.34
r142 2 44 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.84 $X2=5.8 $Y2=1.985
r143 1 32 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.26
+ $Y=0.37 $X2=5.405 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_1%A_654_392# 1 2 7 8 9 11 12 14 17 19 24 25 26
+ 29 31 32 34 36 37
c107 17 0 3.19186e-20 $X=5.13 $Y=1.575
c108 9 0 9.13148e-20 $X=5.49 $Y=1.765
c109 8 0 1.70198e-19 $X=5.295 $Y=1.26
c110 7 0 1.40957e-19 $X=5.545 $Y=1.26
r111 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.13
+ $Y=1.465 $X2=5.13 $Y2=1.465
r112 34 36 8.97739 $w=3.02e-07 $l=2.13787e-07 $layer=LI1_cond $X=4.985 $Y=1.3
+ $X2=5.097 $Y2=1.465
r113 33 34 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.985 $Y=1.02
+ $X2=4.985 $Y2=1.3
r114 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.9 $Y=0.935
+ $X2=4.985 $Y2=1.02
r115 31 32 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.9 $Y=0.935
+ $X2=4.145 $Y2=0.935
r116 27 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.98 $Y=0.85
+ $X2=4.145 $Y2=0.935
r117 27 29 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=3.98 $Y=0.85
+ $X2=3.98 $Y2=0.58
r118 25 36 12.5232 $w=3.02e-07 $l=3.96447e-07 $layer=LI1_cond $X=4.9 $Y=1.775
+ $X2=5.097 $Y2=1.465
r119 25 26 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=4.9 $Y=1.775
+ $X2=3.745 $Y2=1.775
r120 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.66 $Y=1.86
+ $X2=3.745 $Y2=1.775
r121 23 24 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.66 $Y=1.86
+ $X2=3.66 $Y2=2.18
r122 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.575 $Y=2.265
+ $X2=3.66 $Y2=2.18
r123 19 21 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.575 $Y=2.265
+ $X2=3.425 $Y2=2.265
r124 17 37 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=5.13 $Y=1.575
+ $X2=5.13 $Y2=1.465
r125 17 18 107.776 $w=1.61e-07 $l=3.6e-07 $layer=POLY_cond $X=5.13 $Y=1.67
+ $X2=5.49 $Y2=1.67
r126 15 37 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=5.13 $Y=1.335
+ $X2=5.13 $Y2=1.465
r127 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.62 $Y=1.185
+ $X2=5.62 $Y2=0.74
r128 9 18 4.52116 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=5.49 $Y=1.765
+ $X2=5.49 $Y2=1.67
r129 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.49 $Y=1.765
+ $X2=5.49 $Y2=2.34
r130 8 15 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.295 $Y=1.26
+ $X2=5.13 $Y2=1.335
r131 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.545 $Y=1.26
+ $X2=5.62 $Y2=1.185
r132 7 8 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.545 $Y=1.26
+ $X2=5.295 $Y2=1.26
r133 2 21 600 $w=1.7e-07 $l=3.74566e-07 $layer=licon1_PDIFF $count=1 $X=3.27
+ $Y=1.96 $X2=3.425 $Y2=2.265
r134 1 29 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=3.795
+ $Y=0.37 $X2=3.98 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_1%RESET_B 1 3 4 6 7
c34 1 0 4.25141e-20 $X=6.01 $Y=1.22
r35 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.07
+ $Y=1.385 $X2=6.07 $Y2=1.385
r36 7 11 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=6.06 $Y=1.295 $X2=6.06
+ $Y2=1.385
r37 4 10 77.2841 $w=2.7e-07 $l=3.995e-07 $layer=POLY_cond $X=6.11 $Y=1.765
+ $X2=6.07 $Y2=1.385
r38 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.11 $Y=1.765
+ $X2=6.11 $Y2=2.34
r39 1 10 38.9026 $w=2.7e-07 $l=1.92678e-07 $layer=POLY_cond $X=6.01 $Y=1.22
+ $X2=6.07 $Y2=1.385
r40 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.01 $Y=1.22 $X2=6.01
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_1%VPWR 1 2 3 4 17 21 25 30 31 32 41 48 55 56
+ 59 62 69
r71 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r72 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r73 56 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r74 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r75 53 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.42 $Y2=3.33
r76 53 55 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.96 $Y2=3.33
r77 52 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r78 52 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.04
+ $Y2=3.33
r79 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r80 49 51 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.43 $Y=3.33 $X2=6
+ $Y2=3.33
r81 48 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=3.33
+ $X2=6.42 $Y2=3.33
r82 48 51 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.255 $Y=3.33 $X2=6
+ $Y2=3.33
r83 47 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r84 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r85 43 46 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r86 43 44 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r87 41 49 10.1669 $w=1.7e-07 $l=3.98e-07 $layer=LI1_cond $X=5.032 $Y=3.33
+ $X2=5.43 $Y2=3.33
r88 41 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r89 41 62 9.55358 $w=7.93e-07 $l=6.35e-07 $layer=LI1_cond $X=5.032 $Y=3.33
+ $X2=5.032 $Y2=2.695
r90 41 46 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.635 $Y=3.33
+ $X2=4.56 $Y2=3.33
r91 40 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r92 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r93 37 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r94 37 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r95 36 39 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r96 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r97 34 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.82 $Y2=3.33
r98 34 36 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.2 $Y2=3.33
r99 32 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r100 32 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 30 39 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.3 $Y=3.33
+ $X2=2.16 $Y2=3.33
r102 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.3 $Y=3.33
+ $X2=2.465 $Y2=3.33
r103 29 43 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.63 $Y=3.33
+ $X2=2.64 $Y2=3.33
r104 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=3.33
+ $X2=2.465 $Y2=3.33
r105 25 28 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.42 $Y=2.145
+ $X2=6.42 $Y2=2.825
r106 23 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=3.245
+ $X2=6.42 $Y2=3.33
r107 23 28 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=6.42 $Y=3.245
+ $X2=6.42 $Y2=2.825
r108 19 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=3.245
+ $X2=2.465 $Y2=3.33
r109 19 21 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.465 $Y=3.245
+ $X2=2.465 $Y2=2.945
r110 15 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=3.33
r111 15 17 39.4624 $w=3.28e-07 $l=1.13e-06 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=2.115
r112 4 28 600 $w=1.7e-07 $l=1.09622e-06 $layer=licon1_PDIFF $count=1 $X=6.185
+ $Y=1.84 $X2=6.42 $Y2=2.825
r113 4 25 300 $w=1.7e-07 $l=4.05832e-07 $layer=licon1_PDIFF $count=2 $X=6.185
+ $Y=1.84 $X2=6.42 $Y2=2.145
r114 3 62 300 $w=1.7e-07 $l=6.8815e-07 $layer=licon1_PDIFF $count=2 $X=4.65
+ $Y=2.54 $X2=5.265 $Y2=2.695
r115 2 21 600 $w=1.7e-07 $l=1.09622e-06 $layer=licon1_PDIFF $count=1 $X=2.23
+ $Y=1.96 $X2=2.465 $Y2=2.945
r116 1 17 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.97 $X2=0.82 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_1%Q 1 2 9 13 14 15 16 23 32
r22 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=6.935 $Y=2 $X2=6.935
+ $Y2=2.035
r23 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=6.935 $Y=2.405
+ $X2=6.935 $Y2=2.775
r24 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=6.935 $Y=1.975
+ $X2=6.935 $Y2=2
r25 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=6.935 $Y=1.975
+ $X2=6.935 $Y2=1.82
r26 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=6.935 $Y=2.06
+ $X2=6.935 $Y2=2.405
r27 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=6.935 $Y=2.06
+ $X2=6.935 $Y2=2.035
r28 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.03 $Y=1.13 $X2=7.03
+ $Y2=1.82
r29 7 13 9.39714 $w=3.83e-07 $l=1.92e-07 $layer=LI1_cond $X=6.922 $Y=0.938
+ $X2=6.922 $Y2=1.13
r30 7 9 12.6619 $w=3.83e-07 $l=4.23e-07 $layer=LI1_cond $X=6.922 $Y=0.938
+ $X2=6.922 $Y2=0.515
r31 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=1.84 $X2=6.92 $Y2=1.985
r32 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=1.84 $X2=6.92 $Y2=2.815
r33 1 9 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=6.675
+ $Y=0.37 $X2=6.895 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTN_1%VGND 1 2 3 4 15 19 22 23 25 26 27 29 53 54
+ 58 66 72
c67 19 0 1.72324e-19 $X=6.305 $Y=0.49
c68 15 0 1.70198e-19 $X=4.84 $Y=0.515
r69 70 72 7.43269 $w=4.93e-07 $l=8e-08 $layer=LI1_cond $X=3.12 $Y=0.162 $X2=3.2
+ $Y2=0.162
r70 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r71 68 70 2.05387 $w=4.93e-07 $l=8.5e-08 $layer=LI1_cond $X=3.035 $Y=0.162
+ $X2=3.12 $Y2=0.162
r72 65 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r73 64 68 9.54446 $w=4.93e-07 $l=3.95e-07 $layer=LI1_cond $X=2.64 $Y=0.162
+ $X2=3.035 $Y2=0.162
r74 64 66 12.3861 $w=4.93e-07 $l=2.85e-07 $layer=LI1_cond $X=2.64 $Y=0.162
+ $X2=2.355 $Y2=0.162
r75 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r76 58 61 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.79
+ $Y2=0.325
r77 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r78 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r79 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r80 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r81 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r82 47 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6 $Y2=0
r83 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r84 45 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r85 44 72 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=3.2
+ $Y2=0
r86 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r87 41 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r88 40 66 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.355
+ $Y2=0
r89 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r90 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r91 38 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r92 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r93 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r94 35 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r95 35 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r96 32 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r97 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r98 29 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r99 29 31 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.24
+ $Y2=0
r100 27 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r101 27 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r102 25 50 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=6
+ $Y2=0
r103 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=6.305
+ $Y2=0
r104 24 53 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=6.47 $Y=0 $X2=6.96
+ $Y2=0
r105 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.47 $Y=0 $X2=6.305
+ $Y2=0
r106 22 44 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.67 $Y=0 $X2=4.56
+ $Y2=0
r107 22 23 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.67 $Y=0 $X2=4.84
+ $Y2=0
r108 21 47 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=5.01 $Y=0 $X2=5.04
+ $Y2=0
r109 21 23 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.01 $Y=0 $X2=4.84
+ $Y2=0
r110 17 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.305 $Y=0.085
+ $X2=6.305 $Y2=0
r111 17 19 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=6.305 $Y=0.085
+ $X2=6.305 $Y2=0.49
r112 13 23 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.84 $Y=0.085
+ $X2=4.84 $Y2=0
r113 13 15 14.575 $w=3.38e-07 $l=4.3e-07 $layer=LI1_cond $X=4.84 $Y=0.085
+ $X2=4.84 $Y2=0.515
r114 4 19 91 $w=1.7e-07 $l=2.73496e-07 $layer=licon1_NDIFF $count=2 $X=6.085
+ $Y=0.37 $X2=6.305 $Y2=0.49
r115 3 15 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.695
+ $Y=0.37 $X2=4.84 $Y2=0.515
r116 2 68 91 $w=1.7e-07 $l=7.76338e-07 $layer=licon1_NDIFF $count=2 $X=2.3
+ $Y=0.41 $X2=3.035 $Y2=0.325
r117 1 61 182 $w=1.7e-07 $l=4.51802e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.68 $X2=0.79 $Y2=0.325
.ends

