* File: sky130_fd_sc_ls__bufbuf_16.spice
* Created: Fri Aug 28 13:07:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__bufbuf_16.pex.spice"
.subckt sky130_fd_sc_ls__bufbuf_16  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1049 N_VGND_M1049_d N_A_M1049_g N_A_27_368#_M1049_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1025 N_VGND_M1049_d N_A_27_368#_M1025_g N_A_203_74#_M1025_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1029 N_VGND_M1029_d N_A_27_368#_M1029_g N_A_203_74#_M1025_s VNB NSHORT L=0.15
+ W=0.74 AD=0.10545 AS=0.1036 PD=1.025 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1050 N_VGND_M1029_d N_A_27_368#_M1050_g N_A_203_74#_M1050_s VNB NSHORT L=0.15
+ W=0.74 AD=0.10545 AS=0.2109 PD=1.025 PS=2.05 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_588_74#_M1000_d N_A_203_74#_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.3 SB=75009.8 A=0.111 P=1.78 MULT=1
MM1006 N_A_588_74#_M1000_d N_A_203_74#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75009.4 A=0.111 P=1.78 MULT=1
MM1023 N_A_588_74#_M1023_d N_A_203_74#_M1023_g N_VGND_M1006_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.2 SB=75008.9 A=0.111 P=1.78 MULT=1
MM1027 N_A_588_74#_M1023_d N_A_203_74#_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75008.4 A=0.111 P=1.78 MULT=1
MM1041 N_A_588_74#_M1041_d N_A_203_74#_M1041_g N_VGND_M1027_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75002.1 SB=75007.9 A=0.111 P=1.78 MULT=1
MM1048 N_A_588_74#_M1041_d N_A_203_74#_M1048_g N_VGND_M1048_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.6 SB=75007.5 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1048_s N_A_588_74#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003
+ SB=75007.1 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A_588_74#_M1004_g N_X_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.4
+ SB=75006.7 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1004_d N_A_588_74#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.9
+ SB=75006.2 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A_588_74#_M1011_g N_X_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.3
+ SB=75005.8 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1011_d N_A_588_74#_M1012_g N_X_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.7
+ SB=75005.4 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_588_74#_M1013_g N_X_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.1
+ SB=75004.9 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1013_d N_A_588_74#_M1014_g N_X_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75005.6
+ SB=75004.4 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_A_588_74#_M1018_g N_X_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.1
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1018_d N_A_588_74#_M1021_g N_X_M1021_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75006.6
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1022_d N_A_588_74#_M1022_g N_X_M1021_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75007
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1022_d N_A_588_74#_M1024_g N_X_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75007.5
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1034 N_VGND_M1034_d N_A_588_74#_M1034_g N_X_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75007.9
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1037 N_VGND_M1034_d N_A_588_74#_M1037_g N_X_M1037_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75008.4
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1040 N_VGND_M1040_d N_A_588_74#_M1040_g N_X_M1037_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1332 AS=0.1036 PD=1.1 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75008.9
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1042 N_VGND_M1040_d N_A_588_74#_M1042_g N_X_M1042_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1332 AS=0.1036 PD=1.1 PS=1.02 NRD=12.972 NRS=0 M=1 R=4.93333 SA=75009.4
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1045 N_VGND_M1045_d N_A_588_74#_M1045_g N_X_M1042_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75009.8
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1030 N_VPWR_M1030_d N_A_M1030_g N_A_27_368#_M1030_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1001 N_A_203_74#_M1001_d N_A_27_368#_M1001_g N_VPWR_M1030_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1031 N_A_203_74#_M1001_d N_A_27_368#_M1031_g N_VPWR_M1031_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1043 N_A_203_74#_M1043_d N_A_27_368#_M1043_g N_VPWR_M1031_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_A_203_74#_M1005_g N_A_588_74#_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75009.8 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1016_d N_A_203_74#_M1016_g N_A_588_74#_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75009.3 A=0.168 P=2.54 MULT=1
MM1028 N_VPWR_M1016_d N_A_203_74#_M1028_g N_A_588_74#_M1028_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75008.9 A=0.168 P=2.54 MULT=1
MM1032 N_VPWR_M1032_d N_A_203_74#_M1032_g N_A_588_74#_M1028_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.1736 AS=0.168 PD=1.43 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75008.4 A=0.168 P=2.54 MULT=1
MM1036 N_VPWR_M1032_d N_A_203_74#_M1036_g N_A_588_74#_M1036_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.1736 AS=0.168 PD=1.43 PS=1.42 NRD=3.5066 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75008 A=0.168 P=2.54 MULT=1
MM1046 N_VPWR_M1046_d N_A_203_74#_M1046_g N_A_588_74#_M1036_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.1736 AS=0.168 PD=1.43 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75007.5 A=0.168 P=2.54 MULT=1
MM1003 N_X_M1003_d N_A_588_74#_M1003_g N_VPWR_M1046_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.1736 PD=1.42 PS=1.43 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75002.9 SB=75007.1 A=0.168 P=2.54 MULT=1
MM1008 N_X_M1003_d N_A_588_74#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.4 SB=75006.6 A=0.168 P=2.54 MULT=1
MM1009 N_X_M1009_d N_A_588_74#_M1009_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.9 SB=75006.1 A=0.168 P=2.54 MULT=1
MM1010 N_X_M1009_d N_A_588_74#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.3 SB=75005.7 A=0.168 P=2.54 MULT=1
MM1015 N_X_M1015_d N_A_588_74#_M1015_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.8 SB=75005.2 A=0.168 P=2.54 MULT=1
MM1017 N_X_M1015_d N_A_588_74#_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.2 SB=75004.8 A=0.168 P=2.54 MULT=1
MM1019 N_X_M1019_d N_A_588_74#_M1019_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.7 SB=75004.3 A=0.168 P=2.54 MULT=1
MM1020 N_X_M1019_d N_A_588_74#_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.1 SB=75003.9 A=0.168 P=2.54 MULT=1
MM1026 N_X_M1026_d N_A_588_74#_M1026_g N_VPWR_M1020_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.6 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1033 N_X_M1026_d N_A_588_74#_M1033_g N_VPWR_M1033_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75007
+ SB=75003 A=0.168 P=2.54 MULT=1
MM1035 N_X_M1035_d N_A_588_74#_M1035_g N_VPWR_M1033_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.5 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1038 N_X_M1035_d N_A_588_74#_M1038_g N_VPWR_M1038_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.9 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1039 N_X_M1039_d N_A_588_74#_M1039_g N_VPWR_M1038_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75008.4 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1044 N_X_M1039_d N_A_588_74#_M1044_g N_VPWR_M1044_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75008.8 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1047 N_X_M1047_d N_A_588_74#_M1047_g N_VPWR_M1044_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75009.3 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1051 N_X_M1047_d N_A_588_74#_M1051_g N_VPWR_M1051_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.3304 PD=1.47 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75009.8 SB=75000.2 A=0.168 P=2.54 MULT=1
DX52_noxref VNB VPB NWDIODE A=24.8124 P=30.4
c_120 VNB 0 1.53678e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__bufbuf_16.pxi.spice"
*
.ends
*
*
