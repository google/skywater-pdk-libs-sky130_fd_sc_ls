* File: sky130_fd_sc_ls__o2111ai_1.pxi.spice
* Created: Wed Sep  2 11:16:49 2020
* 
x_PM_SKY130_FD_SC_LS__O2111AI_1%D1 N_D1_c_49_n N_D1_M1003_g N_D1_c_50_n
+ N_D1_M1006_g D1 PM_SKY130_FD_SC_LS__O2111AI_1%D1
x_PM_SKY130_FD_SC_LS__O2111AI_1%C1 N_C1_c_74_n N_C1_M1007_g N_C1_c_75_n
+ N_C1_M1005_g C1 C1 C1 PM_SKY130_FD_SC_LS__O2111AI_1%C1
x_PM_SKY130_FD_SC_LS__O2111AI_1%B1 N_B1_c_108_n N_B1_M1001_g N_B1_c_109_n
+ N_B1_M1000_g B1 N_B1_c_110_n PM_SKY130_FD_SC_LS__O2111AI_1%B1
x_PM_SKY130_FD_SC_LS__O2111AI_1%A2 N_A2_c_137_n N_A2_M1002_g N_A2_c_138_n
+ N_A2_M1008_g A2 PM_SKY130_FD_SC_LS__O2111AI_1%A2
x_PM_SKY130_FD_SC_LS__O2111AI_1%A1 N_A1_c_166_n N_A1_M1009_g N_A1_c_167_n
+ N_A1_M1004_g A1 PM_SKY130_FD_SC_LS__O2111AI_1%A1
x_PM_SKY130_FD_SC_LS__O2111AI_1%VPWR N_VPWR_M1003_s N_VPWR_M1005_d
+ N_VPWR_M1009_d N_VPWR_c_190_n N_VPWR_c_191_n N_VPWR_c_192_n N_VPWR_c_193_n
+ N_VPWR_c_194_n N_VPWR_c_195_n VPWR N_VPWR_c_196_n N_VPWR_c_197_n
+ N_VPWR_c_198_n N_VPWR_c_189_n PM_SKY130_FD_SC_LS__O2111AI_1%VPWR
x_PM_SKY130_FD_SC_LS__O2111AI_1%Y N_Y_M1006_s N_Y_M1003_d N_Y_M1000_d
+ N_Y_c_229_n N_Y_c_232_n N_Y_c_233_n N_Y_c_234_n N_Y_c_235_n N_Y_c_230_n
+ N_Y_c_236_n Y Y Y N_Y_c_237_n PM_SKY130_FD_SC_LS__O2111AI_1%Y
x_PM_SKY130_FD_SC_LS__O2111AI_1%A_368_74# N_A_368_74#_M1001_d
+ N_A_368_74#_M1004_d N_A_368_74#_c_285_n N_A_368_74#_c_282_n
+ N_A_368_74#_c_283_n N_A_368_74#_c_284_n
+ PM_SKY130_FD_SC_LS__O2111AI_1%A_368_74#
x_PM_SKY130_FD_SC_LS__O2111AI_1%VGND N_VGND_M1002_d N_VGND_c_310_n VGND
+ N_VGND_c_311_n N_VGND_c_312_n N_VGND_c_313_n N_VGND_c_314_n
+ PM_SKY130_FD_SC_LS__O2111AI_1%VGND
cc_1 VNB N_D1_c_49_n 0.042283f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.765
cc_2 VNB N_D1_c_50_n 0.0217968f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.22
cc_3 VNB D1 0.00350742f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_C1_c_74_n 0.0172466f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.765
cc_5 VNB N_C1_c_75_n 0.0372066f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.22
cc_6 VNB C1 0.00553803f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB N_B1_c_108_n 0.0190408f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.765
cc_8 VNB N_B1_c_109_n 0.0343061f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.22
cc_9 VNB N_B1_c_110_n 0.0102576f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.385
cc_10 VNB N_A2_c_137_n 0.0186396f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.765
cc_11 VNB N_A2_c_138_n 0.035316f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.22
cc_12 VNB A2 0.0144016f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_13 VNB N_A1_c_166_n 0.06837f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.765
cc_14 VNB N_A1_c_167_n 0.0247091f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.22
cc_15 VNB A1 0.00922063f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_16 VNB N_VPWR_c_189_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_229_n 0.0309816f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.385
cc_18 VNB N_Y_c_230_n 0.0331431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_368_74#_c_282_n 0.00289626f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.385
cc_20 VNB N_A_368_74#_c_283_n 0.00716806f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.385
cc_21 VNB N_A_368_74#_c_284_n 0.021252f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.385
cc_22 VNB N_VGND_c_310_n 0.00739995f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.74
cc_23 VNB N_VGND_c_311_n 0.0659727f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.385
cc_24 VNB N_VGND_c_312_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_313_n 0.219739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_314_n 0.00786346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VPB N_D1_c_49_n 0.0242032f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.765
cc_28 VPB N_C1_c_75_n 0.0234011f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.22
cc_29 VPB N_B1_c_109_n 0.0237827f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.22
cc_30 VPB N_A2_c_138_n 0.0231209f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.22
cc_31 VPB N_A1_c_166_n 0.029309f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.765
cc_32 VPB N_VPWR_c_190_n 0.0476314f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.295
cc_33 VPB N_VPWR_c_191_n 0.00980878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_192_n 0.012808f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_193_n 0.0559106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_194_n 0.0142356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_195_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_196_n 0.0212158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_197_n 0.0314247f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_198_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_189_n 0.0818387f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_Y_c_229_n 0.00311325f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.385
cc_43 VPB N_Y_c_232_n 0.0157847f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.295
cc_44 VPB N_Y_c_233_n 0.0148348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_Y_c_234_n 0.0165547f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_Y_c_235_n 0.00290171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_Y_c_236_n 0.00785442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_Y_c_237_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 N_D1_c_50_n N_C1_c_74_n 0.0499419f $X=0.835 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_50 N_D1_c_49_n N_C1_c_75_n 0.042231f $X=0.82 $Y=1.765 $X2=0 $Y2=0
cc_51 D1 N_C1_c_75_n 3.85374e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_52 N_D1_c_50_n C1 0.0100911f $X=0.835 $Y=1.22 $X2=0 $Y2=0
cc_53 D1 C1 0.028682f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_54 N_D1_c_49_n N_VPWR_c_190_n 0.0227729f $X=0.82 $Y=1.765 $X2=0 $Y2=0
cc_55 N_D1_c_49_n N_VPWR_c_196_n 0.00445602f $X=0.82 $Y=1.765 $X2=0 $Y2=0
cc_56 N_D1_c_49_n N_VPWR_c_189_n 0.00861803f $X=0.82 $Y=1.765 $X2=0 $Y2=0
cc_57 N_D1_c_49_n N_Y_c_229_n 0.0112146f $X=0.82 $Y=1.765 $X2=0 $Y2=0
cc_58 N_D1_c_50_n N_Y_c_229_n 0.00317526f $X=0.835 $Y=1.22 $X2=0 $Y2=0
cc_59 D1 N_Y_c_229_n 0.0186037f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_60 N_D1_c_49_n N_Y_c_232_n 0.0153438f $X=0.82 $Y=1.765 $X2=0 $Y2=0
cc_61 D1 N_Y_c_232_n 0.0221856f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_62 N_D1_c_49_n N_Y_c_230_n 0.00110132f $X=0.82 $Y=1.765 $X2=0 $Y2=0
cc_63 N_D1_c_50_n N_Y_c_230_n 0.0105771f $X=0.835 $Y=1.22 $X2=0 $Y2=0
cc_64 D1 N_Y_c_230_n 0.0150353f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_65 N_D1_c_49_n N_Y_c_236_n 0.00250598f $X=0.82 $Y=1.765 $X2=0 $Y2=0
cc_66 D1 N_Y_c_236_n 0.00234631f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_67 N_D1_c_49_n N_Y_c_237_n 0.0175796f $X=0.82 $Y=1.765 $X2=0 $Y2=0
cc_68 N_D1_c_50_n N_VGND_c_311_n 0.00433162f $X=0.835 $Y=1.22 $X2=0 $Y2=0
cc_69 N_D1_c_50_n N_VGND_c_313_n 0.00822327f $X=0.835 $Y=1.22 $X2=0 $Y2=0
cc_70 N_C1_c_74_n N_B1_c_108_n 0.0274744f $X=1.225 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_71 C1 N_B1_c_108_n 0.00865512f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_72 N_C1_c_75_n N_B1_c_109_n 0.0415974f $X=1.27 $Y=1.765 $X2=0 $Y2=0
cc_73 C1 N_B1_c_109_n 3.45051e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_74 N_C1_c_75_n N_B1_c_110_n 0.00198614f $X=1.27 $Y=1.765 $X2=0 $Y2=0
cc_75 C1 N_B1_c_110_n 0.0299123f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_76 N_C1_c_75_n N_VPWR_c_191_n 0.0105538f $X=1.27 $Y=1.765 $X2=0 $Y2=0
cc_77 N_C1_c_75_n N_VPWR_c_196_n 0.00326636f $X=1.27 $Y=1.765 $X2=0 $Y2=0
cc_78 N_C1_c_75_n N_VPWR_c_189_n 0.0047469f $X=1.27 $Y=1.765 $X2=0 $Y2=0
cc_79 N_C1_c_75_n N_Y_c_234_n 0.00692056f $X=1.27 $Y=1.765 $X2=0 $Y2=0
cc_80 C1 N_Y_c_234_n 0.00850845f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_81 N_C1_c_74_n N_Y_c_230_n 9.85906e-19 $X=1.225 $Y=1.22 $X2=0 $Y2=0
cc_82 C1 N_Y_c_230_n 0.030281f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_83 N_C1_c_75_n N_Y_c_236_n 0.00618089f $X=1.27 $Y=1.765 $X2=0 $Y2=0
cc_84 C1 N_Y_c_236_n 0.0199629f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_85 N_C1_c_75_n N_Y_c_237_n 0.0218603f $X=1.27 $Y=1.765 $X2=0 $Y2=0
cc_86 C1 A_182_74# 0.00751072f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_87 C1 A_260_74# 0.00953457f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_88 C1 N_A_368_74#_c_285_n 0.00723659f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_89 N_C1_c_74_n N_A_368_74#_c_282_n 7.73661e-19 $X=1.225 $Y=1.22 $X2=0 $Y2=0
cc_90 C1 N_A_368_74#_c_282_n 0.0160909f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_91 N_C1_c_74_n N_VGND_c_311_n 0.00303293f $X=1.225 $Y=1.22 $X2=0 $Y2=0
cc_92 C1 N_VGND_c_311_n 0.00877891f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_93 N_C1_c_74_n N_VGND_c_313_n 0.00372419f $X=1.225 $Y=1.22 $X2=0 $Y2=0
cc_94 C1 N_VGND_c_313_n 0.0110375f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_95 N_B1_c_108_n N_A2_c_137_n 0.0193073f $X=1.765 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_96 N_B1_c_109_n N_A2_c_138_n 0.0411695f $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_97 N_B1_c_110_n N_A2_c_138_n 4.15266e-19 $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_98 N_B1_c_109_n A2 4.1351e-19 $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_99 N_B1_c_110_n A2 0.0249496f $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_100 N_B1_c_109_n N_VPWR_c_191_n 0.00363267f $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_101 N_B1_c_109_n N_VPWR_c_197_n 0.00461464f $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_102 N_B1_c_109_n N_VPWR_c_189_n 0.00909489f $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_103 N_B1_c_109_n N_Y_c_234_n 0.0202121f $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_104 N_B1_c_110_n N_Y_c_234_n 0.0295555f $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_105 N_B1_c_109_n N_Y_c_235_n 4.36072e-19 $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_106 N_B1_c_109_n N_Y_c_237_n 4.95897e-19 $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_107 N_B1_c_108_n N_A_368_74#_c_285_n 0.0027133f $X=1.765 $Y=1.22 $X2=0 $Y2=0
cc_108 N_B1_c_109_n N_A_368_74#_c_285_n 8.89733e-19 $X=1.9 $Y=1.765 $X2=0 $Y2=0
cc_109 N_B1_c_110_n N_A_368_74#_c_285_n 0.011699f $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_110 N_B1_c_108_n N_A_368_74#_c_282_n 0.0082564f $X=1.765 $Y=1.22 $X2=0 $Y2=0
cc_111 N_B1_c_108_n N_VGND_c_310_n 5.94017e-19 $X=1.765 $Y=1.22 $X2=0 $Y2=0
cc_112 N_B1_c_108_n N_VGND_c_311_n 0.00445602f $X=1.765 $Y=1.22 $X2=0 $Y2=0
cc_113 N_B1_c_108_n N_VGND_c_313_n 0.00859779f $X=1.765 $Y=1.22 $X2=0 $Y2=0
cc_114 N_A2_c_138_n N_A1_c_166_n 0.0821501f $X=2.375 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_115 A2 N_A1_c_166_n 0.00906015f $X=2.555 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_116 N_A2_c_137_n N_A1_c_167_n 0.0198738f $X=2.275 $Y=1.22 $X2=0 $Y2=0
cc_117 A2 N_A1_c_167_n 3.9318e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_118 N_A2_c_138_n A1 2.10483e-19 $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_119 A2 A1 0.0290366f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_120 N_A2_c_138_n N_VPWR_c_193_n 0.00397156f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A2_c_138_n N_VPWR_c_197_n 0.00445602f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A2_c_138_n N_VPWR_c_189_n 0.00858784f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A2_c_138_n N_Y_c_234_n 0.00786791f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_124 A2 N_Y_c_234_n 0.00963966f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_125 N_A2_c_138_n N_Y_c_235_n 0.0201405f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A2_c_137_n N_A_368_74#_c_282_n 0.00267906f $X=2.275 $Y=1.22 $X2=0 $Y2=0
cc_127 N_A2_c_137_n N_A_368_74#_c_283_n 0.0128517f $X=2.275 $Y=1.22 $X2=0 $Y2=0
cc_128 N_A2_c_138_n N_A_368_74#_c_283_n 0.00101205f $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_129 A2 N_A_368_74#_c_283_n 0.0398068f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A2_c_137_n N_A_368_74#_c_284_n 8.66094e-19 $X=2.275 $Y=1.22 $X2=0 $Y2=0
cc_131 N_A2_c_137_n N_VGND_c_310_n 0.00759f $X=2.275 $Y=1.22 $X2=0 $Y2=0
cc_132 N_A2_c_137_n N_VGND_c_311_n 0.00383152f $X=2.275 $Y=1.22 $X2=0 $Y2=0
cc_133 N_A2_c_137_n N_VGND_c_313_n 0.0038476f $X=2.275 $Y=1.22 $X2=0 $Y2=0
cc_134 N_A1_c_166_n N_VPWR_c_193_n 0.03076f $X=2.83 $Y=1.765 $X2=0 $Y2=0
cc_135 A1 N_VPWR_c_193_n 0.017696f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_136 N_A1_c_166_n N_VPWR_c_197_n 0.00413917f $X=2.83 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A1_c_166_n N_VPWR_c_189_n 0.00817855f $X=2.83 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A1_c_166_n N_Y_c_234_n 6.72262e-19 $X=2.83 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A1_c_166_n N_Y_c_235_n 0.00322942f $X=2.83 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A1_c_166_n N_A_368_74#_c_283_n 0.00199248f $X=2.83 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A1_c_167_n N_A_368_74#_c_283_n 0.013911f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_142 A1 N_A_368_74#_c_283_n 0.0252927f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_143 N_A1_c_167_n N_A_368_74#_c_284_n 0.00854971f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_144 N_A1_c_167_n N_VGND_c_310_n 0.00499784f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_145 N_A1_c_167_n N_VGND_c_312_n 0.00434272f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_146 N_A1_c_167_n N_VGND_c_313_n 0.00449889f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_147 N_VPWR_M1003_s N_Y_c_232_n 0.00346832f $X=0.4 $Y=1.84 $X2=0 $Y2=0
cc_148 N_VPWR_c_190_n N_Y_c_232_n 0.025036f $X=0.545 $Y=2.145 $X2=0 $Y2=0
cc_149 N_VPWR_M1005_d N_Y_c_234_n 0.00644688f $X=1.345 $Y=1.84 $X2=0 $Y2=0
cc_150 N_VPWR_c_191_n N_Y_c_234_n 0.0229431f $X=1.65 $Y=2.145 $X2=0 $Y2=0
cc_151 N_VPWR_c_193_n N_Y_c_234_n 0.00203979f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_152 N_VPWR_c_191_n N_Y_c_235_n 0.00158095f $X=1.65 $Y=2.145 $X2=0 $Y2=0
cc_153 N_VPWR_c_193_n N_Y_c_235_n 0.029941f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_154 N_VPWR_c_197_n N_Y_c_235_n 0.0145938f $X=2.89 $Y=3.33 $X2=0 $Y2=0
cc_155 N_VPWR_c_189_n N_Y_c_235_n 0.0120466f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_156 N_VPWR_c_190_n N_Y_c_237_n 0.0368013f $X=0.545 $Y=2.145 $X2=0 $Y2=0
cc_157 N_VPWR_c_191_n N_Y_c_237_n 0.0729358f $X=1.65 $Y=2.145 $X2=0 $Y2=0
cc_158 N_VPWR_c_196_n N_Y_c_237_n 0.0189233f $X=1.485 $Y=3.33 $X2=0 $Y2=0
cc_159 N_VPWR_c_189_n N_Y_c_237_n 0.0153506f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_160 N_Y_c_230_n N_VGND_c_311_n 0.0296309f $X=0.62 $Y=0.515 $X2=0 $Y2=0
cc_161 N_Y_c_230_n N_VGND_c_313_n 0.024582f $X=0.62 $Y=0.515 $X2=0 $Y2=0
cc_162 N_A_368_74#_c_283_n N_VGND_M1002_d 0.00792129f $X=2.915 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_163 N_A_368_74#_c_282_n N_VGND_c_310_n 0.0105237f $X=1.99 $Y=0.515 $X2=0
+ $Y2=0
cc_164 N_A_368_74#_c_283_n N_VGND_c_310_n 0.0207516f $X=2.915 $Y=0.925 $X2=0
+ $Y2=0
cc_165 N_A_368_74#_c_284_n N_VGND_c_310_n 0.0102004f $X=3.08 $Y=0.515 $X2=0
+ $Y2=0
cc_166 N_A_368_74#_c_282_n N_VGND_c_311_n 0.0145621f $X=1.99 $Y=0.515 $X2=0
+ $Y2=0
cc_167 N_A_368_74#_c_284_n N_VGND_c_312_n 0.0145323f $X=3.08 $Y=0.515 $X2=0
+ $Y2=0
cc_168 N_A_368_74#_c_282_n N_VGND_c_313_n 0.0120343f $X=1.99 $Y=0.515 $X2=0
+ $Y2=0
cc_169 N_A_368_74#_c_283_n N_VGND_c_313_n 0.0115465f $X=2.915 $Y=0.925 $X2=0
+ $Y2=0
cc_170 N_A_368_74#_c_284_n N_VGND_c_313_n 0.0119861f $X=3.08 $Y=0.515 $X2=0
+ $Y2=0
