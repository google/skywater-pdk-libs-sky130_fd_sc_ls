* File: sky130_fd_sc_ls__nor4bb_1.spice
* Created: Wed Sep  2 11:16:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nor4bb_1.pex.spice"
.subckt sky130_fd_sc_ls__nor4bb_1  VNB VPB C_N A B D_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D_N	D_N
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_C_N_M1003_g N_A_27_112#_M1003_s VNB NSHORT L=0.15 W=0.55
+ AD=0.142488 AS=0.3025 PD=1.04457 PS=2.2 NRD=30 NRS=0 M=1 R=3.66667 SA=75000.5
+ SB=75003.8 A=0.0825 P=1.4 MULT=1
MM1009 N_Y_M1009_d N_A_M1009_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.74 AD=0.1295
+ AS=0.191712 PD=1.09 PS=1.40543 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.9
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_B_M1008_g N_Y_M1009_d VNB NSHORT L=0.15 W=0.74
+ AD=0.25715 AS=0.1295 PD=1.435 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.4
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1006_d N_A_27_112#_M1006_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.25715 PD=1.09 PS=1.435 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A_611_244#_M1005_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.74
+ AD=0.38024 AS=0.1295 PD=1.89876 PS=1.09 NRD=18.648 NRS=0 M=1 R=4.93333
+ SA=75002.7 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1002 N_A_611_244#_M1002_d N_D_N_M1002_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.55 AD=0.15675 AS=0.28261 PD=1.67 PS=1.41124 NRD=0 NRS=18 M=1 R=3.66667
+ SA=75004 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1007 N_VPWR_M1007_d N_C_N_M1007_g N_A_27_112#_M1007_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.437721 AS=0.2478 PD=1.82143 PS=2.27 NRD=109.296 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75002.9 A=0.126 P=1.98 MULT=1
MM1000 A_313_368# N_A_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.12 AD=0.1512
+ AS=0.583629 PD=1.39 PS=2.42857 NRD=14.0658 NRS=17.5724 M=1 R=7.46667
+ SA=75001.1 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1010 A_397_368# N_B_M1010_g A_313_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.2884
+ AS=0.1512 PD=1.635 PS=1.39 NRD=35.6176 NRS=14.0658 M=1 R=7.46667 SA=75001.5
+ SB=75001.5 A=0.168 P=2.54 MULT=1
MM1001 A_530_368# N_A_27_112#_M1001_g A_397_368# VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2352 AS=0.2884 PD=1.54 PS=1.635 NRD=27.2451 NRS=35.6176 M=1 R=7.46667
+ SA=75002.2 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1011_d N_A_611_244#_M1011_g A_530_368# VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.2352 PD=2.83 PS=1.54 NRD=1.7533 NRS=27.2451 M=1 R=7.46667
+ SA=75002.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1004 N_A_611_244#_M1004_d N_D_N_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.231 PD=2.27 PS=2.23 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.2 A=0.126 P=1.98 MULT=1
DX12_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ls__nor4bb_1.pxi.spice"
*
.ends
*
*
