* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__and2b_2 A_N B VGND VNB VPB VPWR X
X0 VPWR a_198_48# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VPWR B a_198_48# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_505_74# a_27_74# a_198_48# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 VGND a_198_48# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 a_27_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X5 X a_198_48# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 X a_198_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 VGND B a_505_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 a_27_74# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X9 a_198_48# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends
