* File: sky130_fd_sc_ls__o21a_2.pex.spice
* Created: Wed Sep  2 11:17:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O21A_2%A1 1 3 4 6 8 9 10
c23 10 0 1.25174e-19 $X=0.72 $Y=1.295
c24 1 0 1.4014e-19 $X=0.7 $Y=1.22
r25 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.385 $X2=0.61 $Y2=1.385
r26 10 15 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.61 $Y2=1.365
r27 9 15 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.61 $Y2=1.365
r28 8 14 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.625 $Y=1.385
+ $X2=0.61 $Y2=1.385
r29 4 8 107.404 $w=1.72e-07 $l=3.82492e-07 $layer=POLY_cond $X=0.725 $Y=1.765
+ $X2=0.72 $Y2=1.385
r30 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.725 $Y=1.765
+ $X2=0.725 $Y2=2.34
r31 1 8 47.1543 $w=1.72e-07 $l=1.74714e-07 $layer=POLY_cond $X=0.7 $Y=1.22
+ $X2=0.72 $Y2=1.385
r32 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.7 $Y=1.22 $X2=0.7
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_2%A2 1 3 4 6 7
c27 7 0 1.79042e-19 $X=1.2 $Y=1.295
c28 4 0 1.25174e-19 $X=1.31 $Y=1.22
r29 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.385 $X2=1.22 $Y2=1.385
r30 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.22 $Y=1.295 $X2=1.22
+ $Y2=1.385
r31 4 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.31 $Y=1.22
+ $X2=1.22 $Y2=1.385
r32 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.31 $Y=1.22 $X2=1.31
+ $Y2=0.74
r33 1 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=1.145 $Y=1.765
+ $X2=1.22 $Y2=1.385
r34 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.145 $Y=1.765
+ $X2=1.145 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_2%B1 1 3 4 6 7 11
c36 4 0 3.89014e-20 $X=1.785 $Y=1.22
c37 1 0 9.63186e-20 $X=1.715 $Y=1.765
r38 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.385 $X2=1.79 $Y2=1.385
r39 7 11 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.79 $Y2=1.365
r40 4 10 38.9026 $w=2.7e-07 $l=1.67481e-07 $layer=POLY_cond $X=1.785 $Y=1.22
+ $X2=1.79 $Y2=1.385
r41 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.785 $Y=1.22 $X2=1.785
+ $Y2=0.74
r42 1 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=1.715 $Y=1.765
+ $X2=1.79 $Y2=1.385
r43 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.715 $Y=1.765
+ $X2=1.715 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_2%A_244_368# 1 2 7 9 10 12 13 15 16 17 18 20 23
+ 27 28 31 34 36 37 41
r74 46 47 6.5877 $w=4.39e-07 $l=6e-08 $layer=POLY_cond $X=2.855 $Y=1.492
+ $X2=2.915 $Y2=1.492
r75 42 46 41.1731 $w=4.39e-07 $l=3.75e-07 $layer=POLY_cond $X=2.48 $Y=1.492
+ $X2=2.855 $Y2=1.492
r76 42 44 8.23462 $w=4.39e-07 $l=7.5e-08 $layer=POLY_cond $X=2.48 $Y=1.492
+ $X2=2.405 $Y2=1.492
r77 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.48
+ $Y=1.385 $X2=2.48 $Y2=1.385
r78 38 41 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.21 $Y=1.385
+ $X2=2.48 $Y2=1.385
r79 35 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=1.55
+ $X2=2.21 $Y2=1.385
r80 35 36 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.21 $Y=1.55
+ $X2=2.21 $Y2=1.72
r81 34 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=1.22
+ $X2=2.21 $Y2=1.385
r82 34 37 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.21 $Y=1.22
+ $X2=2.21 $Y2=1.01
r83 29 37 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=2.1 $Y=0.815
+ $X2=2.1 $Y2=1.01
r84 29 31 9.16044 $w=3.88e-07 $l=3.1e-07 $layer=LI1_cond $X=2.1 $Y=0.815 $X2=2.1
+ $Y2=0.505
r85 27 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.125 $Y=1.805
+ $X2=2.21 $Y2=1.72
r86 27 28 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.125 $Y=1.805
+ $X2=1.655 $Y2=1.805
r87 23 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.49 $Y=1.985
+ $X2=1.49 $Y2=2.695
r88 21 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.49 $Y=1.89
+ $X2=1.655 $Y2=1.805
r89 21 23 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.49 $Y=1.89
+ $X2=1.49 $Y2=1.985
r90 18 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.345 $Y=1.22
+ $X2=3.345 $Y2=0.74
r91 17 47 30.5413 $w=4.39e-07 $l=2.31482e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.915 $Y2=1.492
r92 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.27 $Y=1.295
+ $X2=3.345 $Y2=1.22
r93 16 17 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.27 $Y=1.295
+ $X2=2.99 $Y2=1.295
r94 13 47 28.1521 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.915 $Y=1.22
+ $X2=2.915 $Y2=1.492
r95 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.915 $Y=1.22
+ $X2=2.915 $Y2=0.74
r96 10 46 28.1521 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=1.492
r97 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=2.4
r98 7 44 28.1521 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=1.492
r99 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=2.4
r100 2 25 400 $w=1.7e-07 $l=9.80752e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=1.84 $X2=1.49 $Y2=2.695
r101 2 23 400 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=1.84 $X2=1.49 $Y2=1.985
r102 1 31 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=1.86
+ $Y=0.37 $X2=2 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_2%VPWR 1 2 3 12 18 24 27 28 29 35 42 49 50 53
+ 56
r42 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 50 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r46 47 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.13 $Y2=3.33
r47 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.6 $Y2=3.33
r48 46 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 46 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 43 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.13 $Y2=3.33
r52 43 45 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 42 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=3.13 $Y2=3.33
r54 42 45 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r58 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 35 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=2.13 $Y2=3.33
r60 35 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 33 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 29 54 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r64 29 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 27 32 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.335 $Y=3.33
+ $X2=0.24 $Y2=3.33
r66 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.335 $Y=3.33
+ $X2=0.5 $Y2=3.33
r67 26 37 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=0.665 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.665 $Y=3.33
+ $X2=0.5 $Y2=3.33
r69 22 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=3.245
+ $X2=3.13 $Y2=3.33
r70 22 24 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=3.13 $Y=3.245
+ $X2=3.13 $Y2=2.225
r71 18 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.13 $Y=2.145
+ $X2=2.13 $Y2=2.825
r72 16 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=3.245
+ $X2=2.13 $Y2=3.33
r73 16 21 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.13 $Y=3.245
+ $X2=2.13 $Y2=2.825
r74 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.5 $Y=1.985 $X2=0.5
+ $Y2=2.695
r75 10 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.5 $Y=3.245 $X2=0.5
+ $Y2=3.33
r76 10 15 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=0.5 $Y=3.245 $X2=0.5
+ $Y2=2.695
r77 3 24 300 $w=1.7e-07 $l=4.74579e-07 $layer=licon1_PDIFF $count=2 $X=2.93
+ $Y=1.84 $X2=3.13 $Y2=2.225
r78 2 21 400 $w=1.7e-07 $l=1.14242e-06 $layer=licon1_PDIFF $count=1 $X=1.79
+ $Y=1.84 $X2=2.13 $Y2=2.825
r79 2 18 400 $w=1.7e-07 $l=4.68295e-07 $layer=licon1_PDIFF $count=1 $X=1.79
+ $Y=1.84 $X2=2.13 $Y2=2.145
r80 1 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.355
+ $Y=1.84 $X2=0.5 $Y2=2.695
r81 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.355
+ $Y=1.84 $X2=0.5 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_2%X 1 2 9 13 14 15 16 22 33
c30 22 0 9.63186e-20 $X=3.13 $Y=1.72
r31 22 33 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=3.13 $Y=1.72
+ $X2=3.13 $Y2=1.665
r32 16 22 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=3.12 $Y=1.805
+ $X2=3.13 $Y2=1.805
r33 16 33 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.13 $Y=1.65
+ $X2=3.13 $Y2=1.665
r34 15 16 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.13 $Y=1.295
+ $X2=3.13 $Y2=1.65
r35 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.13 $Y=0.925
+ $X2=3.13 $Y2=1.295
r36 13 14 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.13 $Y=0.515
+ $X2=3.13 $Y2=0.925
r37 9 11 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.63 $Y=1.985
+ $X2=2.63 $Y2=2.815
r38 7 16 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.63 $Y=1.805
+ $X2=3.12 $Y2=1.805
r39 7 9 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.63 $Y=1.89 $X2=2.63
+ $Y2=1.985
r40 2 11 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=2.815
r41 2 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=1.985
r42 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.99
+ $Y=0.37 $X2=3.13 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_2%A_54_74# 1 2 7 9 11 13 15
r26 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.84 $X2=1.57
+ $Y2=0.925
r27 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.57 $Y=0.84
+ $X2=1.57 $Y2=0.505
r28 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=0.925
+ $X2=0.415 $Y2=0.925
r29 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=0.925
+ $X2=1.57 $Y2=0.925
r30 11 12 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.405 $Y=0.925
+ $X2=0.58 $Y2=0.925
r31 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.415 $Y=0.84 $X2=0.415
+ $Y2=0.925
r32 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.415 $Y=0.84
+ $X2=0.415 $Y2=0.505
r33 2 20 182 $w=1.7e-07 $l=6.40859e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.37 $X2=1.57 $Y2=0.925
r34 2 15 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.37 $X2=1.57 $Y2=0.505
r35 1 18 182 $w=1.7e-07 $l=6.23298e-07 $layer=licon1_NDIFF $count=1 $X=0.27
+ $Y=0.37 $X2=0.415 $Y2=0.925
r36 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.27
+ $Y=0.37 $X2=0.415 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LS__O21A_2%VGND 1 2 3 12 16 18 20 22 24 29 34 40 43 47
r44 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r45 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 38 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r48 38 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r49 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r50 35 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.63
+ $Y2=0
r51 35 37 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=3.12
+ $Y2=0
r52 34 46 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=3.475 $Y=0 $X2=3.657
+ $Y2=0
r53 34 37 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.475 $Y=0 $X2=3.12
+ $Y2=0
r54 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r55 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r56 30 40 11.0851 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=0.992
+ $Y2=0
r57 30 32 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=2.16
+ $Y2=0
r58 29 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.63
+ $Y2=0
r59 29 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.16
+ $Y2=0
r60 27 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r61 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r62 24 40 11.0851 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=0.75 $Y=0 $X2=0.992
+ $Y2=0
r63 24 26 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=0.75 $Y=0 $X2=0.72
+ $Y2=0
r64 22 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r65 22 41 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r66 18 46 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.6 $Y=0.085
+ $X2=3.657 $Y2=0
r67 18 20 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=3.6 $Y=0.085 $X2=3.6
+ $Y2=0.515
r68 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0
r69 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0.515
r70 10 40 1.99554 $w=4.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.992 $Y=0.085
+ $X2=0.992 $Y2=0
r71 10 12 10.6044 $w=4.83e-07 $l=4.3e-07 $layer=LI1_cond $X=0.992 $Y=0.085
+ $X2=0.992 $Y2=0.515
r72 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.42
+ $Y=0.37 $X2=3.56 $Y2=0.515
r73 2 16 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=2.485
+ $Y=0.37 $X2=2.63 $Y2=0.515
r74 1 12 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=0.775
+ $Y=0.37 $X2=0.99 $Y2=0.515
.ends

