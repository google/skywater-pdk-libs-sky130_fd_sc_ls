* File: sky130_fd_sc_ls__and2_4.spice
* Created: Wed Sep  2 10:54:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__and2_4.pex.spice"
.subckt sky130_fd_sc_ls__and2_4  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_X_M1000_d N_A_83_269#_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1002 N_X_M1000_d N_A_83_269#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1010 N_X_M1010_d N_A_83_269#_M1010_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1591 AS=0.1036 PD=1.17 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1015 N_X_M1010_d N_A_83_269#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1591 AS=0.13883 PD=1.17 PS=1.17971 NRD=12.972 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1003 N_A_504_119#_M1003_d N_B_M1003_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0976 AS=0.12007 PD=0.945 PS=1.02029 NRD=0 NRS=14.988 M=1 R=4.26667
+ SA=75002.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1001 N_A_83_269#_M1001_d N_A_M1001_g N_A_504_119#_M1003_d VNB NSHORT L=0.15
+ W=0.64 AD=0.104 AS=0.0976 PD=0.965 PS=0.945 NRD=8.436 NRS=4.68 M=1 R=4.26667
+ SA=75002.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1006 N_A_83_269#_M1001_d N_A_M1006_g N_A_504_119#_M1006_s VNB NSHORT L=0.15
+ W=0.64 AD=0.104 AS=0.096 PD=0.965 PS=0.94 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.1
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1007 N_A_504_119#_M1006_s N_B_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.64
+ AD=0.096 AS=0.1824 PD=0.94 PS=1.85 NRD=3.744 NRS=0 M=1 R=4.26667 SA=75003.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_A_83_269#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_83_269#_M1011_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1012 N_VPWR_M1011_d N_A_83_269#_M1012_g N_X_M1012_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.1792 PD=1.42 PS=1.44 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1013_d N_A_83_269#_M1013_g N_X_M1012_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.228486 AS=0.1792 PD=1.72 PS=1.44 NRD=1.7533 NRS=5.2599 M=1 R=7.46667
+ SA=75001.6 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1013_d N_B_M1005_g N_A_83_269#_M1005_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.171364 AS=0.1365 PD=1.29 PS=1.165 NRD=22.852 NRS=2.3443 M=1 R=5.6
+ SA=75002.1 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_A_83_269#_M1005_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1365 AS=0.1365 PD=1.165 PS=1.165 NRD=8.1952 NRS=8.1952 M=1 R=5.6
+ SA=75002.6 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1014 N_VPWR_M1004_d N_A_M1014_g N_A_83_269#_M1014_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1365 AS=0.126 PD=1.165 PS=1.14 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75003.1
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_B_M1009_g N_A_83_269#_M1014_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2478 AS=0.126 PD=2.27 PS=1.14 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75003.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.742 P=13.12
c_83 VPB 0 2.91098e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__and2_4.pxi.spice"
*
.ends
*
*
