* File: sky130_fd_sc_ls__o31a_4.spice
* Created: Wed Sep  2 11:22:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o31a_4.pex.spice"
.subckt sky130_fd_sc_ls__o31a_4  VNB VPB B1 A3 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* A3	A3
* B1	B1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_86_260#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_86_260#_M1007_g N_X_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.10915 AS=0.1036 PD=1.035 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1007_d N_A_86_260#_M1016_g N_X_M1016_s VNB NSHORT L=0.15 W=0.74
+ AD=0.10915 AS=0.1036 PD=1.035 PS=1.02 NRD=2.424 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_A_86_260#_M1018_g N_X_M1016_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_492_125#_M1008_d N_B1_M1008_g N_A_86_260#_M1008_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1952 AS=0.1056 PD=1.89 PS=0.97 NRD=3.744 NRS=9.372 M=1 R=4.26667
+ SA=75000.2 SB=75003.6 A=0.096 P=1.58 MULT=1
MM1022 N_A_492_125#_M1022_d N_B1_M1022_g N_A_86_260#_M1008_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1408 AS=0.1056 PD=1.08 PS=0.97 NRD=14.988 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1019 N_VGND_M1019_d N_A3_M1019_g N_A_492_125#_M1022_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1408 PD=0.92 PS=1.08 NRD=0 NRS=14.988 M=1 R=4.26667 SA=75001.3
+ SB=75002.5 A=0.096 P=1.58 MULT=1
MM1021 N_VGND_M1019_d N_A3_M1021_g N_A_492_125#_M1021_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.7
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g N_A_492_125#_M1021_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.2
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1013 N_VGND_M1010_d N_A1_M1013_g N_A_492_125#_M1013_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75002.6
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1017 N_VGND_M1017_d N_A1_M1017_g N_A_492_125#_M1013_s VNB NSHORT L=0.15 W=0.64
+ AD=0.112 AS=0.112 PD=0.99 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.1
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1014 N_VGND_M1017_d N_A2_M1014_g N_A_492_125#_M1014_s VNB NSHORT L=0.15 W=0.64
+ AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75003.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_A_86_260#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1004_d N_A_86_260#_M1004_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75002 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1004_d N_A_86_260#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1015 N_VPWR_M1015_d N_A_86_260#_M1015_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.222098 AS=0.168 PD=1.59019 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1006 N_A_86_260#_M1006_d N_B1_M1006_g N_VPWR_M1015_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.198302 PD=1.3 PS=1.41981 NRD=1.9503 NRS=19.0302 M=1 R=6.66667
+ SA=75002.1 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1012 N_A_86_260#_M1006_d N_B1_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75002.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_A_699_392#_M1001_d N_A3_M1001_g N_A_86_260#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.6 A=0.15 P=2.3 MULT=1
MM1020 N_A_699_392#_M1020_d N_A3_M1020_g N_A_86_260#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1002 N_A_968_392#_M1002_d N_A2_M1002_g N_A_699_392#_M1020_d VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_968_392#_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.15 PD=1.35 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.6
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1005_d N_A1_M1011_g N_A_968_392#_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.17 PD=1.35 PS=1.34 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75002.1 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1023 N_A_968_392#_M1011_s N_A2_M1023_g N_A_699_392#_M1023_s VPB PHIGHVT L=0.15
+ W=1 AD=0.17 AS=0.305 PD=1.34 PS=2.61 NRD=9.8303 NRS=3.9203 M=1 R=6.66667
+ SA=75002.6 SB=75000.2 A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.206 P=17.92
c_73 VNB 0 1.74626e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__o31a_4.pxi.spice"
*
.ends
*
*
