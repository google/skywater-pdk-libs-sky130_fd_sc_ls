* File: sky130_fd_sc_ls__dfbbn_2.pxi.spice
* Created: Wed Sep  2 11:00:30 2020
* 
x_PM_SKY130_FD_SC_LS__DFBBN_2%CLK_N N_CLK_N_M1032_g N_CLK_N_c_293_n
+ N_CLK_N_M1028_g CLK_N N_CLK_N_c_294_n PM_SKY130_FD_SC_LS__DFBBN_2%CLK_N
x_PM_SKY130_FD_SC_LS__DFBBN_2%D N_D_M1015_g N_D_c_324_n N_D_c_328_n N_D_M1039_g
+ D D N_D_c_326_n PM_SKY130_FD_SC_LS__DFBBN_2%D
x_PM_SKY130_FD_SC_LS__DFBBN_2%A_473_405# N_A_473_405#_M1035_d
+ N_A_473_405#_M1040_s N_A_473_405#_M1011_d N_A_473_405#_M1031_g
+ N_A_473_405#_c_374_n N_A_473_405#_M1024_g N_A_473_405#_M1000_g
+ N_A_473_405#_c_375_n N_A_473_405#_M1002_g N_A_473_405#_c_376_n
+ N_A_473_405#_c_377_n N_A_473_405#_c_378_n N_A_473_405#_c_379_n
+ N_A_473_405#_c_368_n N_A_473_405#_c_369_n N_A_473_405#_c_370_n
+ N_A_473_405#_c_444_p N_A_473_405#_c_381_n N_A_473_405#_c_371_n
+ N_A_473_405#_c_372_n N_A_473_405#_c_384_n N_A_473_405#_c_385_n
+ N_A_473_405#_c_386_n PM_SKY130_FD_SC_LS__DFBBN_2%A_473_405#
x_PM_SKY130_FD_SC_LS__DFBBN_2%A_200_74# N_A_200_74#_M1033_d N_A_200_74#_M1029_d
+ N_A_200_74#_c_559_n N_A_200_74#_M1042_g N_A_200_74#_M1023_g
+ N_A_200_74#_c_543_n N_A_200_74#_M1041_g N_A_200_74#_c_544_n
+ N_A_200_74#_M1001_g N_A_200_74#_c_561_n N_A_200_74#_c_545_n
+ N_A_200_74#_c_562_n N_A_200_74#_c_563_n N_A_200_74#_c_564_n
+ N_A_200_74#_c_565_n N_A_200_74#_c_579_n N_A_200_74#_c_566_n
+ N_A_200_74#_c_546_n N_A_200_74#_c_547_n N_A_200_74#_c_548_n
+ N_A_200_74#_c_549_n N_A_200_74#_c_568_n N_A_200_74#_c_550_n
+ N_A_200_74#_c_551_n N_A_200_74#_c_570_n N_A_200_74#_c_552_n
+ N_A_200_74#_c_553_n N_A_200_74#_c_554_n N_A_200_74#_c_583_n
+ N_A_200_74#_c_555_n N_A_200_74#_c_556_n N_A_200_74#_c_557_n
+ N_A_200_74#_c_558_n PM_SKY130_FD_SC_LS__DFBBN_2%A_200_74#
x_PM_SKY130_FD_SC_LS__DFBBN_2%A_601_119# N_A_601_119#_M1037_d
+ N_A_601_119#_M1042_d N_A_601_119#_c_771_n N_A_601_119#_c_778_n
+ N_A_601_119#_c_779_n N_A_601_119#_M1040_g N_A_601_119#_c_772_n
+ N_A_601_119#_M1035_g N_A_601_119#_c_773_n N_A_601_119#_c_794_n
+ N_A_601_119#_c_803_n N_A_601_119#_c_781_n N_A_601_119#_c_774_n
+ N_A_601_119#_c_775_n N_A_601_119#_c_776_n
+ PM_SKY130_FD_SC_LS__DFBBN_2%A_601_119#
x_PM_SKY130_FD_SC_LS__DFBBN_2%A_975_322# N_A_975_322#_M1022_s
+ N_A_975_322#_M1021_s N_A_975_322#_c_878_n N_A_975_322#_M1017_g
+ N_A_975_322#_M1005_g N_A_975_322#_M1019_g N_A_975_322#_c_880_n
+ N_A_975_322#_c_900_n N_A_975_322#_M1036_g N_A_975_322#_c_881_n
+ N_A_975_322#_c_882_n N_A_975_322#_c_883_n N_A_975_322#_c_884_n
+ N_A_975_322#_c_885_n N_A_975_322#_c_886_n N_A_975_322#_c_887_n
+ N_A_975_322#_c_888_n N_A_975_322#_c_889_n N_A_975_322#_c_890_n
+ N_A_975_322#_c_891_n N_A_975_322#_c_892_n N_A_975_322#_c_893_n
+ N_A_975_322#_c_894_n N_A_975_322#_c_902_n N_A_975_322#_c_903_n
+ N_A_975_322#_c_895_n N_A_975_322#_c_982_p N_A_975_322#_c_896_n
+ N_A_975_322#_c_897_n PM_SKY130_FD_SC_LS__DFBBN_2%A_975_322#
x_PM_SKY130_FD_SC_LS__DFBBN_2%SET_B N_SET_B_c_1063_n N_SET_B_M1011_g
+ N_SET_B_M1003_g N_SET_B_c_1065_n N_SET_B_M1030_g N_SET_B_M1009_g
+ N_SET_B_c_1067_n N_SET_B_c_1072_n N_SET_B_c_1073_n SET_B N_SET_B_c_1068_n
+ N_SET_B_c_1076_n PM_SKY130_FD_SC_LS__DFBBN_2%SET_B
x_PM_SKY130_FD_SC_LS__DFBBN_2%A_27_74# N_A_27_74#_M1032_s N_A_27_74#_M1028_s
+ N_A_27_74#_M1033_g N_A_27_74#_c_1192_n N_A_27_74#_M1029_g N_A_27_74#_c_1193_n
+ N_A_27_74#_c_1194_n N_A_27_74#_M1037_g N_A_27_74#_c_1196_n N_A_27_74#_c_1209_n
+ N_A_27_74#_c_1210_n N_A_27_74#_c_1211_n N_A_27_74#_c_1212_n N_A_27_74#_M1043_g
+ N_A_27_74#_M1034_g N_A_27_74#_c_1198_n N_A_27_74#_c_1199_n N_A_27_74#_c_1213_n
+ N_A_27_74#_c_1214_n N_A_27_74#_M1010_g N_A_27_74#_c_1200_n N_A_27_74#_c_1201_n
+ N_A_27_74#_c_1216_n N_A_27_74#_c_1217_n N_A_27_74#_c_1218_n
+ N_A_27_74#_c_1202_n N_A_27_74#_c_1203_n N_A_27_74#_c_1204_n
+ N_A_27_74#_c_1232_n N_A_27_74#_c_1205_n N_A_27_74#_c_1206_n
+ N_A_27_74#_c_1207_n PM_SKY130_FD_SC_LS__DFBBN_2%A_27_74#
x_PM_SKY130_FD_SC_LS__DFBBN_2%A_1555_410# N_A_1555_410#_M1019_d
+ N_A_1555_410#_M1030_s N_A_1555_410#_M1014_d N_A_1555_410#_c_1392_n
+ N_A_1555_410#_M1004_g N_A_1555_410#_c_1393_n N_A_1555_410#_M1018_g
+ N_A_1555_410#_c_1395_n N_A_1555_410#_M1012_g N_A_1555_410#_c_1383_n
+ N_A_1555_410#_M1027_g N_A_1555_410#_c_1396_n N_A_1555_410#_M1020_g
+ N_A_1555_410#_c_1384_n N_A_1555_410#_M1038_g N_A_1555_410#_c_1385_n
+ N_A_1555_410#_c_1386_n N_A_1555_410#_c_1387_n N_A_1555_410#_M1013_g
+ N_A_1555_410#_M1025_g N_A_1555_410#_c_1400_n N_A_1555_410#_c_1401_n
+ N_A_1555_410#_c_1402_n N_A_1555_410#_c_1458_n N_A_1555_410#_c_1403_n
+ N_A_1555_410#_c_1389_n N_A_1555_410#_c_1404_n N_A_1555_410#_c_1405_n
+ N_A_1555_410#_c_1406_n N_A_1555_410#_c_1407_n N_A_1555_410#_c_1408_n
+ N_A_1555_410#_c_1409_n N_A_1555_410#_c_1430_n N_A_1555_410#_c_1390_n
+ N_A_1555_410#_c_1391_n PM_SKY130_FD_SC_LS__DFBBN_2%A_1555_410#
x_PM_SKY130_FD_SC_LS__DFBBN_2%A_1335_112# N_A_1335_112#_M1034_d
+ N_A_1335_112#_M1041_d N_A_1335_112#_M1008_g N_A_1335_112#_c_1606_n
+ N_A_1335_112#_M1014_g N_A_1335_112#_c_1607_n N_A_1335_112#_c_1611_n
+ N_A_1335_112#_c_1612_n N_A_1335_112#_c_1613_n N_A_1335_112#_c_1608_n
+ N_A_1335_112#_c_1615_n N_A_1335_112#_c_1659_n N_A_1335_112#_c_1616_n
+ N_A_1335_112#_c_1609_n N_A_1335_112#_c_1618_n N_A_1335_112#_c_1619_n
+ N_A_1335_112#_c_1620_n N_A_1335_112#_c_1621_n
+ PM_SKY130_FD_SC_LS__DFBBN_2%A_1335_112#
x_PM_SKY130_FD_SC_LS__DFBBN_2%RESET_B N_RESET_B_c_1744_n N_RESET_B_M1021_g
+ N_RESET_B_c_1745_n N_RESET_B_M1022_g RESET_B N_RESET_B_c_1746_n
+ PM_SKY130_FD_SC_LS__DFBBN_2%RESET_B
x_PM_SKY130_FD_SC_LS__DFBBN_2%A_2516_368# N_A_2516_368#_M1025_s
+ N_A_2516_368#_M1013_s N_A_2516_368#_c_1780_n N_A_2516_368#_M1007_g
+ N_A_2516_368#_M1006_g N_A_2516_368#_c_1781_n N_A_2516_368#_M1016_g
+ N_A_2516_368#_M1026_g N_A_2516_368#_c_1782_n N_A_2516_368#_c_1783_n
+ N_A_2516_368#_c_1776_n N_A_2516_368#_c_1777_n N_A_2516_368#_c_1784_n
+ N_A_2516_368#_c_1778_n N_A_2516_368#_c_1779_n
+ PM_SKY130_FD_SC_LS__DFBBN_2%A_2516_368#
x_PM_SKY130_FD_SC_LS__DFBBN_2%VPWR N_VPWR_M1028_d N_VPWR_M1039_d N_VPWR_M1017_d
+ N_VPWR_M1002_s N_VPWR_M1004_d N_VPWR_M1030_d N_VPWR_M1021_d N_VPWR_M1020_s
+ N_VPWR_M1013_d N_VPWR_M1016_s N_VPWR_c_1854_n N_VPWR_c_1855_n N_VPWR_c_1856_n
+ N_VPWR_c_1857_n N_VPWR_c_1858_n N_VPWR_c_1859_n N_VPWR_c_1860_n
+ N_VPWR_c_1861_n N_VPWR_c_1862_n N_VPWR_c_1863_n N_VPWR_c_1864_n
+ N_VPWR_c_1865_n N_VPWR_c_1866_n N_VPWR_c_1867_n N_VPWR_c_1868_n
+ N_VPWR_c_1869_n N_VPWR_c_1870_n VPWR N_VPWR_c_1871_n N_VPWR_c_1872_n
+ N_VPWR_c_1873_n N_VPWR_c_1874_n N_VPWR_c_1875_n N_VPWR_c_1876_n
+ N_VPWR_c_1877_n N_VPWR_c_1878_n N_VPWR_c_1879_n N_VPWR_c_1880_n
+ N_VPWR_c_1881_n N_VPWR_c_1853_n PM_SKY130_FD_SC_LS__DFBBN_2%VPWR
x_PM_SKY130_FD_SC_LS__DFBBN_2%A_311_119# N_A_311_119#_M1015_s
+ N_A_311_119#_M1023_d N_A_311_119#_M1039_s N_A_311_119#_M1043_d
+ N_A_311_119#_c_2026_n N_A_311_119#_c_2045_n N_A_311_119#_c_2027_n
+ N_A_311_119#_c_2028_n N_A_311_119#_c_2029_n N_A_311_119#_c_2030_n
+ N_A_311_119#_c_2037_n N_A_311_119#_c_2038_n N_A_311_119#_c_2039_n
+ N_A_311_119#_c_2031_n N_A_311_119#_c_2032_n N_A_311_119#_c_2033_n
+ N_A_311_119#_c_2034_n N_A_311_119#_c_2035_n
+ PM_SKY130_FD_SC_LS__DFBBN_2%A_311_119#
x_PM_SKY130_FD_SC_LS__DFBBN_2%Q_N N_Q_N_M1027_s N_Q_N_M1012_d N_Q_N_c_2157_n
+ N_Q_N_c_2155_n N_Q_N_c_2171_n Q_N Q_N Q_N PM_SKY130_FD_SC_LS__DFBBN_2%Q_N
x_PM_SKY130_FD_SC_LS__DFBBN_2%Q N_Q_M1006_d N_Q_M1007_d N_Q_c_2193_n
+ N_Q_c_2194_n N_Q_c_2196_n N_Q_c_2198_n Q Q Q PM_SKY130_FD_SC_LS__DFBBN_2%Q
x_PM_SKY130_FD_SC_LS__DFBBN_2%VGND N_VGND_M1032_d N_VGND_M1015_d N_VGND_M1003_d
+ N_VGND_M1018_d N_VGND_M1022_d N_VGND_M1038_d N_VGND_M1025_d N_VGND_M1026_s
+ N_VGND_c_2229_n N_VGND_c_2230_n N_VGND_c_2231_n N_VGND_c_2232_n
+ N_VGND_c_2233_n N_VGND_c_2234_n N_VGND_c_2235_n N_VGND_c_2236_n VGND
+ N_VGND_c_2237_n N_VGND_c_2238_n N_VGND_c_2239_n N_VGND_c_2240_n
+ N_VGND_c_2241_n N_VGND_c_2242_n N_VGND_c_2243_n N_VGND_c_2244_n
+ N_VGND_c_2245_n N_VGND_c_2246_n N_VGND_c_2247_n N_VGND_c_2248_n
+ N_VGND_c_2249_n N_VGND_c_2250_n N_VGND_c_2251_n N_VGND_c_2252_n
+ PM_SKY130_FD_SC_LS__DFBBN_2%VGND
x_PM_SKY130_FD_SC_LS__DFBBN_2%A_867_125# N_A_867_125#_M1035_s
+ N_A_867_125#_M1005_d N_A_867_125#_c_2376_n N_A_867_125#_c_2377_n
+ N_A_867_125#_c_2378_n N_A_867_125#_c_2379_n
+ PM_SKY130_FD_SC_LS__DFBBN_2%A_867_125#
x_PM_SKY130_FD_SC_LS__DFBBN_2%A_1832_74# N_A_1832_74#_M1009_d
+ N_A_1832_74#_M1008_d N_A_1832_74#_c_2416_n N_A_1832_74#_c_2410_n
+ N_A_1832_74#_c_2411_n N_A_1832_74#_c_2412_n
+ PM_SKY130_FD_SC_LS__DFBBN_2%A_1832_74#
cc_1 VNB N_CLK_N_M1032_g 0.0292041f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_CLK_N_c_293_n 0.0461135f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_3 VNB N_CLK_N_c_294_n 0.016346f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_4 VNB N_D_M1015_g 0.0218268f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_5 VNB N_D_c_324_n 0.00965277f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_6 VNB D 0.00754307f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_7 VNB N_D_c_326_n 0.04446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_473_405#_M1031_g 0.0389929f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_9 VNB N_A_473_405#_M1000_g 0.0363908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_473_405#_c_368_n 0.00254694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_473_405#_c_369_n 0.00356345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_473_405#_c_370_n 0.00167311f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_473_405#_c_371_n 0.00142582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_473_405#_c_372_n 0.014186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_200_74#_c_543_n 0.00999107f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.465
cc_16 VNB N_A_200_74#_c_544_n 0.021122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_200_74#_c_545_n 0.0114485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_200_74#_c_546_n 0.00467856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_200_74#_c_547_n 0.00205587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_200_74#_c_548_n 0.00377088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_200_74#_c_549_n 0.0107632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_200_74#_c_550_n 0.0100185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_200_74#_c_551_n 0.00932659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_200_74#_c_552_n 0.00439927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_200_74#_c_553_n 0.0476318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_200_74#_c_554_n 0.0406152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_200_74#_c_555_n 0.0020871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_200_74#_c_556_n 0.034084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_200_74#_c_557_n 0.00495044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_200_74#_c_558_n 0.0162715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_601_119#_c_771_n 0.0284123f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_32 VNB N_A_601_119#_c_772_n 0.0141357f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_33 VNB N_A_601_119#_c_773_n 0.0368475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_601_119#_c_774_n 0.0080484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_601_119#_c_775_n 0.00105081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_601_119#_c_776_n 0.00758961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_975_322#_c_878_n 0.00886992f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_38 VNB N_A_975_322#_M1005_g 0.0322965f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_39 VNB N_A_975_322#_c_880_n 0.00627748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_975_322#_c_881_n 0.00170742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_975_322#_c_882_n 0.018117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_975_322#_c_883_n 5.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_975_322#_c_884_n 0.00348971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_975_322#_c_885_n 0.049584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_975_322#_c_886_n 0.00300857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_975_322#_c_887_n 0.00289067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_975_322#_c_888_n 0.0144768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_975_322#_c_889_n 8.92125e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_975_322#_c_890_n 0.00663725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_975_322#_c_891_n 0.0318897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_975_322#_c_892_n 0.00993441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_975_322#_c_893_n 0.0107497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_975_322#_c_894_n 0.00688916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_975_322#_c_895_n 4.96706e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_975_322#_c_896_n 0.00214173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_975_322#_c_897_n 0.0156811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_SET_B_c_1063_n 0.0072424f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_58 VNB N_SET_B_M1003_g 0.0336951f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_59 VNB N_SET_B_c_1065_n 0.0173889f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_60 VNB N_SET_B_M1009_g 0.0302798f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.465
cc_61 VNB N_SET_B_c_1067_n 0.00458063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_SET_B_c_1068_n 0.0014129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_27_74#_M1033_g 0.0195304f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.465
cc_64 VNB N_A_27_74#_c_1192_n 0.0366902f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_65 VNB N_A_27_74#_c_1193_n 0.134018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_27_74#_c_1194_n 0.0113774f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.665
cc_67 VNB N_A_27_74#_M1037_g 0.0477822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_27_74#_c_1196_n 0.263846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_27_74#_M1034_g 0.0299979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_27_74#_c_1198_n 0.0503085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_27_74#_c_1199_n 0.00907112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_27_74#_c_1200_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_27_74#_c_1201_n 0.0188481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_27_74#_c_1202_n 0.0247745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_27_74#_c_1203_n 0.00333636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_27_74#_c_1204_n 0.00916851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_27_74#_c_1205_n 0.0033318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_27_74#_c_1206_n 7.84349e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_27_74#_c_1207_n 0.00267302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1555_410#_M1018_g 0.0422621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1555_410#_c_1383_n 0.0171089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1555_410#_c_1384_n 0.0172736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1555_410#_c_1385_n 0.0480337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1555_410#_c_1386_n 0.0357841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1555_410#_c_1387_n 0.0138262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1555_410#_M1025_g 0.03301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1555_410#_c_1389_n 0.0128564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1555_410#_c_1390_n 0.00358533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1555_410#_c_1391_n 0.00185235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1335_112#_M1008_g 0.0335173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1335_112#_c_1606_n 0.0189776f $X=-0.19 $Y=-0.245 $X2=0.33
+ $Y2=1.465
cc_92 VNB N_A_1335_112#_c_1607_n 0.0105465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1335_112#_c_1608_n 0.0074943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1335_112#_c_1609_n 0.00337646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_RESET_B_c_1744_n 0.0285916f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_96 VNB N_RESET_B_c_1745_n 0.0193585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_RESET_B_c_1746_n 0.00461828f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_98 VNB N_A_2516_368#_M1006_g 0.0205325f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_99 VNB N_A_2516_368#_M1026_g 0.0227577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2516_368#_c_1776_n 0.0138925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_2516_368#_c_1777_n 0.0109236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_2516_368#_c_1778_n 0.00101278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_2516_368#_c_1779_n 0.055377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VPWR_c_1853_n 0.601534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_311_119#_c_2026_n 0.0125638f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=1.665
cc_106 VNB N_A_311_119#_c_2027_n 0.00190227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_311_119#_c_2028_n 0.00165852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_311_119#_c_2029_n 0.0091336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_311_119#_c_2030_n 0.00381631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_311_119#_c_2031_n 0.00817927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_311_119#_c_2032_n 0.0025518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_311_119#_c_2033_n 0.00200249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_311_119#_c_2034_n 0.0115642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_311_119#_c_2035_n 0.00951758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_Q_N_c_2155_n 8.47293e-19 $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_116 VNB Q_N 0.00279061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_Q_c_2193_n 0.00214054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_Q_c_2194_n 0.0188601f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_119 VNB N_VGND_c_2229_n 0.00222691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2230_n 0.00955289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2231_n 0.00678165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2232_n 0.01013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2233_n 0.0262467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2234_n 0.00938091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2235_n 0.0115487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2236_n 0.0226839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2237_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2238_n 0.0307998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2239_n 0.0768126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2240_n 0.0662733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2241_n 0.0200226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2242_n 0.019905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2243_n 0.0168561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2244_n 0.00501873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2245_n 0.00526018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2246_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2247_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2248_n 0.040772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2249_n 0.0315104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2250_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2251_n 0.00528956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2252_n 0.717897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_A_867_125#_c_2376_n 0.00598735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_A_867_125#_c_2377_n 0.0198023f $X=-0.19 $Y=-0.245 $X2=0.33
+ $Y2=1.465
cc_145 VNB N_A_867_125#_c_2378_n 0.00343796f $X=-0.19 $Y=-0.245 $X2=0.33
+ $Y2=1.465
cc_146 VNB N_A_867_125#_c_2379_n 0.00475019f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=1.665
cc_147 VNB N_A_1832_74#_c_2410_n 0.00162646f $X=-0.19 $Y=-0.245 $X2=0.33
+ $Y2=1.465
cc_148 VNB N_A_1832_74#_c_2411_n 0.00542253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_A_1832_74#_c_2412_n 0.0030118f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=1.665
cc_150 VPB N_CLK_N_c_293_n 0.0289622f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_151 VPB N_CLK_N_c_294_n 0.00727431f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_152 VPB N_D_c_324_n 0.0391307f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_153 VPB N_D_c_328_n 0.0227778f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_154 VPB N_A_473_405#_M1031_g 0.020268f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_155 VPB N_A_473_405#_c_374_n 0.0492991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_473_405#_c_375_n 0.0177302f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_473_405#_c_376_n 0.00180276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_473_405#_c_377_n 0.0220831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_473_405#_c_378_n 0.00131809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_473_405#_c_379_n 0.00502838f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_473_405#_c_368_n 0.0031906f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_473_405#_c_381_n 0.00789632f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_473_405#_c_371_n 0.00618103f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_473_405#_c_372_n 0.0444742f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_473_405#_c_384_n 0.00562746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_473_405#_c_385_n 0.00195558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_473_405#_c_386_n 0.00831545f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_200_74#_c_559_n 0.0506207f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_169 VPB N_A_200_74#_c_543_n 0.0452928f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.465
cc_170 VPB N_A_200_74#_c_561_n 0.011188f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_200_74#_c_562_n 0.0118289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_200_74#_c_563_n 0.00442365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_200_74#_c_564_n 0.00581697f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_200_74#_c_565_n 0.0203135f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_200_74#_c_566_n 0.00414584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_200_74#_c_548_n 0.00124778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_200_74#_c_568_n 0.00970887f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_200_74#_c_550_n 0.0030323f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_200_74#_c_570_n 2.5096e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_601_119#_c_771_n 0.00394935f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_181 VPB N_A_601_119#_c_778_n 0.00805961f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_182 VPB N_A_601_119#_c_779_n 0.0227156f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_601_119#_c_773_n 0.0286451f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_601_119#_c_781_n 0.00551783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_601_119#_c_776_n 0.00746621f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_975_322#_c_878_n 0.0443399f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_187 VPB N_A_975_322#_c_880_n 0.00773999f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_975_322#_c_900_n 0.023562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_975_322#_c_893_n 0.00634404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_975_322#_c_902_n 0.00425184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_975_322#_c_903_n 0.00393056f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_975_322#_c_895_n 0.0021807f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_SET_B_c_1063_n 0.0500271f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_194 VPB N_SET_B_c_1065_n 0.0375544f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_195 VPB N_SET_B_c_1067_n 0.00237939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_SET_B_c_1072_n 0.0354504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_SET_B_c_1073_n 0.00274556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB SET_B 0.00143942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_SET_B_c_1068_n 0.00165254f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_SET_B_c_1076_n 0.00115456f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_27_74#_c_1192_n 0.0258938f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_202 VPB N_A_27_74#_c_1209_n 0.0359501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_27_74#_c_1210_n 0.00648852f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_27_74#_c_1211_n 0.0326387f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_27_74#_c_1212_n 0.0220289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_27_74#_c_1213_n 0.0238245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_27_74#_c_1214_n 0.0221135f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_27_74#_c_1201_n 0.00752409f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_27_74#_c_1216_n 0.0116114f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_27_74#_c_1217_n 0.00805193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_27_74#_c_1218_n 0.0357063f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_27_74#_c_1206_n 0.00278492f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1555_410#_c_1392_n 0.0171656f $X=-0.19 $Y=1.66 $X2=0.375
+ $Y2=1.465
cc_214 VPB N_A_1555_410#_c_1393_n 0.0107571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_1555_410#_M1018_g 0.0040972f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1555_410#_c_1395_n 0.0168357f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1555_410#_c_1396_n 0.0174986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_1555_410#_c_1385_n 0.0281536f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_1555_410#_c_1386_n 0.0246364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_1555_410#_c_1387_n 0.0256466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_1555_410#_c_1400_n 0.0216656f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_1555_410#_c_1401_n 0.00185087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1555_410#_c_1402_n 0.0667315f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1555_410#_c_1403_n 0.0168669f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1555_410#_c_1404_n 0.00116731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1555_410#_c_1405_n 0.00302121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1555_410#_c_1406_n 0.0116305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1555_410#_c_1407_n 0.00122019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_1555_410#_c_1408_n 0.00620857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_1555_410#_c_1409_n 0.00590798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_1555_410#_c_1390_n 0.00195054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_1335_112#_c_1606_n 0.0402764f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_233 VPB N_A_1335_112#_c_1611_n 0.00336771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_1335_112#_c_1612_n 0.011416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_1335_112#_c_1613_n 0.00138366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_1335_112#_c_1608_n 0.00168665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_1335_112#_c_1615_n 0.00507963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_1335_112#_c_1616_n 0.00362369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_1335_112#_c_1609_n 0.00901319f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_1335_112#_c_1618_n 0.00122055f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_1335_112#_c_1619_n 0.00271803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_1335_112#_c_1620_n 0.00241115f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_1335_112#_c_1621_n 0.00853468f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_RESET_B_c_1744_n 0.0303249f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_245 VPB N_RESET_B_c_1746_n 0.00416237f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_246 VPB N_A_2516_368#_c_1780_n 0.0160425f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_247 VPB N_A_2516_368#_c_1781_n 0.0164199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_2516_368#_c_1782_n 0.00303355f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_2516_368#_c_1783_n 0.0123996f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_2516_368#_c_1784_n 0.00176f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_2516_368#_c_1779_n 0.0148059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1854_n 0.00770537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1855_n 0.00830666f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1856_n 0.00658128f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1857_n 0.010011f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1858_n 0.0223371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1859_n 0.0172425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1860_n 0.016172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1861_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1862_n 0.0450285f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1863_n 0.0366957f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1864_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1865_n 0.0635348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1866_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1867_n 0.0199677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1868_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1869_n 0.0143811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1870_n 0.0459699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1871_n 0.0197879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1872_n 0.0196646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1873_n 0.0477054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1874_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1875_n 0.0208242f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1876_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1877_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1878_n 0.0139421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1879_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1880_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1881_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1853_n 0.191421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_311_119#_c_2026_n 0.0148481f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.665
cc_282 VPB N_A_311_119#_c_2037_n 0.0102982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_311_119#_c_2038_n 0.0123143f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_A_311_119#_c_2039_n 0.00419923f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_311_119#_c_2032_n 0.00341626f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_Q_N_c_2157_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_Q_N_c_2155_n 0.00127472f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_288 VPB N_Q_c_2194_n 0.00393307f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_289 VPB N_Q_c_2196_n 0.00501111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB Q 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_291 N_CLK_N_c_293_n N_A_200_74#_c_561_n 6.23412e-19 $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_292 N_CLK_N_c_293_n N_A_27_74#_c_1192_n 0.0473578f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_293 N_CLK_N_c_294_n N_A_27_74#_c_1192_n 2.76539e-19 $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_294 N_CLK_N_M1032_g N_A_27_74#_c_1194_n 0.0271107f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_295 N_CLK_N_c_293_n N_A_27_74#_c_1217_n 0.0016558f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_296 N_CLK_N_c_294_n N_A_27_74#_c_1217_n 0.0249655f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_297 N_CLK_N_c_293_n N_A_27_74#_c_1218_n 0.0104891f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_298 N_CLK_N_M1032_g N_A_27_74#_c_1202_n 0.00159319f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_299 N_CLK_N_M1032_g N_A_27_74#_c_1203_n 0.0145993f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_300 N_CLK_N_c_293_n N_A_27_74#_c_1203_n 9.73098e-19 $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_301 N_CLK_N_c_294_n N_A_27_74#_c_1203_n 0.00971403f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_302 N_CLK_N_c_293_n N_A_27_74#_c_1204_n 0.00158295f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_303 N_CLK_N_c_294_n N_A_27_74#_c_1204_n 0.0209549f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_304 N_CLK_N_c_293_n N_A_27_74#_c_1232_n 0.0139266f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_305 N_CLK_N_c_294_n N_A_27_74#_c_1232_n 0.00433199f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_306 N_CLK_N_M1032_g N_A_27_74#_c_1205_n 0.00383463f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_307 N_CLK_N_c_293_n N_A_27_74#_c_1206_n 0.00487653f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_308 N_CLK_N_c_294_n N_A_27_74#_c_1206_n 0.0113335f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_309 N_CLK_N_c_293_n N_A_27_74#_c_1207_n 0.00235667f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_310 N_CLK_N_c_294_n N_A_27_74#_c_1207_n 0.0269075f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_311 N_CLK_N_c_293_n N_VPWR_c_1854_n 0.00486623f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_312 N_CLK_N_c_293_n N_VPWR_c_1871_n 0.00445602f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_313 N_CLK_N_c_293_n N_VPWR_c_1853_n 0.00861134f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_314 N_CLK_N_M1032_g N_VGND_c_2229_n 0.0125189f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_315 N_CLK_N_M1032_g N_VGND_c_2237_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_316 N_CLK_N_M1032_g N_VGND_c_2252_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_317 N_D_M1015_g N_A_473_405#_M1031_g 0.0145675f $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_318 N_D_c_324_n N_A_473_405#_M1031_g 0.0158704f $X=2.01 $Y=2.35 $X2=0 $Y2=0
cc_319 D N_A_473_405#_M1031_g 0.0133258f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_320 N_D_c_326_n N_A_473_405#_M1031_g 0.0213733f $X=2.12 $Y=1.345 $X2=0 $Y2=0
cc_321 N_D_c_324_n N_A_473_405#_c_374_n 0.015988f $X=2.01 $Y=2.35 $X2=0 $Y2=0
cc_322 N_D_c_328_n N_A_473_405#_c_374_n 0.011617f $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_323 N_D_c_328_n N_A_473_405#_c_376_n 2.4885e-19 $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_324 N_D_c_324_n N_A_473_405#_c_384_n 4.05702e-19 $X=2.01 $Y=2.35 $X2=0 $Y2=0
cc_325 N_D_c_328_n N_A_200_74#_c_561_n 0.00318693f $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_326 N_D_M1015_g N_A_200_74#_c_545_n 0.00293016f $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_327 N_D_c_328_n N_A_200_74#_c_562_n 0.0102018f $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_328 N_D_c_324_n N_A_200_74#_c_564_n 0.0117083f $X=2.01 $Y=2.35 $X2=0 $Y2=0
cc_329 N_D_c_328_n N_A_200_74#_c_564_n 0.0157085f $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_330 D N_A_200_74#_c_565_n 0.0470514f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_331 N_D_c_326_n N_A_200_74#_c_565_n 0.00357357f $X=2.12 $Y=1.345 $X2=0 $Y2=0
cc_332 N_D_c_324_n N_A_200_74#_c_579_n 0.00803832f $X=2.01 $Y=2.35 $X2=0 $Y2=0
cc_333 D N_A_200_74#_c_579_n 0.0133696f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_334 N_D_c_326_n N_A_200_74#_c_579_n 5.80967e-19 $X=2.12 $Y=1.345 $X2=0 $Y2=0
cc_335 D N_A_200_74#_c_546_n 0.00354331f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_336 D N_A_200_74#_c_583_n 0.00643738f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_337 D N_A_200_74#_c_557_n 0.0135499f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_338 N_D_c_326_n N_A_27_74#_c_1192_n 0.00191984f $X=2.12 $Y=1.345 $X2=0 $Y2=0
cc_339 N_D_M1015_g N_A_27_74#_c_1193_n 0.00999521f $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_340 D N_A_27_74#_M1037_g 0.00262641f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_341 N_D_c_328_n N_VPWR_c_1855_n 0.00177169f $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_342 N_D_c_328_n N_VPWR_c_1863_n 9.62598e-19 $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_343 N_D_M1015_g N_A_311_119#_c_2026_n 0.0127716f $X=1.915 $Y=0.805 $X2=0
+ $Y2=0
cc_344 N_D_c_324_n N_A_311_119#_c_2026_n 0.021905f $X=2.01 $Y=2.35 $X2=0 $Y2=0
cc_345 N_D_c_328_n N_A_311_119#_c_2026_n 0.00575009f $X=2.01 $Y=2.44 $X2=0 $Y2=0
cc_346 D N_A_311_119#_c_2026_n 0.0262091f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_347 N_D_M1015_g N_A_311_119#_c_2045_n 0.0110649f $X=1.915 $Y=0.805 $X2=0
+ $Y2=0
cc_348 D N_A_311_119#_c_2045_n 0.0544193f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_349 N_D_c_326_n N_A_311_119#_c_2045_n 0.0069224f $X=2.12 $Y=1.345 $X2=0 $Y2=0
cc_350 N_D_M1015_g N_A_311_119#_c_2027_n 7.90383e-19 $X=1.915 $Y=0.805 $X2=0
+ $Y2=0
cc_351 N_D_M1015_g N_A_311_119#_c_2033_n 0.00775522f $X=1.915 $Y=0.805 $X2=0
+ $Y2=0
cc_352 N_D_M1015_g N_VGND_c_2230_n 0.00256919f $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_353 N_D_M1015_g N_VGND_c_2252_n 9.39239e-19 $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_354 N_A_473_405#_c_374_n N_A_200_74#_c_559_n 0.0519381f $X=2.605 $Y=2.44
+ $X2=0 $Y2=0
cc_355 N_A_473_405#_c_376_n N_A_200_74#_c_559_n 0.00695333f $X=2.72 $Y=2.905
+ $X2=0 $Y2=0
cc_356 N_A_473_405#_c_377_n N_A_200_74#_c_559_n 0.0125924f $X=4.185 $Y=2.99
+ $X2=0 $Y2=0
cc_357 N_A_473_405#_c_384_n N_A_200_74#_c_559_n 0.00219513f $X=2.72 $Y=2.19
+ $X2=0 $Y2=0
cc_358 N_A_473_405#_M1000_g N_A_200_74#_c_543_n 0.00111182f $X=6.125 $Y=0.9
+ $X2=0 $Y2=0
cc_359 N_A_473_405#_c_375_n N_A_200_74#_c_543_n 0.0464592f $X=6.485 $Y=2.045
+ $X2=0 $Y2=0
cc_360 N_A_473_405#_c_371_n N_A_200_74#_c_543_n 9.50289e-19 $X=6.215 $Y=1.795
+ $X2=0 $Y2=0
cc_361 N_A_473_405#_c_372_n N_A_200_74#_c_543_n 0.026425f $X=6.215 $Y=1.795
+ $X2=0 $Y2=0
cc_362 N_A_473_405#_M1031_g N_A_200_74#_c_564_n 0.00289829f $X=2.57 $Y=0.805
+ $X2=0 $Y2=0
cc_363 N_A_473_405#_c_374_n N_A_200_74#_c_564_n 0.00224895f $X=2.605 $Y=2.44
+ $X2=0 $Y2=0
cc_364 N_A_473_405#_c_376_n N_A_200_74#_c_564_n 0.00512793f $X=2.72 $Y=2.905
+ $X2=0 $Y2=0
cc_365 N_A_473_405#_c_384_n N_A_200_74#_c_564_n 0.0195339f $X=2.72 $Y=2.19 $X2=0
+ $Y2=0
cc_366 N_A_473_405#_M1031_g N_A_200_74#_c_565_n 0.0111042f $X=2.57 $Y=0.805
+ $X2=0 $Y2=0
cc_367 N_A_473_405#_c_374_n N_A_200_74#_c_565_n 0.00418988f $X=2.605 $Y=2.44
+ $X2=0 $Y2=0
cc_368 N_A_473_405#_c_384_n N_A_200_74#_c_565_n 0.0329615f $X=2.72 $Y=2.19 $X2=0
+ $Y2=0
cc_369 N_A_473_405#_M1031_g N_A_200_74#_c_566_n 0.00512098f $X=2.57 $Y=0.805
+ $X2=0 $Y2=0
cc_370 N_A_473_405#_c_374_n N_A_200_74#_c_566_n 2.96042e-19 $X=2.605 $Y=2.44
+ $X2=0 $Y2=0
cc_371 N_A_473_405#_c_377_n N_A_200_74#_c_566_n 0.00315571f $X=4.185 $Y=2.99
+ $X2=0 $Y2=0
cc_372 N_A_473_405#_c_384_n N_A_200_74#_c_566_n 0.0262106f $X=2.72 $Y=2.19 $X2=0
+ $Y2=0
cc_373 N_A_473_405#_M1031_g N_A_200_74#_c_546_n 0.00173341f $X=2.57 $Y=0.805
+ $X2=0 $Y2=0
cc_374 N_A_473_405#_M1000_g N_A_200_74#_c_547_n 4.59312e-19 $X=6.125 $Y=0.9
+ $X2=0 $Y2=0
cc_375 N_A_473_405#_M1000_g N_A_200_74#_c_548_n 0.00337066f $X=6.125 $Y=0.9
+ $X2=0 $Y2=0
cc_376 N_A_473_405#_c_371_n N_A_200_74#_c_548_n 0.010434f $X=6.215 $Y=1.795
+ $X2=0 $Y2=0
cc_377 N_A_473_405#_c_372_n N_A_200_74#_c_548_n 0.00120462f $X=6.215 $Y=1.795
+ $X2=0 $Y2=0
cc_378 N_A_473_405#_M1000_g N_A_200_74#_c_554_n 0.00635926f $X=6.125 $Y=0.9
+ $X2=0 $Y2=0
cc_379 N_A_473_405#_c_368_n N_A_200_74#_c_554_n 0.0119957f $X=4.69 $Y=2.305
+ $X2=0 $Y2=0
cc_380 N_A_473_405#_c_369_n N_A_200_74#_c_554_n 0.0294005f $X=4.905 $Y=0.95
+ $X2=0 $Y2=0
cc_381 N_A_473_405#_c_371_n N_A_200_74#_c_554_n 0.00209182f $X=6.215 $Y=1.795
+ $X2=0 $Y2=0
cc_382 N_A_473_405#_c_372_n N_A_200_74#_c_554_n 0.00354269f $X=6.215 $Y=1.795
+ $X2=0 $Y2=0
cc_383 N_A_473_405#_M1031_g N_A_200_74#_c_557_n 6.41937e-19 $X=2.57 $Y=0.805
+ $X2=0 $Y2=0
cc_384 N_A_473_405#_c_377_n N_A_601_119#_M1042_d 0.00250812f $X=4.185 $Y=2.99
+ $X2=0 $Y2=0
cc_385 N_A_473_405#_c_368_n N_A_601_119#_c_771_n 0.0149084f $X=4.69 $Y=2.305
+ $X2=0 $Y2=0
cc_386 N_A_473_405#_c_369_n N_A_601_119#_c_771_n 0.00142228f $X=4.905 $Y=0.95
+ $X2=0 $Y2=0
cc_387 N_A_473_405#_c_368_n N_A_601_119#_c_778_n 0.00293098f $X=4.69 $Y=2.305
+ $X2=0 $Y2=0
cc_388 N_A_473_405#_c_377_n N_A_601_119#_c_779_n 0.00690373f $X=4.185 $Y=2.99
+ $X2=0 $Y2=0
cc_389 N_A_473_405#_c_379_n N_A_601_119#_c_779_n 0.0100662f $X=4.395 $Y=2.905
+ $X2=0 $Y2=0
cc_390 N_A_473_405#_c_368_n N_A_601_119#_c_779_n 0.00866773f $X=4.69 $Y=2.305
+ $X2=0 $Y2=0
cc_391 N_A_473_405#_c_385_n N_A_601_119#_c_779_n 0.0112004f $X=4.35 $Y=2.39
+ $X2=0 $Y2=0
cc_392 N_A_473_405#_c_369_n N_A_601_119#_c_772_n 0.0143026f $X=4.905 $Y=0.95
+ $X2=0 $Y2=0
cc_393 N_A_473_405#_c_370_n N_A_601_119#_c_772_n 0.00485412f $X=4.91 $Y=0.86
+ $X2=0 $Y2=0
cc_394 N_A_473_405#_c_385_n N_A_601_119#_c_773_n 0.00164109f $X=4.35 $Y=2.39
+ $X2=0 $Y2=0
cc_395 N_A_473_405#_c_376_n N_A_601_119#_c_794_n 0.00873904f $X=2.72 $Y=2.905
+ $X2=0 $Y2=0
cc_396 N_A_473_405#_c_377_n N_A_601_119#_c_794_n 0.0253034f $X=4.185 $Y=2.99
+ $X2=0 $Y2=0
cc_397 N_A_473_405#_c_376_n N_A_601_119#_c_781_n 0.00639528f $X=2.72 $Y=2.905
+ $X2=0 $Y2=0
cc_398 N_A_473_405#_M1031_g N_A_601_119#_c_775_n 2.98275e-19 $X=2.57 $Y=0.805
+ $X2=0 $Y2=0
cc_399 N_A_473_405#_c_377_n N_A_975_322#_c_878_n 5.64795e-19 $X=4.185 $Y=2.99
+ $X2=0 $Y2=0
cc_400 N_A_473_405#_c_379_n N_A_975_322#_c_878_n 0.00178304f $X=4.395 $Y=2.905
+ $X2=0 $Y2=0
cc_401 N_A_473_405#_c_368_n N_A_975_322#_c_878_n 0.00752208f $X=4.69 $Y=2.305
+ $X2=0 $Y2=0
cc_402 N_A_473_405#_c_369_n N_A_975_322#_c_878_n 0.00421385f $X=4.905 $Y=0.95
+ $X2=0 $Y2=0
cc_403 N_A_473_405#_c_444_p N_A_975_322#_c_878_n 0.0163009f $X=5.565 $Y=2.405
+ $X2=0 $Y2=0
cc_404 N_A_473_405#_c_385_n N_A_975_322#_c_878_n 4.07331e-19 $X=4.35 $Y=2.39
+ $X2=0 $Y2=0
cc_405 N_A_473_405#_c_386_n N_A_975_322#_c_878_n 6.96418e-19 $X=5.73 $Y=2.405
+ $X2=0 $Y2=0
cc_406 N_A_473_405#_c_368_n N_A_975_322#_M1005_g 0.00188131f $X=4.69 $Y=2.305
+ $X2=0 $Y2=0
cc_407 N_A_473_405#_c_369_n N_A_975_322#_M1005_g 0.00763463f $X=4.905 $Y=0.95
+ $X2=0 $Y2=0
cc_408 N_A_473_405#_c_370_n N_A_975_322#_M1005_g 0.00439649f $X=4.91 $Y=0.86
+ $X2=0 $Y2=0
cc_409 N_A_473_405#_c_368_n N_A_975_322#_c_881_n 0.00699031f $X=4.69 $Y=2.305
+ $X2=0 $Y2=0
cc_410 N_A_473_405#_M1000_g N_A_975_322#_c_882_n 0.0127894f $X=6.125 $Y=0.9
+ $X2=0 $Y2=0
cc_411 N_A_473_405#_c_371_n N_A_975_322#_c_882_n 0.0239276f $X=6.215 $Y=1.795
+ $X2=0 $Y2=0
cc_412 N_A_473_405#_c_372_n N_A_975_322#_c_882_n 0.00301153f $X=6.215 $Y=1.795
+ $X2=0 $Y2=0
cc_413 N_A_473_405#_c_368_n N_A_975_322#_c_883_n 0.00754708f $X=4.69 $Y=2.305
+ $X2=0 $Y2=0
cc_414 N_A_473_405#_c_369_n N_A_975_322#_c_883_n 3.48023e-19 $X=4.905 $Y=0.95
+ $X2=0 $Y2=0
cc_415 N_A_473_405#_M1000_g N_A_975_322#_c_884_n 0.00615644f $X=6.125 $Y=0.9
+ $X2=0 $Y2=0
cc_416 N_A_473_405#_c_368_n N_A_975_322#_c_895_n 0.024558f $X=4.69 $Y=2.305
+ $X2=0 $Y2=0
cc_417 N_A_473_405#_c_369_n N_A_975_322#_c_895_n 0.0015534f $X=4.905 $Y=0.95
+ $X2=0 $Y2=0
cc_418 N_A_473_405#_c_444_p N_A_975_322#_c_895_n 0.0106544f $X=5.565 $Y=2.405
+ $X2=0 $Y2=0
cc_419 N_A_473_405#_c_444_p N_SET_B_c_1063_n 0.00936169f $X=5.565 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_420 N_A_473_405#_c_381_n N_SET_B_c_1063_n 0.00108043f $X=6.215 $Y=2.32
+ $X2=-0.19 $Y2=-0.245
cc_421 N_A_473_405#_c_371_n N_SET_B_c_1063_n 0.005367f $X=6.215 $Y=1.795
+ $X2=-0.19 $Y2=-0.245
cc_422 N_A_473_405#_c_372_n N_SET_B_c_1063_n 0.0131884f $X=6.215 $Y=1.795
+ $X2=-0.19 $Y2=-0.245
cc_423 N_A_473_405#_c_386_n N_SET_B_c_1063_n 0.00728739f $X=5.73 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_424 N_A_473_405#_M1000_g N_SET_B_M1003_g 0.0315389f $X=6.125 $Y=0.9 $X2=0
+ $Y2=0
cc_425 N_A_473_405#_c_369_n N_SET_B_M1003_g 3.79105e-19 $X=4.905 $Y=0.95 $X2=0
+ $Y2=0
cc_426 N_A_473_405#_c_375_n N_SET_B_c_1072_n 0.00731159f $X=6.485 $Y=2.045 $X2=0
+ $Y2=0
cc_427 N_A_473_405#_c_381_n N_SET_B_c_1072_n 0.0152534f $X=6.215 $Y=2.32 $X2=0
+ $Y2=0
cc_428 N_A_473_405#_c_371_n N_SET_B_c_1072_n 0.0218749f $X=6.215 $Y=1.795 $X2=0
+ $Y2=0
cc_429 N_A_473_405#_c_372_n N_SET_B_c_1072_n 0.00799711f $X=6.215 $Y=1.795 $X2=0
+ $Y2=0
cc_430 N_A_473_405#_M1011_d N_SET_B_c_1073_n 2.31732e-19 $X=5.58 $Y=2.12 $X2=0
+ $Y2=0
cc_431 N_A_473_405#_c_368_n N_SET_B_c_1073_n 0.00505032f $X=4.69 $Y=2.305 $X2=0
+ $Y2=0
cc_432 N_A_473_405#_c_444_p N_SET_B_c_1073_n 0.00373413f $X=5.565 $Y=2.405 $X2=0
+ $Y2=0
cc_433 N_A_473_405#_c_371_n N_SET_B_c_1073_n 5.57939e-19 $X=6.215 $Y=1.795 $X2=0
+ $Y2=0
cc_434 N_A_473_405#_M1011_d N_SET_B_c_1068_n 0.00139233f $X=5.58 $Y=2.12 $X2=0
+ $Y2=0
cc_435 N_A_473_405#_c_368_n N_SET_B_c_1068_n 0.00289955f $X=4.69 $Y=2.305 $X2=0
+ $Y2=0
cc_436 N_A_473_405#_c_444_p N_SET_B_c_1068_n 0.0179641f $X=5.565 $Y=2.405 $X2=0
+ $Y2=0
cc_437 N_A_473_405#_c_371_n N_SET_B_c_1068_n 0.0232504f $X=6.215 $Y=1.795 $X2=0
+ $Y2=0
cc_438 N_A_473_405#_c_372_n N_SET_B_c_1068_n 0.00143947f $X=6.215 $Y=1.795 $X2=0
+ $Y2=0
cc_439 N_A_473_405#_M1031_g N_A_27_74#_c_1193_n 0.00997995f $X=2.57 $Y=0.805
+ $X2=0 $Y2=0
cc_440 N_A_473_405#_M1031_g N_A_27_74#_M1037_g 0.0821317f $X=2.57 $Y=0.805 $X2=0
+ $Y2=0
cc_441 N_A_473_405#_M1000_g N_A_27_74#_c_1196_n 0.00894529f $X=6.125 $Y=0.9
+ $X2=0 $Y2=0
cc_442 N_A_473_405#_c_377_n N_A_27_74#_c_1212_n 0.0136872f $X=4.185 $Y=2.99
+ $X2=0 $Y2=0
cc_443 N_A_473_405#_c_379_n N_A_27_74#_c_1212_n 0.00461053f $X=4.395 $Y=2.905
+ $X2=0 $Y2=0
cc_444 N_A_473_405#_M1000_g N_A_27_74#_M1034_g 0.0255423f $X=6.125 $Y=0.9 $X2=0
+ $Y2=0
cc_445 N_A_473_405#_c_372_n N_A_27_74#_c_1199_n 0.00259785f $X=6.215 $Y=1.795
+ $X2=0 $Y2=0
cc_446 N_A_473_405#_c_375_n N_A_1335_112#_c_1619_n 0.0028817f $X=6.485 $Y=2.045
+ $X2=0 $Y2=0
cc_447 N_A_473_405#_c_371_n N_A_1335_112#_c_1619_n 0.00340601f $X=6.215 $Y=1.795
+ $X2=0 $Y2=0
cc_448 N_A_473_405#_c_444_p N_VPWR_M1017_d 0.00908618f $X=5.565 $Y=2.405 $X2=0
+ $Y2=0
cc_449 N_A_473_405#_c_381_n N_VPWR_M1002_s 0.00489622f $X=6.215 $Y=2.32 $X2=0
+ $Y2=0
cc_450 N_A_473_405#_c_371_n N_VPWR_M1002_s 0.00288115f $X=6.215 $Y=1.795 $X2=0
+ $Y2=0
cc_451 N_A_473_405#_c_374_n N_VPWR_c_1855_n 0.00469074f $X=2.605 $Y=2.44 $X2=0
+ $Y2=0
cc_452 N_A_473_405#_c_376_n N_VPWR_c_1855_n 0.0266436f $X=2.72 $Y=2.905 $X2=0
+ $Y2=0
cc_453 N_A_473_405#_c_378_n N_VPWR_c_1855_n 0.0135904f $X=2.805 $Y=2.99 $X2=0
+ $Y2=0
cc_454 N_A_473_405#_c_384_n N_VPWR_c_1855_n 0.00817548f $X=2.72 $Y=2.19 $X2=0
+ $Y2=0
cc_455 N_A_473_405#_c_377_n N_VPWR_c_1856_n 0.00614778f $X=4.185 $Y=2.99 $X2=0
+ $Y2=0
cc_456 N_A_473_405#_c_379_n N_VPWR_c_1856_n 0.0084925f $X=4.395 $Y=2.905 $X2=0
+ $Y2=0
cc_457 N_A_473_405#_c_444_p N_VPWR_c_1856_n 0.0205767f $X=5.565 $Y=2.405 $X2=0
+ $Y2=0
cc_458 N_A_473_405#_c_386_n N_VPWR_c_1856_n 0.0122284f $X=5.73 $Y=2.405 $X2=0
+ $Y2=0
cc_459 N_A_473_405#_c_375_n N_VPWR_c_1857_n 0.0106074f $X=6.485 $Y=2.045 $X2=0
+ $Y2=0
cc_460 N_A_473_405#_c_381_n N_VPWR_c_1857_n 0.0198925f $X=6.215 $Y=2.32 $X2=0
+ $Y2=0
cc_461 N_A_473_405#_c_386_n N_VPWR_c_1857_n 0.023773f $X=5.73 $Y=2.405 $X2=0
+ $Y2=0
cc_462 N_A_473_405#_c_374_n N_VPWR_c_1865_n 0.00420085f $X=2.605 $Y=2.44 $X2=0
+ $Y2=0
cc_463 N_A_473_405#_c_377_n N_VPWR_c_1865_n 0.118578f $X=4.185 $Y=2.99 $X2=0
+ $Y2=0
cc_464 N_A_473_405#_c_378_n N_VPWR_c_1865_n 0.0122392f $X=2.805 $Y=2.99 $X2=0
+ $Y2=0
cc_465 N_A_473_405#_c_386_n N_VPWR_c_1867_n 0.0142535f $X=5.73 $Y=2.405 $X2=0
+ $Y2=0
cc_466 N_A_473_405#_c_375_n N_VPWR_c_1870_n 0.00413917f $X=6.485 $Y=2.045 $X2=0
+ $Y2=0
cc_467 N_A_473_405#_c_374_n N_VPWR_c_1853_n 0.00376497f $X=2.605 $Y=2.44 $X2=0
+ $Y2=0
cc_468 N_A_473_405#_c_375_n N_VPWR_c_1853_n 0.00817532f $X=6.485 $Y=2.045 $X2=0
+ $Y2=0
cc_469 N_A_473_405#_c_377_n N_VPWR_c_1853_n 0.0677251f $X=4.185 $Y=2.99 $X2=0
+ $Y2=0
cc_470 N_A_473_405#_c_378_n N_VPWR_c_1853_n 0.00661913f $X=2.805 $Y=2.99 $X2=0
+ $Y2=0
cc_471 N_A_473_405#_c_444_p N_VPWR_c_1853_n 0.0220533f $X=5.565 $Y=2.405 $X2=0
+ $Y2=0
cc_472 N_A_473_405#_c_381_n N_VPWR_c_1853_n 9.09039e-19 $X=6.215 $Y=2.32 $X2=0
+ $Y2=0
cc_473 N_A_473_405#_c_385_n N_VPWR_c_1853_n 0.00631965f $X=4.35 $Y=2.39 $X2=0
+ $Y2=0
cc_474 N_A_473_405#_c_386_n N_VPWR_c_1853_n 0.0119151f $X=5.73 $Y=2.405 $X2=0
+ $Y2=0
cc_475 N_A_473_405#_c_377_n N_A_311_119#_M1043_d 0.00530205f $X=4.185 $Y=2.99
+ $X2=0 $Y2=0
cc_476 N_A_473_405#_M1031_g N_A_311_119#_c_2045_n 0.00943189f $X=2.57 $Y=0.805
+ $X2=0 $Y2=0
cc_477 N_A_473_405#_M1031_g N_A_311_119#_c_2027_n 0.00811923f $X=2.57 $Y=0.805
+ $X2=0 $Y2=0
cc_478 N_A_473_405#_c_377_n N_A_311_119#_c_2037_n 0.0189889f $X=4.185 $Y=2.99
+ $X2=0 $Y2=0
cc_479 N_A_473_405#_c_379_n N_A_311_119#_c_2037_n 0.0184494f $X=4.395 $Y=2.905
+ $X2=0 $Y2=0
cc_480 N_A_473_405#_c_368_n N_A_311_119#_c_2037_n 0.00472472f $X=4.69 $Y=2.305
+ $X2=0 $Y2=0
cc_481 N_A_473_405#_c_385_n N_A_311_119#_c_2037_n 0.0145503f $X=4.35 $Y=2.39
+ $X2=0 $Y2=0
cc_482 N_A_473_405#_M1040_s N_A_311_119#_c_2038_n 0.00258597f $X=4.22 $Y=2.12
+ $X2=0 $Y2=0
cc_483 N_A_473_405#_c_368_n N_A_311_119#_c_2038_n 0.0136799f $X=4.69 $Y=2.305
+ $X2=0 $Y2=0
cc_484 N_A_473_405#_c_385_n N_A_311_119#_c_2038_n 0.0219082f $X=4.35 $Y=2.39
+ $X2=0 $Y2=0
cc_485 N_A_473_405#_c_369_n N_A_311_119#_c_2031_n 0.0056021f $X=4.905 $Y=0.95
+ $X2=0 $Y2=0
cc_486 N_A_473_405#_c_368_n N_A_311_119#_c_2032_n 0.0462789f $X=4.69 $Y=2.305
+ $X2=0 $Y2=0
cc_487 N_A_473_405#_M1031_g N_A_311_119#_c_2033_n 8.39015e-19 $X=2.57 $Y=0.805
+ $X2=0 $Y2=0
cc_488 N_A_473_405#_c_369_n N_A_311_119#_c_2035_n 0.0110901f $X=4.905 $Y=0.95
+ $X2=0 $Y2=0
cc_489 N_A_473_405#_c_376_n A_536_503# 0.00433065f $X=2.72 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_490 N_A_473_405#_c_377_n A_536_503# 0.00331953f $X=4.185 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_491 N_A_473_405#_c_368_n A_930_424# 0.00217075f $X=4.69 $Y=2.305 $X2=-0.19
+ $Y2=-0.245
cc_492 N_A_473_405#_c_444_p A_930_424# 0.00506866f $X=5.565 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_493 N_A_473_405#_c_385_n A_930_424# 0.00179016f $X=4.35 $Y=2.39 $X2=-0.19
+ $Y2=-0.245
cc_494 N_A_473_405#_M1031_g N_VGND_c_2230_n 0.0018517f $X=2.57 $Y=0.805 $X2=0
+ $Y2=0
cc_495 N_A_473_405#_M1000_g N_VGND_c_2231_n 0.00809789f $X=6.125 $Y=0.9 $X2=0
+ $Y2=0
cc_496 N_A_473_405#_M1031_g N_VGND_c_2252_n 7.22543e-19 $X=2.57 $Y=0.805 $X2=0
+ $Y2=0
cc_497 N_A_473_405#_M1000_g N_VGND_c_2252_n 7.97988e-19 $X=6.125 $Y=0.9 $X2=0
+ $Y2=0
cc_498 N_A_473_405#_c_370_n N_A_867_125#_c_2376_n 0.0136817f $X=4.91 $Y=0.86
+ $X2=0 $Y2=0
cc_499 N_A_473_405#_c_370_n N_A_867_125#_c_2377_n 0.026256f $X=4.91 $Y=0.86
+ $X2=0 $Y2=0
cc_500 N_A_473_405#_M1000_g N_A_867_125#_c_2379_n 2.03891e-19 $X=6.125 $Y=0.9
+ $X2=0 $Y2=0
cc_501 N_A_473_405#_c_370_n N_A_867_125#_c_2379_n 0.0137573f $X=4.91 $Y=0.86
+ $X2=0 $Y2=0
cc_502 N_A_200_74#_c_554_n N_A_601_119#_c_771_n 0.00634081f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_503 N_A_200_74#_c_546_n N_A_601_119#_c_773_n 8.68299e-19 $X=3.117 $Y=1.685
+ $X2=0 $Y2=0
cc_504 N_A_200_74#_c_554_n N_A_601_119#_c_773_n 0.00643501f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_505 N_A_200_74#_c_559_n N_A_601_119#_c_794_n 0.00328982f $X=3.025 $Y=2.44
+ $X2=0 $Y2=0
cc_506 N_A_200_74#_c_566_n N_A_601_119#_c_794_n 0.00776399f $X=3.07 $Y=2.19
+ $X2=0 $Y2=0
cc_507 N_A_200_74#_c_554_n N_A_601_119#_c_803_n 0.00614621f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_508 N_A_200_74#_c_556_n N_A_601_119#_c_803_n 0.00234121f $X=3.38 $Y=1.29
+ $X2=0 $Y2=0
cc_509 N_A_200_74#_c_557_n N_A_601_119#_c_803_n 0.0140588f $X=3.38 $Y=1.29 $X2=0
+ $Y2=0
cc_510 N_A_200_74#_c_558_n N_A_601_119#_c_803_n 0.00984914f $X=3.38 $Y=1.125
+ $X2=0 $Y2=0
cc_511 N_A_200_74#_c_559_n N_A_601_119#_c_781_n 0.00336111f $X=3.025 $Y=2.44
+ $X2=0 $Y2=0
cc_512 N_A_200_74#_c_566_n N_A_601_119#_c_781_n 0.0374872f $X=3.07 $Y=2.19 $X2=0
+ $Y2=0
cc_513 N_A_200_74#_c_570_n N_A_601_119#_c_781_n 0.00486729f $X=3.102 $Y=1.77
+ $X2=0 $Y2=0
cc_514 N_A_200_74#_c_546_n N_A_601_119#_c_774_n 3.54416e-19 $X=3.117 $Y=1.685
+ $X2=0 $Y2=0
cc_515 N_A_200_74#_c_554_n N_A_601_119#_c_774_n 0.0133834f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_516 N_A_200_74#_c_583_n N_A_601_119#_c_774_n 3.70253e-19 $X=3.265 $Y=1.295
+ $X2=0 $Y2=0
cc_517 N_A_200_74#_c_556_n N_A_601_119#_c_774_n 0.00224713f $X=3.38 $Y=1.29
+ $X2=0 $Y2=0
cc_518 N_A_200_74#_c_557_n N_A_601_119#_c_774_n 0.0240518f $X=3.38 $Y=1.29 $X2=0
+ $Y2=0
cc_519 N_A_200_74#_c_558_n N_A_601_119#_c_774_n 0.00514335f $X=3.38 $Y=1.125
+ $X2=0 $Y2=0
cc_520 N_A_200_74#_c_554_n N_A_601_119#_c_775_n 2.62589e-19 $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_521 N_A_200_74#_c_583_n N_A_601_119#_c_775_n 0.00277796f $X=3.265 $Y=1.295
+ $X2=0 $Y2=0
cc_522 N_A_200_74#_c_556_n N_A_601_119#_c_775_n 0.00145122f $X=3.38 $Y=1.29
+ $X2=0 $Y2=0
cc_523 N_A_200_74#_c_557_n N_A_601_119#_c_775_n 0.0187249f $X=3.38 $Y=1.29 $X2=0
+ $Y2=0
cc_524 N_A_200_74#_c_558_n N_A_601_119#_c_775_n 0.0090522f $X=3.38 $Y=1.125
+ $X2=0 $Y2=0
cc_525 N_A_200_74#_c_546_n N_A_601_119#_c_776_n 0.0113226f $X=3.117 $Y=1.685
+ $X2=0 $Y2=0
cc_526 N_A_200_74#_c_570_n N_A_601_119#_c_776_n 0.00932708f $X=3.102 $Y=1.77
+ $X2=0 $Y2=0
cc_527 N_A_200_74#_c_554_n N_A_601_119#_c_776_n 0.0152385f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_528 N_A_200_74#_c_556_n N_A_601_119#_c_776_n 9.10257e-19 $X=3.38 $Y=1.29
+ $X2=0 $Y2=0
cc_529 N_A_200_74#_c_557_n N_A_601_119#_c_776_n 0.0111996f $X=3.38 $Y=1.29 $X2=0
+ $Y2=0
cc_530 N_A_200_74#_c_554_n N_A_975_322#_c_878_n 0.00452129f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_531 N_A_200_74#_c_554_n N_A_975_322#_M1005_g 0.00695811f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_532 N_A_200_74#_c_547_n N_A_975_322#_c_882_n 0.00439286f $X=6.95 $Y=1.41
+ $X2=0 $Y2=0
cc_533 N_A_200_74#_c_548_n N_A_975_322#_c_882_n 0.00255362f $X=6.95 $Y=1.745
+ $X2=0 $Y2=0
cc_534 N_A_200_74#_c_554_n N_A_975_322#_c_882_n 0.050214f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_535 N_A_200_74#_c_555_n N_A_975_322#_c_882_n 3.46995e-19 $X=6.96 $Y=1.295
+ $X2=0 $Y2=0
cc_536 N_A_200_74#_c_554_n N_A_975_322#_c_883_n 0.00737607f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_537 N_A_200_74#_c_547_n N_A_975_322#_c_884_n 0.00355597f $X=6.95 $Y=1.41
+ $X2=0 $Y2=0
cc_538 N_A_200_74#_c_554_n N_A_975_322#_c_884_n 0.0135266f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_539 N_A_200_74#_c_555_n N_A_975_322#_c_884_n 2.91867e-19 $X=6.96 $Y=1.295
+ $X2=0 $Y2=0
cc_540 N_A_200_74#_c_544_n N_A_975_322#_c_885_n 0.00455188f $X=8.125 $Y=1.22
+ $X2=0 $Y2=0
cc_541 N_A_200_74#_c_544_n N_A_975_322#_c_887_n 0.00114059f $X=8.125 $Y=1.22
+ $X2=0 $Y2=0
cc_542 N_A_200_74#_c_554_n N_A_975_322#_c_895_n 0.0041092f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_543 N_A_200_74#_c_554_n N_SET_B_M1003_g 0.00638662f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_544 N_A_200_74#_c_543_n N_SET_B_c_1072_n 0.00945489f $X=6.905 $Y=2.045 $X2=0
+ $Y2=0
cc_545 N_A_200_74#_c_548_n N_SET_B_c_1072_n 0.00963642f $X=6.95 $Y=1.745 $X2=0
+ $Y2=0
cc_546 N_A_200_74#_c_549_n N_SET_B_c_1072_n 0.00691152f $X=7.685 $Y=1.295 $X2=0
+ $Y2=0
cc_547 N_A_200_74#_c_555_n N_SET_B_c_1072_n 0.0121439f $X=6.96 $Y=1.295 $X2=0
+ $Y2=0
cc_548 N_A_200_74#_c_554_n N_SET_B_c_1073_n 0.0112743f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_549 N_A_200_74#_c_554_n N_SET_B_c_1068_n 0.00143342f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_550 N_A_200_74#_c_545_n N_A_27_74#_M1033_g 0.00206322f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_551 N_A_200_74#_c_550_n N_A_27_74#_M1033_g 0.00229974f $X=1.225 $Y=1.82 $X2=0
+ $Y2=0
cc_552 N_A_200_74#_c_561_n N_A_27_74#_c_1192_n 0.0110388f $X=1.17 $Y=2.815 $X2=0
+ $Y2=0
cc_553 N_A_200_74#_c_563_n N_A_27_74#_c_1192_n 0.00456398f $X=1.445 $Y=2.99
+ $X2=0 $Y2=0
cc_554 N_A_200_74#_c_568_n N_A_27_74#_c_1192_n 0.0056203f $X=1.17 $Y=1.985 $X2=0
+ $Y2=0
cc_555 N_A_200_74#_c_550_n N_A_27_74#_c_1192_n 0.00804745f $X=1.225 $Y=1.82
+ $X2=0 $Y2=0
cc_556 N_A_200_74#_c_551_n N_A_27_74#_c_1192_n 0.00203031f $X=1.25 $Y=1.13 $X2=0
+ $Y2=0
cc_557 N_A_200_74#_c_545_n N_A_27_74#_c_1193_n 0.00837633f $X=1.14 $Y=0.515
+ $X2=0 $Y2=0
cc_558 N_A_200_74#_c_546_n N_A_27_74#_M1037_g 0.00416694f $X=3.117 $Y=1.685
+ $X2=0 $Y2=0
cc_559 N_A_200_74#_c_583_n N_A_27_74#_M1037_g 0.00283946f $X=3.265 $Y=1.295
+ $X2=0 $Y2=0
cc_560 N_A_200_74#_c_556_n N_A_27_74#_M1037_g 0.021337f $X=3.38 $Y=1.29 $X2=0
+ $Y2=0
cc_561 N_A_200_74#_c_557_n N_A_27_74#_M1037_g 0.00397504f $X=3.38 $Y=1.29 $X2=0
+ $Y2=0
cc_562 N_A_200_74#_c_558_n N_A_27_74#_M1037_g 0.0131066f $X=3.38 $Y=1.125 $X2=0
+ $Y2=0
cc_563 N_A_200_74#_c_558_n N_A_27_74#_c_1196_n 0.00882199f $X=3.38 $Y=1.125
+ $X2=0 $Y2=0
cc_564 N_A_200_74#_c_546_n N_A_27_74#_c_1209_n 0.00494396f $X=3.117 $Y=1.685
+ $X2=0 $Y2=0
cc_565 N_A_200_74#_c_570_n N_A_27_74#_c_1209_n 0.00657744f $X=3.102 $Y=1.77
+ $X2=0 $Y2=0
cc_566 N_A_200_74#_c_556_n N_A_27_74#_c_1209_n 0.0215947f $X=3.38 $Y=1.29 $X2=0
+ $Y2=0
cc_567 N_A_200_74#_c_557_n N_A_27_74#_c_1209_n 0.00223168f $X=3.38 $Y=1.29 $X2=0
+ $Y2=0
cc_568 N_A_200_74#_c_559_n N_A_27_74#_c_1210_n 0.0213562f $X=3.025 $Y=2.44 $X2=0
+ $Y2=0
cc_569 N_A_200_74#_c_565_n N_A_27_74#_c_1210_n 0.00879974f $X=2.975 $Y=1.77
+ $X2=0 $Y2=0
cc_570 N_A_200_74#_c_570_n N_A_27_74#_c_1210_n 0.00123436f $X=3.102 $Y=1.77
+ $X2=0 $Y2=0
cc_571 N_A_200_74#_c_559_n N_A_27_74#_c_1211_n 0.0205153f $X=3.025 $Y=2.44 $X2=0
+ $Y2=0
cc_572 N_A_200_74#_c_566_n N_A_27_74#_c_1211_n 0.00147896f $X=3.07 $Y=2.19 $X2=0
+ $Y2=0
cc_573 N_A_200_74#_c_570_n N_A_27_74#_c_1211_n 2.79334e-19 $X=3.102 $Y=1.77
+ $X2=0 $Y2=0
cc_574 N_A_200_74#_c_559_n N_A_27_74#_c_1212_n 0.0124214f $X=3.025 $Y=2.44 $X2=0
+ $Y2=0
cc_575 N_A_200_74#_c_543_n N_A_27_74#_c_1198_n 0.0176671f $X=6.905 $Y=2.045
+ $X2=0 $Y2=0
cc_576 N_A_200_74#_c_544_n N_A_27_74#_c_1198_n 4.59884e-19 $X=8.125 $Y=1.22
+ $X2=0 $Y2=0
cc_577 N_A_200_74#_c_547_n N_A_27_74#_c_1198_n 0.0145524f $X=6.95 $Y=1.41 $X2=0
+ $Y2=0
cc_578 N_A_200_74#_c_549_n N_A_27_74#_c_1198_n 0.0147998f $X=7.685 $Y=1.295
+ $X2=0 $Y2=0
cc_579 N_A_200_74#_c_553_n N_A_27_74#_c_1198_n 0.0209136f $X=7.85 $Y=1.385 $X2=0
+ $Y2=0
cc_580 N_A_200_74#_c_554_n N_A_27_74#_c_1198_n 0.00183941f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_581 N_A_200_74#_c_554_n N_A_27_74#_c_1199_n 0.00777034f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_582 N_A_200_74#_c_543_n N_A_27_74#_c_1213_n 0.0113011f $X=6.905 $Y=2.045
+ $X2=0 $Y2=0
cc_583 N_A_200_74#_c_543_n N_A_27_74#_c_1214_n 0.0140197f $X=6.905 $Y=2.045
+ $X2=0 $Y2=0
cc_584 N_A_200_74#_c_543_n N_A_27_74#_c_1201_n 0.0207914f $X=6.905 $Y=2.045
+ $X2=0 $Y2=0
cc_585 N_A_200_74#_c_548_n N_A_27_74#_c_1201_n 0.00543189f $X=6.95 $Y=1.745
+ $X2=0 $Y2=0
cc_586 N_A_200_74#_c_549_n N_A_27_74#_c_1201_n 0.00618964f $X=7.685 $Y=1.295
+ $X2=0 $Y2=0
cc_587 N_A_200_74#_c_552_n N_A_27_74#_c_1201_n 5.52136e-19 $X=7.81 $Y=1.295
+ $X2=0 $Y2=0
cc_588 N_A_200_74#_c_543_n N_A_27_74#_c_1216_n 0.00101556f $X=6.905 $Y=2.045
+ $X2=0 $Y2=0
cc_589 N_A_200_74#_c_549_n N_A_27_74#_c_1216_n 3.32419e-19 $X=7.685 $Y=1.295
+ $X2=0 $Y2=0
cc_590 N_A_200_74#_c_561_n N_A_27_74#_c_1218_n 0.00480111f $X=1.17 $Y=2.815
+ $X2=0 $Y2=0
cc_591 N_A_200_74#_c_551_n N_A_27_74#_c_1203_n 0.00142346f $X=1.25 $Y=1.13 $X2=0
+ $Y2=0
cc_592 N_A_200_74#_c_550_n N_A_27_74#_c_1205_n 0.00465906f $X=1.225 $Y=1.82
+ $X2=0 $Y2=0
cc_593 N_A_200_74#_c_568_n N_A_27_74#_c_1206_n 0.00581222f $X=1.17 $Y=1.985
+ $X2=0 $Y2=0
cc_594 N_A_200_74#_c_550_n N_A_27_74#_c_1206_n 0.00543374f $X=1.225 $Y=1.82
+ $X2=0 $Y2=0
cc_595 N_A_200_74#_c_568_n N_A_27_74#_c_1207_n 0.00761489f $X=1.17 $Y=1.985
+ $X2=0 $Y2=0
cc_596 N_A_200_74#_c_550_n N_A_27_74#_c_1207_n 0.0253261f $X=1.225 $Y=1.82 $X2=0
+ $Y2=0
cc_597 N_A_200_74#_c_551_n N_A_27_74#_c_1207_n 0.00413233f $X=1.25 $Y=1.13 $X2=0
+ $Y2=0
cc_598 N_A_200_74#_c_544_n N_A_1555_410#_M1018_g 0.040507f $X=8.125 $Y=1.22
+ $X2=0 $Y2=0
cc_599 N_A_200_74#_c_553_n N_A_1555_410#_M1018_g 0.00365403f $X=7.85 $Y=1.385
+ $X2=0 $Y2=0
cc_600 N_A_200_74#_c_553_n N_A_1555_410#_c_1402_n 0.00788658f $X=7.85 $Y=1.385
+ $X2=0 $Y2=0
cc_601 N_A_200_74#_c_544_n N_A_1335_112#_c_1607_n 0.00978321f $X=8.125 $Y=1.22
+ $X2=0 $Y2=0
cc_602 N_A_200_74#_c_547_n N_A_1335_112#_c_1607_n 0.0235121f $X=6.95 $Y=1.41
+ $X2=0 $Y2=0
cc_603 N_A_200_74#_c_549_n N_A_1335_112#_c_1607_n 0.0452891f $X=7.685 $Y=1.295
+ $X2=0 $Y2=0
cc_604 N_A_200_74#_c_552_n N_A_1335_112#_c_1607_n 0.0205478f $X=7.81 $Y=1.295
+ $X2=0 $Y2=0
cc_605 N_A_200_74#_c_553_n N_A_1335_112#_c_1607_n 0.00492308f $X=7.85 $Y=1.385
+ $X2=0 $Y2=0
cc_606 N_A_200_74#_c_554_n N_A_1335_112#_c_1607_n 0.00583385f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_607 N_A_200_74#_c_555_n N_A_1335_112#_c_1607_n 0.00233818f $X=6.96 $Y=1.295
+ $X2=0 $Y2=0
cc_608 N_A_200_74#_c_543_n N_A_1335_112#_c_1611_n 0.0138618f $X=6.905 $Y=2.045
+ $X2=0 $Y2=0
cc_609 N_A_200_74#_c_549_n N_A_1335_112#_c_1612_n 0.0102854f $X=7.685 $Y=1.295
+ $X2=0 $Y2=0
cc_610 N_A_200_74#_c_552_n N_A_1335_112#_c_1612_n 0.0179961f $X=7.81 $Y=1.295
+ $X2=0 $Y2=0
cc_611 N_A_200_74#_c_553_n N_A_1335_112#_c_1612_n 0.00502433f $X=7.85 $Y=1.385
+ $X2=0 $Y2=0
cc_612 N_A_200_74#_c_543_n N_A_1335_112#_c_1613_n 0.00104254f $X=6.905 $Y=2.045
+ $X2=0 $Y2=0
cc_613 N_A_200_74#_c_548_n N_A_1335_112#_c_1613_n 0.0143366f $X=6.95 $Y=1.745
+ $X2=0 $Y2=0
cc_614 N_A_200_74#_c_549_n N_A_1335_112#_c_1613_n 0.0077037f $X=7.685 $Y=1.295
+ $X2=0 $Y2=0
cc_615 N_A_200_74#_c_544_n N_A_1335_112#_c_1608_n 0.00925103f $X=8.125 $Y=1.22
+ $X2=0 $Y2=0
cc_616 N_A_200_74#_c_552_n N_A_1335_112#_c_1608_n 0.0266406f $X=7.81 $Y=1.295
+ $X2=0 $Y2=0
cc_617 N_A_200_74#_c_553_n N_A_1335_112#_c_1608_n 0.00728664f $X=7.85 $Y=1.385
+ $X2=0 $Y2=0
cc_618 N_A_200_74#_c_543_n N_A_1335_112#_c_1619_n 0.00579767f $X=6.905 $Y=2.045
+ $X2=0 $Y2=0
cc_619 N_A_200_74#_c_548_n N_A_1335_112#_c_1619_n 0.00913898f $X=6.95 $Y=1.745
+ $X2=0 $Y2=0
cc_620 N_A_200_74#_c_543_n N_A_1335_112#_c_1620_n 0.00292038f $X=6.905 $Y=2.045
+ $X2=0 $Y2=0
cc_621 N_A_200_74#_c_548_n N_A_1335_112#_c_1620_n 0.0014655f $X=6.95 $Y=1.745
+ $X2=0 $Y2=0
cc_622 N_A_200_74#_c_561_n N_VPWR_c_1854_n 0.0409363f $X=1.17 $Y=2.815 $X2=0
+ $Y2=0
cc_623 N_A_200_74#_c_563_n N_VPWR_c_1854_n 0.0119328f $X=1.445 $Y=2.99 $X2=0
+ $Y2=0
cc_624 N_A_200_74#_c_562_n N_VPWR_c_1855_n 0.0128702f $X=1.955 $Y=2.99 $X2=0
+ $Y2=0
cc_625 N_A_200_74#_c_565_n N_VPWR_c_1855_n 0.00209656f $X=2.975 $Y=1.77 $X2=0
+ $Y2=0
cc_626 N_A_200_74#_c_543_n N_VPWR_c_1857_n 0.00146626f $X=6.905 $Y=2.045 $X2=0
+ $Y2=0
cc_627 N_A_200_74#_c_562_n N_VPWR_c_1863_n 0.0449818f $X=1.955 $Y=2.99 $X2=0
+ $Y2=0
cc_628 N_A_200_74#_c_563_n N_VPWR_c_1863_n 0.0314532f $X=1.445 $Y=2.99 $X2=0
+ $Y2=0
cc_629 N_A_200_74#_c_559_n N_VPWR_c_1865_n 9.44495e-19 $X=3.025 $Y=2.44 $X2=0
+ $Y2=0
cc_630 N_A_200_74#_c_543_n N_VPWR_c_1870_n 0.00445602f $X=6.905 $Y=2.045 $X2=0
+ $Y2=0
cc_631 N_A_200_74#_c_543_n N_VPWR_c_1853_n 0.00858989f $X=6.905 $Y=2.045 $X2=0
+ $Y2=0
cc_632 N_A_200_74#_c_562_n N_VPWR_c_1853_n 0.025776f $X=1.955 $Y=2.99 $X2=0
+ $Y2=0
cc_633 N_A_200_74#_c_563_n N_VPWR_c_1853_n 0.0170323f $X=1.445 $Y=2.99 $X2=0
+ $Y2=0
cc_634 N_A_200_74#_c_562_n N_A_311_119#_M1039_s 0.0074246f $X=1.955 $Y=2.99
+ $X2=0 $Y2=0
cc_635 N_A_200_74#_c_562_n N_A_311_119#_c_2026_n 0.012787f $X=1.955 $Y=2.99
+ $X2=0 $Y2=0
cc_636 N_A_200_74#_c_564_n N_A_311_119#_c_2026_n 0.0624288f $X=2.04 $Y=2.905
+ $X2=0 $Y2=0
cc_637 N_A_200_74#_c_579_n N_A_311_119#_c_2026_n 0.0135851f $X=2.125 $Y=1.77
+ $X2=0 $Y2=0
cc_638 N_A_200_74#_c_550_n N_A_311_119#_c_2026_n 0.0857106f $X=1.225 $Y=1.82
+ $X2=0 $Y2=0
cc_639 N_A_200_74#_c_565_n N_A_311_119#_c_2045_n 7.39332e-19 $X=2.975 $Y=1.77
+ $X2=0 $Y2=0
cc_640 N_A_200_74#_c_554_n N_A_311_119#_c_2029_n 0.0061077f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_641 N_A_200_74#_c_554_n N_A_311_119#_c_2030_n 2.86461e-19 $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_642 N_A_200_74#_c_558_n N_A_311_119#_c_2030_n 0.00639522f $X=3.38 $Y=1.125
+ $X2=0 $Y2=0
cc_643 N_A_200_74#_c_554_n N_A_311_119#_c_2038_n 0.00348442f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_644 N_A_200_74#_c_554_n N_A_311_119#_c_2039_n 7.52032e-19 $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_645 N_A_200_74#_c_554_n N_A_311_119#_c_2031_n 0.00117028f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_646 N_A_200_74#_c_558_n N_A_311_119#_c_2031_n 0.0043128f $X=3.38 $Y=1.125
+ $X2=0 $Y2=0
cc_647 N_A_200_74#_c_554_n N_A_311_119#_c_2032_n 0.00767715f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_648 N_A_200_74#_c_545_n N_A_311_119#_c_2033_n 0.0857106f $X=1.14 $Y=0.515
+ $X2=0 $Y2=0
cc_649 N_A_200_74#_c_558_n N_A_311_119#_c_2034_n 0.00150382f $X=3.38 $Y=1.125
+ $X2=0 $Y2=0
cc_650 N_A_200_74#_c_554_n N_A_311_119#_c_2035_n 0.0166026f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_651 N_A_200_74#_c_545_n N_VGND_c_2229_n 0.0165488f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_652 N_A_200_74#_c_545_n N_VGND_c_2230_n 0.00796378f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_653 N_A_200_74#_c_554_n N_VGND_c_2231_n 0.00876862f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_654 N_A_200_74#_c_545_n N_VGND_c_2238_n 0.017299f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_655 N_A_200_74#_c_545_n N_VGND_c_2252_n 0.0127744f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_656 N_A_200_74#_c_554_n N_A_867_125#_c_2376_n 0.00640173f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_657 N_A_200_74#_c_554_n N_A_867_125#_c_2379_n 0.00876862f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_658 N_A_601_119#_c_771_n N_A_975_322#_c_878_n 0.0204332f $X=4.575 $Y=1.795
+ $X2=0 $Y2=0
cc_659 N_A_601_119#_c_778_n N_A_975_322#_c_878_n 0.00522408f $X=4.575 $Y=1.955
+ $X2=0 $Y2=0
cc_660 N_A_601_119#_c_779_n N_A_975_322#_c_878_n 0.0455164f $X=4.575 $Y=2.045
+ $X2=0 $Y2=0
cc_661 N_A_601_119#_c_771_n N_A_975_322#_M1005_g 0.00562136f $X=4.575 $Y=1.795
+ $X2=0 $Y2=0
cc_662 N_A_601_119#_c_772_n N_A_975_322#_M1005_g 0.0225897f $X=4.695 $Y=1.25
+ $X2=0 $Y2=0
cc_663 N_A_601_119#_c_771_n N_A_975_322#_c_883_n 2.65013e-19 $X=4.575 $Y=1.795
+ $X2=0 $Y2=0
cc_664 N_A_601_119#_c_771_n N_A_975_322#_c_895_n 2.95261e-19 $X=4.575 $Y=1.795
+ $X2=0 $Y2=0
cc_665 N_A_601_119#_c_775_n N_A_27_74#_M1037_g 0.00456431f $X=3.145 $Y=0.775
+ $X2=0 $Y2=0
cc_666 N_A_601_119#_c_772_n N_A_27_74#_c_1196_n 0.00737233f $X=4.695 $Y=1.25
+ $X2=0 $Y2=0
cc_667 N_A_601_119#_c_773_n N_A_27_74#_c_1209_n 0.00850319f $X=4.485 $Y=1.63
+ $X2=0 $Y2=0
cc_668 N_A_601_119#_c_781_n N_A_27_74#_c_1209_n 0.00230071f $X=3.485 $Y=2.565
+ $X2=0 $Y2=0
cc_669 N_A_601_119#_c_776_n N_A_27_74#_c_1209_n 0.00975615f $X=3.8 $Y=1.63 $X2=0
+ $Y2=0
cc_670 N_A_601_119#_c_781_n N_A_27_74#_c_1211_n 0.0182295f $X=3.485 $Y=2.565
+ $X2=0 $Y2=0
cc_671 N_A_601_119#_c_794_n N_A_27_74#_c_1212_n 0.0042982f $X=3.4 $Y=2.65 $X2=0
+ $Y2=0
cc_672 N_A_601_119#_c_781_n N_A_27_74#_c_1212_n 0.00489265f $X=3.485 $Y=2.565
+ $X2=0 $Y2=0
cc_673 N_A_601_119#_c_779_n N_VPWR_c_1856_n 0.00123641f $X=4.575 $Y=2.045 $X2=0
+ $Y2=0
cc_674 N_A_601_119#_c_779_n N_VPWR_c_1865_n 0.00333127f $X=4.575 $Y=2.045 $X2=0
+ $Y2=0
cc_675 N_A_601_119#_c_779_n N_VPWR_c_1853_n 0.00391696f $X=4.575 $Y=2.045 $X2=0
+ $Y2=0
cc_676 N_A_601_119#_c_803_n N_A_311_119#_M1023_d 0.011379f $X=3.715 $Y=0.87
+ $X2=0 $Y2=0
cc_677 N_A_601_119#_c_774_n N_A_311_119#_M1023_d 0.00189353f $X=3.8 $Y=1.465
+ $X2=0 $Y2=0
cc_678 N_A_601_119#_c_775_n N_A_311_119#_c_2045_n 0.00837589f $X=3.145 $Y=0.775
+ $X2=0 $Y2=0
cc_679 N_A_601_119#_c_775_n N_A_311_119#_c_2027_n 0.0159264f $X=3.145 $Y=0.775
+ $X2=0 $Y2=0
cc_680 N_A_601_119#_c_803_n N_A_311_119#_c_2029_n 0.0137866f $X=3.715 $Y=0.87
+ $X2=0 $Y2=0
cc_681 N_A_601_119#_c_803_n N_A_311_119#_c_2030_n 0.0161654f $X=3.715 $Y=0.87
+ $X2=0 $Y2=0
cc_682 N_A_601_119#_c_779_n N_A_311_119#_c_2037_n 0.00210001f $X=4.575 $Y=2.045
+ $X2=0 $Y2=0
cc_683 N_A_601_119#_c_794_n N_A_311_119#_c_2037_n 0.0133758f $X=3.4 $Y=2.65
+ $X2=0 $Y2=0
cc_684 N_A_601_119#_c_781_n N_A_311_119#_c_2037_n 0.031388f $X=3.485 $Y=2.565
+ $X2=0 $Y2=0
cc_685 N_A_601_119#_c_779_n N_A_311_119#_c_2038_n 0.00394305f $X=4.575 $Y=2.045
+ $X2=0 $Y2=0
cc_686 N_A_601_119#_c_773_n N_A_311_119#_c_2038_n 0.00537953f $X=4.485 $Y=1.63
+ $X2=0 $Y2=0
cc_687 N_A_601_119#_c_776_n N_A_311_119#_c_2038_n 0.00770413f $X=3.8 $Y=1.63
+ $X2=0 $Y2=0
cc_688 N_A_601_119#_c_773_n N_A_311_119#_c_2039_n 0.00122678f $X=4.485 $Y=1.63
+ $X2=0 $Y2=0
cc_689 N_A_601_119#_c_781_n N_A_311_119#_c_2039_n 0.0137412f $X=3.485 $Y=2.565
+ $X2=0 $Y2=0
cc_690 N_A_601_119#_c_776_n N_A_311_119#_c_2039_n 0.0217036f $X=3.8 $Y=1.63
+ $X2=0 $Y2=0
cc_691 N_A_601_119#_c_772_n N_A_311_119#_c_2031_n 0.00313522f $X=4.695 $Y=1.25
+ $X2=0 $Y2=0
cc_692 N_A_601_119#_c_803_n N_A_311_119#_c_2031_n 0.0136457f $X=3.715 $Y=0.87
+ $X2=0 $Y2=0
cc_693 N_A_601_119#_c_774_n N_A_311_119#_c_2031_n 0.0126048f $X=3.8 $Y=1.465
+ $X2=0 $Y2=0
cc_694 N_A_601_119#_c_771_n N_A_311_119#_c_2032_n 0.00354361f $X=4.575 $Y=1.795
+ $X2=0 $Y2=0
cc_695 N_A_601_119#_c_778_n N_A_311_119#_c_2032_n 0.00384782f $X=4.575 $Y=1.955
+ $X2=0 $Y2=0
cc_696 N_A_601_119#_c_773_n N_A_311_119#_c_2032_n 0.0204395f $X=4.485 $Y=1.63
+ $X2=0 $Y2=0
cc_697 N_A_601_119#_c_774_n N_A_311_119#_c_2032_n 0.0064903f $X=3.8 $Y=1.465
+ $X2=0 $Y2=0
cc_698 N_A_601_119#_c_776_n N_A_311_119#_c_2032_n 0.0245905f $X=3.8 $Y=1.63
+ $X2=0 $Y2=0
cc_699 N_A_601_119#_c_803_n N_A_311_119#_c_2034_n 0.0057043f $X=3.715 $Y=0.87
+ $X2=0 $Y2=0
cc_700 N_A_601_119#_c_775_n N_A_311_119#_c_2034_n 0.0198509f $X=3.145 $Y=0.775
+ $X2=0 $Y2=0
cc_701 N_A_601_119#_c_771_n N_A_311_119#_c_2035_n 8.48211e-19 $X=4.575 $Y=1.795
+ $X2=0 $Y2=0
cc_702 N_A_601_119#_c_772_n N_A_311_119#_c_2035_n 8.79985e-19 $X=4.695 $Y=1.25
+ $X2=0 $Y2=0
cc_703 N_A_601_119#_c_773_n N_A_311_119#_c_2035_n 0.00550757f $X=4.485 $Y=1.63
+ $X2=0 $Y2=0
cc_704 N_A_601_119#_c_774_n N_A_311_119#_c_2035_n 0.0129342f $X=3.8 $Y=1.465
+ $X2=0 $Y2=0
cc_705 N_A_601_119#_c_776_n N_A_311_119#_c_2035_n 0.0026112f $X=3.8 $Y=1.63
+ $X2=0 $Y2=0
cc_706 N_A_601_119#_c_771_n N_A_867_125#_c_2376_n 0.00164879f $X=4.575 $Y=1.795
+ $X2=0 $Y2=0
cc_707 N_A_601_119#_c_772_n N_A_867_125#_c_2376_n 0.00470519f $X=4.695 $Y=1.25
+ $X2=0 $Y2=0
cc_708 N_A_601_119#_c_773_n N_A_867_125#_c_2376_n 0.00254899f $X=4.485 $Y=1.63
+ $X2=0 $Y2=0
cc_709 N_A_601_119#_c_772_n N_A_867_125#_c_2377_n 0.00313969f $X=4.695 $Y=1.25
+ $X2=0 $Y2=0
cc_710 N_A_975_322#_c_878_n N_SET_B_c_1063_n 0.050395f $X=4.995 $Y=2.045
+ $X2=-0.19 $Y2=-0.245
cc_711 N_A_975_322#_c_882_n N_SET_B_c_1063_n 0.00124312f $X=6.245 $Y=1.375
+ $X2=-0.19 $Y2=-0.245
cc_712 N_A_975_322#_c_895_n N_SET_B_c_1063_n 0.00170888f $X=5.16 $Y=1.775
+ $X2=-0.19 $Y2=-0.245
cc_713 N_A_975_322#_c_878_n N_SET_B_M1003_g 6.31035e-19 $X=4.995 $Y=2.045 $X2=0
+ $Y2=0
cc_714 N_A_975_322#_M1005_g N_SET_B_M1003_g 0.0293097f $X=5.125 $Y=0.9 $X2=0
+ $Y2=0
cc_715 N_A_975_322#_c_881_n N_SET_B_M1003_g 0.00271041f $X=5.16 $Y=1.61 $X2=0
+ $Y2=0
cc_716 N_A_975_322#_c_882_n N_SET_B_M1003_g 0.0123891f $X=6.245 $Y=1.375 $X2=0
+ $Y2=0
cc_717 N_A_975_322#_c_895_n N_SET_B_M1003_g 3.82123e-19 $X=5.16 $Y=1.775 $X2=0
+ $Y2=0
cc_718 N_A_975_322#_c_880_n N_SET_B_c_1065_n 0.0104509f $X=9.58 $Y=1.795 $X2=0
+ $Y2=0
cc_719 N_A_975_322#_c_900_n N_SET_B_c_1065_n 0.0289362f $X=9.58 $Y=1.885 $X2=0
+ $Y2=0
cc_720 N_A_975_322#_c_888_n N_SET_B_c_1065_n 0.00422763f $X=9.37 $Y=1.095 $X2=0
+ $Y2=0
cc_721 N_A_975_322#_c_887_n N_SET_B_M1009_g 7.92189e-19 $X=8.53 $Y=1.01 $X2=0
+ $Y2=0
cc_722 N_A_975_322#_c_888_n N_SET_B_M1009_g 0.015521f $X=9.37 $Y=1.095 $X2=0
+ $Y2=0
cc_723 N_A_975_322#_c_890_n N_SET_B_M1009_g 0.0024163f $X=9.535 $Y=1.385 $X2=0
+ $Y2=0
cc_724 N_A_975_322#_c_891_n N_SET_B_M1009_g 0.0210337f $X=9.535 $Y=1.385 $X2=0
+ $Y2=0
cc_725 N_A_975_322#_c_897_n N_SET_B_M1009_g 0.0271518f $X=9.535 $Y=1.22 $X2=0
+ $Y2=0
cc_726 N_A_975_322#_c_880_n N_SET_B_c_1067_n 0.00127898f $X=9.58 $Y=1.795 $X2=0
+ $Y2=0
cc_727 N_A_975_322#_c_888_n N_SET_B_c_1067_n 0.020715f $X=9.37 $Y=1.095 $X2=0
+ $Y2=0
cc_728 N_A_975_322#_c_890_n N_SET_B_c_1067_n 0.00638826f $X=9.535 $Y=1.385 $X2=0
+ $Y2=0
cc_729 N_A_975_322#_c_891_n N_SET_B_c_1067_n 3.45029e-19 $X=9.535 $Y=1.385 $X2=0
+ $Y2=0
cc_730 N_A_975_322#_c_882_n N_SET_B_c_1072_n 0.0130036f $X=6.245 $Y=1.375 $X2=0
+ $Y2=0
cc_731 N_A_975_322#_c_878_n N_SET_B_c_1073_n 0.00358206f $X=4.995 $Y=2.045 $X2=0
+ $Y2=0
cc_732 N_A_975_322#_c_882_n N_SET_B_c_1073_n 0.00149199f $X=6.245 $Y=1.375 $X2=0
+ $Y2=0
cc_733 N_A_975_322#_c_895_n N_SET_B_c_1073_n 5.75947e-19 $X=5.16 $Y=1.775 $X2=0
+ $Y2=0
cc_734 N_A_975_322#_c_900_n SET_B 0.00117188f $X=9.58 $Y=1.885 $X2=0 $Y2=0
cc_735 N_A_975_322#_c_878_n N_SET_B_c_1068_n 0.00160104f $X=4.995 $Y=2.045 $X2=0
+ $Y2=0
cc_736 N_A_975_322#_c_882_n N_SET_B_c_1068_n 0.0221898f $X=6.245 $Y=1.375 $X2=0
+ $Y2=0
cc_737 N_A_975_322#_c_895_n N_SET_B_c_1068_n 0.0241405f $X=5.16 $Y=1.775 $X2=0
+ $Y2=0
cc_738 N_A_975_322#_c_880_n N_SET_B_c_1076_n 5.44528e-19 $X=9.58 $Y=1.795 $X2=0
+ $Y2=0
cc_739 N_A_975_322#_c_900_n N_SET_B_c_1076_n 0.00175205f $X=9.58 $Y=1.885 $X2=0
+ $Y2=0
cc_740 N_A_975_322#_M1005_g N_A_27_74#_c_1196_n 0.00737233f $X=5.125 $Y=0.9
+ $X2=0 $Y2=0
cc_741 N_A_975_322#_c_885_n N_A_27_74#_c_1196_n 4.42178e-19 $X=8.445 $Y=0.425
+ $X2=0 $Y2=0
cc_742 N_A_975_322#_c_886_n N_A_27_74#_c_1196_n 0.00404452f $X=6.415 $Y=0.425
+ $X2=0 $Y2=0
cc_743 N_A_975_322#_c_884_n N_A_27_74#_M1034_g 0.0112938f $X=6.33 $Y=1.29 $X2=0
+ $Y2=0
cc_744 N_A_975_322#_c_885_n N_A_27_74#_M1034_g 0.0173467f $X=8.445 $Y=0.425
+ $X2=0 $Y2=0
cc_745 N_A_975_322#_c_882_n N_A_27_74#_c_1199_n 4.12184e-19 $X=6.245 $Y=1.375
+ $X2=0 $Y2=0
cc_746 N_A_975_322#_c_892_n N_A_1555_410#_M1019_d 0.00161973f $X=10.375 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_747 N_A_975_322#_c_982_p N_A_1555_410#_M1019_d 5.72817e-19 $X=9.535 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_748 N_A_975_322#_c_885_n N_A_1555_410#_M1018_g 2.16797e-19 $X=8.445 $Y=0.425
+ $X2=0 $Y2=0
cc_749 N_A_975_322#_c_887_n N_A_1555_410#_M1018_g 0.0146703f $X=8.53 $Y=1.01
+ $X2=0 $Y2=0
cc_750 N_A_975_322#_c_889_n N_A_1555_410#_M1018_g 0.00971159f $X=8.615 $Y=1.095
+ $X2=0 $Y2=0
cc_751 N_A_975_322#_c_900_n N_A_1555_410#_c_1403_n 0.0126852f $X=9.58 $Y=1.885
+ $X2=0 $Y2=0
cc_752 N_A_975_322#_M1022_s N_A_1555_410#_c_1389_n 0.00233929f $X=10.685 $Y=0.82
+ $X2=0 $Y2=0
cc_753 N_A_975_322#_c_894_n N_A_1555_410#_c_1389_n 0.0283623f $X=10.825 $Y=1.095
+ $X2=0 $Y2=0
cc_754 N_A_975_322#_c_896_n N_A_1555_410#_c_1389_n 0.0142342f $X=10.46 $Y=1.095
+ $X2=0 $Y2=0
cc_755 N_A_975_322#_c_902_n N_A_1555_410#_c_1404_n 0.00136016f $X=10.545
+ $Y=2.035 $X2=0 $Y2=0
cc_756 N_A_975_322#_c_900_n N_A_1555_410#_c_1405_n 8.11517e-19 $X=9.58 $Y=1.885
+ $X2=0 $Y2=0
cc_757 N_A_975_322#_M1021_s N_A_1555_410#_c_1406_n 0.0117589f $X=10.625 $Y=1.84
+ $X2=0 $Y2=0
cc_758 N_A_975_322#_c_902_n N_A_1555_410#_c_1406_n 0.0130069f $X=10.545 $Y=2.035
+ $X2=0 $Y2=0
cc_759 N_A_975_322#_c_903_n N_A_1555_410#_c_1406_n 0.0231665f $X=10.755 $Y=2.035
+ $X2=0 $Y2=0
cc_760 N_A_975_322#_c_903_n N_A_1555_410#_c_1407_n 0.00710262f $X=10.755
+ $Y=2.035 $X2=0 $Y2=0
cc_761 N_A_975_322#_c_900_n N_A_1555_410#_c_1409_n 7.46086e-19 $X=9.58 $Y=1.885
+ $X2=0 $Y2=0
cc_762 N_A_975_322#_c_891_n N_A_1555_410#_c_1430_n 3.47622e-19 $X=9.535 $Y=1.385
+ $X2=0 $Y2=0
cc_763 N_A_975_322#_c_892_n N_A_1555_410#_c_1430_n 0.0402386f $X=10.375 $Y=1.095
+ $X2=0 $Y2=0
cc_764 N_A_975_322#_c_982_p N_A_1555_410#_c_1430_n 0.00434233f $X=9.535 $Y=1.095
+ $X2=0 $Y2=0
cc_765 N_A_975_322#_c_894_n N_A_1555_410#_c_1391_n 0.00851086f $X=10.825
+ $Y=1.095 $X2=0 $Y2=0
cc_766 N_A_975_322#_c_890_n N_A_1335_112#_M1008_g 0.00146389f $X=9.535 $Y=1.385
+ $X2=0 $Y2=0
cc_767 N_A_975_322#_c_891_n N_A_1335_112#_M1008_g 0.0205282f $X=9.535 $Y=1.385
+ $X2=0 $Y2=0
cc_768 N_A_975_322#_c_892_n N_A_1335_112#_M1008_g 0.0133931f $X=10.375 $Y=1.095
+ $X2=0 $Y2=0
cc_769 N_A_975_322#_c_893_n N_A_1335_112#_M1008_g 0.00578333f $X=10.46 $Y=1.95
+ $X2=0 $Y2=0
cc_770 N_A_975_322#_c_897_n N_A_1335_112#_M1008_g 0.0229225f $X=9.535 $Y=1.22
+ $X2=0 $Y2=0
cc_771 N_A_975_322#_c_880_n N_A_1335_112#_c_1606_n 0.0168437f $X=9.58 $Y=1.795
+ $X2=0 $Y2=0
cc_772 N_A_975_322#_c_900_n N_A_1335_112#_c_1606_n 0.0519304f $X=9.58 $Y=1.885
+ $X2=0 $Y2=0
cc_773 N_A_975_322#_c_892_n N_A_1335_112#_c_1606_n 0.00206847f $X=10.375
+ $Y=1.095 $X2=0 $Y2=0
cc_774 N_A_975_322#_c_893_n N_A_1335_112#_c_1606_n 0.00500819f $X=10.46 $Y=1.95
+ $X2=0 $Y2=0
cc_775 N_A_975_322#_c_902_n N_A_1335_112#_c_1606_n 0.00347021f $X=10.545
+ $Y=2.035 $X2=0 $Y2=0
cc_776 N_A_975_322#_c_884_n N_A_1335_112#_c_1607_n 0.02006f $X=6.33 $Y=1.29
+ $X2=0 $Y2=0
cc_777 N_A_975_322#_c_885_n N_A_1335_112#_c_1607_n 0.120334f $X=8.445 $Y=0.425
+ $X2=0 $Y2=0
cc_778 N_A_975_322#_c_887_n N_A_1335_112#_c_1607_n 0.0260307f $X=8.53 $Y=1.01
+ $X2=0 $Y2=0
cc_779 N_A_975_322#_c_889_n N_A_1335_112#_c_1608_n 0.0134175f $X=8.615 $Y=1.095
+ $X2=0 $Y2=0
cc_780 N_A_975_322#_c_900_n N_A_1335_112#_c_1659_n 0.0154251f $X=9.58 $Y=1.885
+ $X2=0 $Y2=0
cc_781 N_A_975_322#_c_880_n N_A_1335_112#_c_1609_n 0.00501277f $X=9.58 $Y=1.795
+ $X2=0 $Y2=0
cc_782 N_A_975_322#_c_890_n N_A_1335_112#_c_1609_n 0.00504849f $X=9.535 $Y=1.385
+ $X2=0 $Y2=0
cc_783 N_A_975_322#_c_891_n N_A_1335_112#_c_1609_n 2.79183e-19 $X=9.535 $Y=1.385
+ $X2=0 $Y2=0
cc_784 N_A_975_322#_c_892_n N_A_1335_112#_c_1609_n 0.0217264f $X=10.375 $Y=1.095
+ $X2=0 $Y2=0
cc_785 N_A_975_322#_c_893_n N_A_1335_112#_c_1609_n 0.0323382f $X=10.46 $Y=1.95
+ $X2=0 $Y2=0
cc_786 N_A_975_322#_c_900_n N_A_1335_112#_c_1618_n 0.00933466f $X=9.58 $Y=1.885
+ $X2=0 $Y2=0
cc_787 N_A_975_322#_c_893_n N_A_1335_112#_c_1618_n 0.00213745f $X=10.46 $Y=1.95
+ $X2=0 $Y2=0
cc_788 N_A_975_322#_c_902_n N_A_1335_112#_c_1618_n 0.00385646f $X=10.545
+ $Y=2.035 $X2=0 $Y2=0
cc_789 N_A_975_322#_c_889_n N_A_1335_112#_c_1621_n 0.00444169f $X=8.615 $Y=1.095
+ $X2=0 $Y2=0
cc_790 N_A_975_322#_c_893_n N_RESET_B_c_1744_n 0.0046883f $X=10.46 $Y=1.95
+ $X2=-0.19 $Y2=-0.245
cc_791 N_A_975_322#_c_894_n N_RESET_B_c_1744_n 0.00113847f $X=10.825 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_792 N_A_975_322#_c_903_n N_RESET_B_c_1744_n 0.00326168f $X=10.755 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_793 N_A_975_322#_c_893_n N_RESET_B_c_1745_n 0.00366428f $X=10.46 $Y=1.95
+ $X2=0 $Y2=0
cc_794 N_A_975_322#_c_894_n N_RESET_B_c_1745_n 0.00290255f $X=10.825 $Y=1.095
+ $X2=0 $Y2=0
cc_795 N_A_975_322#_c_893_n N_RESET_B_c_1746_n 0.0346172f $X=10.46 $Y=1.95 $X2=0
+ $Y2=0
cc_796 N_A_975_322#_c_894_n N_RESET_B_c_1746_n 0.018879f $X=10.825 $Y=1.095
+ $X2=0 $Y2=0
cc_797 N_A_975_322#_c_903_n N_RESET_B_c_1746_n 0.0141111f $X=10.755 $Y=2.035
+ $X2=0 $Y2=0
cc_798 N_A_975_322#_c_878_n N_VPWR_c_1856_n 0.00871859f $X=4.995 $Y=2.045 $X2=0
+ $Y2=0
cc_799 N_A_975_322#_c_878_n N_VPWR_c_1865_n 0.00413917f $X=4.995 $Y=2.045 $X2=0
+ $Y2=0
cc_800 N_A_975_322#_c_900_n N_VPWR_c_1873_n 0.00314375f $X=9.58 $Y=1.885 $X2=0
+ $Y2=0
cc_801 N_A_975_322#_c_900_n N_VPWR_c_1878_n 0.00330333f $X=9.58 $Y=1.885 $X2=0
+ $Y2=0
cc_802 N_A_975_322#_c_878_n N_VPWR_c_1853_n 0.00414311f $X=4.995 $Y=2.045 $X2=0
+ $Y2=0
cc_803 N_A_975_322#_c_900_n N_VPWR_c_1853_n 0.00390476f $X=9.58 $Y=1.885 $X2=0
+ $Y2=0
cc_804 N_A_975_322#_c_888_n N_VGND_M1018_d 0.00740764f $X=9.37 $Y=1.095 $X2=0
+ $Y2=0
cc_805 N_A_975_322#_c_882_n N_VGND_c_2231_n 0.0130241f $X=6.245 $Y=1.375 $X2=0
+ $Y2=0
cc_806 N_A_975_322#_c_884_n N_VGND_c_2231_n 0.0235755f $X=6.33 $Y=1.29 $X2=0
+ $Y2=0
cc_807 N_A_975_322#_c_886_n N_VGND_c_2231_n 0.0149762f $X=6.415 $Y=0.425 $X2=0
+ $Y2=0
cc_808 N_A_975_322#_c_885_n N_VGND_c_2232_n 0.0141715f $X=8.445 $Y=0.425 $X2=0
+ $Y2=0
cc_809 N_A_975_322#_c_887_n N_VGND_c_2232_n 0.0186856f $X=8.53 $Y=1.01 $X2=0
+ $Y2=0
cc_810 N_A_975_322#_c_888_n N_VGND_c_2232_n 0.0135869f $X=9.37 $Y=1.095 $X2=0
+ $Y2=0
cc_811 N_A_975_322#_c_885_n N_VGND_c_2240_n 0.0927715f $X=8.445 $Y=0.425 $X2=0
+ $Y2=0
cc_812 N_A_975_322#_c_886_n N_VGND_c_2240_n 0.00789578f $X=6.415 $Y=0.425 $X2=0
+ $Y2=0
cc_813 N_A_975_322#_c_897_n N_VGND_c_2248_n 0.00278271f $X=9.535 $Y=1.22 $X2=0
+ $Y2=0
cc_814 N_A_975_322#_c_885_n N_VGND_c_2252_n 0.0774033f $X=8.445 $Y=0.425 $X2=0
+ $Y2=0
cc_815 N_A_975_322#_c_886_n N_VGND_c_2252_n 0.00563471f $X=6.415 $Y=0.425 $X2=0
+ $Y2=0
cc_816 N_A_975_322#_c_897_n N_VGND_c_2252_n 0.00353984f $X=9.535 $Y=1.22 $X2=0
+ $Y2=0
cc_817 N_A_975_322#_M1005_g N_A_867_125#_c_2377_n 0.00330783f $X=5.125 $Y=0.9
+ $X2=0 $Y2=0
cc_818 N_A_975_322#_M1005_g N_A_867_125#_c_2379_n 0.00537237f $X=5.125 $Y=0.9
+ $X2=0 $Y2=0
cc_819 N_A_975_322#_c_882_n N_A_867_125#_c_2379_n 0.0130241f $X=6.245 $Y=1.375
+ $X2=0 $Y2=0
cc_820 N_A_975_322#_c_884_n A_1240_125# 0.0106247f $X=6.33 $Y=1.29 $X2=-0.19
+ $Y2=-0.245
cc_821 N_A_975_322#_c_888_n N_A_1832_74#_M1009_d 0.00161579f $X=9.37 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_822 N_A_975_322#_c_892_n N_A_1832_74#_M1008_d 0.0034729f $X=10.375 $Y=1.095
+ $X2=0 $Y2=0
cc_823 N_A_975_322#_c_896_n N_A_1832_74#_M1008_d 6.6514e-19 $X=10.46 $Y=1.095
+ $X2=0 $Y2=0
cc_824 N_A_975_322#_c_888_n N_A_1832_74#_c_2416_n 0.0140651f $X=9.37 $Y=1.095
+ $X2=0 $Y2=0
cc_825 N_A_975_322#_c_982_p N_A_1832_74#_c_2416_n 0.00114098f $X=9.535 $Y=1.095
+ $X2=0 $Y2=0
cc_826 N_A_975_322#_c_982_p N_A_1832_74#_c_2412_n 0.00401745f $X=9.535 $Y=1.095
+ $X2=0 $Y2=0
cc_827 N_A_975_322#_c_897_n N_A_1832_74#_c_2412_n 0.0109934f $X=9.535 $Y=1.22
+ $X2=0 $Y2=0
cc_828 N_SET_B_M1003_g N_A_27_74#_c_1196_n 0.00879826f $X=5.625 $Y=0.9 $X2=0
+ $Y2=0
cc_829 N_SET_B_c_1072_n N_A_27_74#_c_1199_n 0.00232724f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_830 N_SET_B_c_1072_n N_A_27_74#_c_1213_n 0.00518867f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_831 N_SET_B_c_1072_n N_A_1555_410#_M1030_s 0.00644023f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_832 SET_B N_A_1555_410#_M1030_s 0.00161567f $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_833 N_SET_B_c_1076_n N_A_1555_410#_M1030_s 0.00105183f $X=8.88 $Y=2.035 $X2=0
+ $Y2=0
cc_834 N_SET_B_c_1065_n N_A_1555_410#_c_1393_n 0.0100531f $X=8.96 $Y=1.885 $X2=0
+ $Y2=0
cc_835 N_SET_B_c_1072_n N_A_1555_410#_c_1393_n 0.00289299f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_836 N_SET_B_c_1076_n N_A_1555_410#_c_1393_n 2.8668e-19 $X=8.88 $Y=2.035 $X2=0
+ $Y2=0
cc_837 N_SET_B_c_1065_n N_A_1555_410#_M1018_g 0.0167528f $X=8.96 $Y=1.885 $X2=0
+ $Y2=0
cc_838 N_SET_B_M1009_g N_A_1555_410#_M1018_g 0.0220493f $X=9.085 $Y=0.74 $X2=0
+ $Y2=0
cc_839 N_SET_B_c_1067_n N_A_1555_410#_M1018_g 0.00280077f $X=8.995 $Y=1.615
+ $X2=0 $Y2=0
cc_840 N_SET_B_c_1065_n N_A_1555_410#_c_1400_n 0.00475092f $X=8.96 $Y=1.885
+ $X2=0 $Y2=0
cc_841 N_SET_B_c_1076_n N_A_1555_410#_c_1400_n 3.42051e-19 $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_842 N_SET_B_c_1065_n N_A_1555_410#_c_1401_n 0.00402606f $X=8.96 $Y=1.885
+ $X2=0 $Y2=0
cc_843 N_SET_B_c_1072_n N_A_1555_410#_c_1401_n 0.0221024f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_844 N_SET_B_c_1072_n N_A_1555_410#_c_1402_n 0.0111728f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_845 N_SET_B_c_1065_n N_A_1555_410#_c_1403_n 0.00834124f $X=8.96 $Y=1.885
+ $X2=0 $Y2=0
cc_846 N_SET_B_c_1072_n N_A_1555_410#_c_1408_n 0.00563301f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_847 N_SET_B_c_1065_n N_A_1555_410#_c_1409_n 0.00451111f $X=8.96 $Y=1.885
+ $X2=0 $Y2=0
cc_848 N_SET_B_c_1072_n N_A_1555_410#_c_1409_n 2.71663e-19 $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_849 N_SET_B_c_1072_n N_A_1335_112#_c_1612_n 0.0396252f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_850 N_SET_B_c_1067_n N_A_1335_112#_c_1608_n 0.0103489f $X=8.995 $Y=1.615
+ $X2=0 $Y2=0
cc_851 N_SET_B_c_1065_n N_A_1335_112#_c_1615_n 0.00383423f $X=8.96 $Y=1.885
+ $X2=0 $Y2=0
cc_852 N_SET_B_c_1072_n N_A_1335_112#_c_1615_n 0.0123221f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_853 SET_B N_A_1335_112#_c_1615_n 0.00328463f $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_854 N_SET_B_c_1076_n N_A_1335_112#_c_1615_n 0.0158868f $X=8.88 $Y=2.035 $X2=0
+ $Y2=0
cc_855 N_SET_B_c_1065_n N_A_1335_112#_c_1659_n 0.0149225f $X=8.96 $Y=1.885 $X2=0
+ $Y2=0
cc_856 N_SET_B_c_1067_n N_A_1335_112#_c_1659_n 0.00370079f $X=8.995 $Y=1.615
+ $X2=0 $Y2=0
cc_857 N_SET_B_c_1072_n N_A_1335_112#_c_1659_n 0.00621792f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_858 SET_B N_A_1335_112#_c_1659_n 0.00838952f $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_859 N_SET_B_c_1076_n N_A_1335_112#_c_1659_n 0.0115811f $X=8.88 $Y=2.035 $X2=0
+ $Y2=0
cc_860 N_SET_B_c_1067_n N_A_1335_112#_c_1609_n 0.00198315f $X=8.995 $Y=1.615
+ $X2=0 $Y2=0
cc_861 N_SET_B_c_1072_n N_A_1335_112#_c_1619_n 0.031922f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_862 N_SET_B_c_1072_n N_A_1335_112#_c_1620_n 0.013405f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_863 N_SET_B_c_1065_n N_A_1335_112#_c_1621_n 5.23151e-19 $X=8.96 $Y=1.885
+ $X2=0 $Y2=0
cc_864 N_SET_B_c_1067_n N_A_1335_112#_c_1621_n 0.00521962f $X=8.995 $Y=1.615
+ $X2=0 $Y2=0
cc_865 N_SET_B_c_1072_n N_A_1335_112#_c_1621_n 0.00138583f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_866 N_SET_B_c_1076_n N_A_1335_112#_c_1621_n 0.00939718f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_867 N_SET_B_c_1073_n N_VPWR_M1017_d 7.43795e-19 $X=5.665 $Y=2.035 $X2=0 $Y2=0
cc_868 N_SET_B_c_1063_n N_VPWR_c_1856_n 0.0048817f $X=5.505 $Y=2.045 $X2=0 $Y2=0
cc_869 N_SET_B_c_1063_n N_VPWR_c_1857_n 0.00334101f $X=5.505 $Y=2.045 $X2=0
+ $Y2=0
cc_870 N_SET_B_c_1072_n N_VPWR_c_1857_n 0.00148621f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_871 N_SET_B_c_1063_n N_VPWR_c_1867_n 0.00445602f $X=5.505 $Y=2.045 $X2=0
+ $Y2=0
cc_872 N_SET_B_c_1065_n N_VPWR_c_1869_n 0.00276611f $X=8.96 $Y=1.885 $X2=0 $Y2=0
cc_873 N_SET_B_c_1065_n N_VPWR_c_1872_n 0.00361132f $X=8.96 $Y=1.885 $X2=0 $Y2=0
cc_874 N_SET_B_c_1065_n N_VPWR_c_1878_n 0.00326445f $X=8.96 $Y=1.885 $X2=0 $Y2=0
cc_875 N_SET_B_c_1063_n N_VPWR_c_1853_n 0.00459317f $X=5.505 $Y=2.045 $X2=0
+ $Y2=0
cc_876 N_SET_B_c_1065_n N_VPWR_c_1853_n 0.00565696f $X=8.96 $Y=1.885 $X2=0 $Y2=0
cc_877 N_SET_B_M1003_g N_VGND_c_2231_n 0.00318941f $X=5.625 $Y=0.9 $X2=0 $Y2=0
cc_878 N_SET_B_M1009_g N_VGND_c_2232_n 0.0039612f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_879 N_SET_B_M1009_g N_VGND_c_2248_n 0.00430908f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_880 N_SET_B_M1003_g N_VGND_c_2252_n 7.94319e-19 $X=5.625 $Y=0.9 $X2=0 $Y2=0
cc_881 N_SET_B_M1009_g N_VGND_c_2252_n 0.00820779f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_882 N_SET_B_M1003_g N_A_867_125#_c_2379_n 0.0080727f $X=5.625 $Y=0.9 $X2=0
+ $Y2=0
cc_883 N_SET_B_M1009_g N_A_1832_74#_c_2416_n 0.00521098f $X=9.085 $Y=0.74 $X2=0
+ $Y2=0
cc_884 N_SET_B_M1009_g N_A_1832_74#_c_2410_n 0.00368587f $X=9.085 $Y=0.74 $X2=0
+ $Y2=0
cc_885 N_A_27_74#_c_1214_n N_A_1555_410#_c_1392_n 0.0276298f $X=7.445 $Y=2.465
+ $X2=0 $Y2=0
cc_886 N_A_27_74#_c_1213_n N_A_1555_410#_c_1393_n 0.00186083f $X=7.445 $Y=2.375
+ $X2=0 $Y2=0
cc_887 N_A_27_74#_c_1216_n N_A_1555_410#_c_1400_n 0.00186083f $X=7.43 $Y=1.94
+ $X2=0 $Y2=0
cc_888 N_A_27_74#_c_1213_n N_A_1555_410#_c_1401_n 0.0011224f $X=7.445 $Y=2.375
+ $X2=0 $Y2=0
cc_889 N_A_27_74#_c_1214_n N_A_1555_410#_c_1401_n 4.58089e-19 $X=7.445 $Y=2.465
+ $X2=0 $Y2=0
cc_890 N_A_27_74#_c_1213_n N_A_1555_410#_c_1402_n 0.0225952f $X=7.445 $Y=2.375
+ $X2=0 $Y2=0
cc_891 N_A_27_74#_c_1214_n N_A_1555_410#_c_1458_n 4.73961e-19 $X=7.445 $Y=2.465
+ $X2=0 $Y2=0
cc_892 N_A_27_74#_M1034_g N_A_1335_112#_c_1607_n 0.00457109f $X=6.6 $Y=0.835
+ $X2=0 $Y2=0
cc_893 N_A_27_74#_c_1198_n N_A_1335_112#_c_1607_n 0.00798476f $X=7.325 $Y=1.26
+ $X2=0 $Y2=0
cc_894 N_A_27_74#_c_1213_n N_A_1335_112#_c_1611_n 0.00103163f $X=7.445 $Y=2.375
+ $X2=0 $Y2=0
cc_895 N_A_27_74#_c_1214_n N_A_1335_112#_c_1611_n 0.0232475f $X=7.445 $Y=2.465
+ $X2=0 $Y2=0
cc_896 N_A_27_74#_c_1201_n N_A_1335_112#_c_1612_n 0.00212009f $X=7.43 $Y=1.79
+ $X2=0 $Y2=0
cc_897 N_A_27_74#_c_1216_n N_A_1335_112#_c_1612_n 0.00488542f $X=7.43 $Y=1.94
+ $X2=0 $Y2=0
cc_898 N_A_27_74#_c_1198_n N_A_1335_112#_c_1613_n 2.53696e-19 $X=7.325 $Y=1.26
+ $X2=0 $Y2=0
cc_899 N_A_27_74#_c_1201_n N_A_1335_112#_c_1613_n 0.00363368f $X=7.43 $Y=1.79
+ $X2=0 $Y2=0
cc_900 N_A_27_74#_c_1216_n N_A_1335_112#_c_1613_n 0.00147317f $X=7.43 $Y=1.94
+ $X2=0 $Y2=0
cc_901 N_A_27_74#_c_1201_n N_A_1335_112#_c_1608_n 0.00361586f $X=7.43 $Y=1.79
+ $X2=0 $Y2=0
cc_902 N_A_27_74#_c_1213_n N_A_1335_112#_c_1619_n 0.00900591f $X=7.445 $Y=2.375
+ $X2=0 $Y2=0
cc_903 N_A_27_74#_c_1213_n N_A_1335_112#_c_1620_n 0.00556844f $X=7.445 $Y=2.375
+ $X2=0 $Y2=0
cc_904 N_A_27_74#_c_1216_n N_A_1335_112#_c_1620_n 0.00339441f $X=7.43 $Y=1.94
+ $X2=0 $Y2=0
cc_905 N_A_27_74#_c_1232_n N_VPWR_M1028_d 0.00454793f $X=0.665 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_906 N_A_27_74#_c_1206_n N_VPWR_M1028_d 0.0015936f $X=0.75 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_907 N_A_27_74#_c_1192_n N_VPWR_c_1854_n 0.00334369f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_908 N_A_27_74#_c_1218_n N_VPWR_c_1854_n 0.0449718f $X=0.27 $Y=2.815 $X2=0
+ $Y2=0
cc_909 N_A_27_74#_c_1232_n N_VPWR_c_1854_n 0.0145152f $X=0.665 $Y=2.035 $X2=0
+ $Y2=0
cc_910 N_A_27_74#_c_1192_n N_VPWR_c_1863_n 0.0044313f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_911 N_A_27_74#_c_1212_n N_VPWR_c_1865_n 9.44495e-19 $X=3.535 $Y=2.44 $X2=0
+ $Y2=0
cc_912 N_A_27_74#_c_1214_n N_VPWR_c_1870_n 0.00366292f $X=7.445 $Y=2.465 $X2=0
+ $Y2=0
cc_913 N_A_27_74#_c_1218_n N_VPWR_c_1871_n 0.0145938f $X=0.27 $Y=2.815 $X2=0
+ $Y2=0
cc_914 N_A_27_74#_c_1192_n N_VPWR_c_1853_n 0.00858246f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_915 N_A_27_74#_c_1214_n N_VPWR_c_1853_n 0.00639614f $X=7.445 $Y=2.465 $X2=0
+ $Y2=0
cc_916 N_A_27_74#_c_1218_n N_VPWR_c_1853_n 0.0120466f $X=0.27 $Y=2.815 $X2=0
+ $Y2=0
cc_917 N_A_27_74#_c_1192_n N_A_311_119#_c_2026_n 0.00166814f $X=0.945 $Y=1.765
+ $X2=0 $Y2=0
cc_918 N_A_27_74#_c_1193_n N_A_311_119#_c_2045_n 0.00196569f $X=2.855 $Y=0.18
+ $X2=0 $Y2=0
cc_919 N_A_27_74#_M1037_g N_A_311_119#_c_2045_n 0.0025009f $X=2.93 $Y=0.805
+ $X2=0 $Y2=0
cc_920 N_A_27_74#_M1037_g N_A_311_119#_c_2027_n 0.00592273f $X=2.93 $Y=0.805
+ $X2=0 $Y2=0
cc_921 N_A_27_74#_c_1193_n N_A_311_119#_c_2028_n 0.00466053f $X=2.855 $Y=0.18
+ $X2=0 $Y2=0
cc_922 N_A_27_74#_c_1196_n N_A_311_119#_c_2029_n 0.00420304f $X=6.525 $Y=0.18
+ $X2=0 $Y2=0
cc_923 N_A_27_74#_M1037_g N_A_311_119#_c_2030_n 0.00142422f $X=2.93 $Y=0.805
+ $X2=0 $Y2=0
cc_924 N_A_27_74#_c_1211_n N_A_311_119#_c_2037_n 0.00649889f $X=3.535 $Y=2.35
+ $X2=0 $Y2=0
cc_925 N_A_27_74#_c_1212_n N_A_311_119#_c_2037_n 0.00595216f $X=3.535 $Y=2.44
+ $X2=0 $Y2=0
cc_926 N_A_27_74#_c_1211_n N_A_311_119#_c_2039_n 0.0037565f $X=3.535 $Y=2.35
+ $X2=0 $Y2=0
cc_927 N_A_27_74#_c_1209_n N_A_311_119#_c_2032_n 0.00376037f $X=3.445 $Y=1.74
+ $X2=0 $Y2=0
cc_928 N_A_27_74#_M1033_g N_A_311_119#_c_2033_n 0.0012846f $X=0.925 $Y=0.74
+ $X2=0 $Y2=0
cc_929 N_A_27_74#_c_1193_n N_A_311_119#_c_2033_n 0.00458356f $X=2.855 $Y=0.18
+ $X2=0 $Y2=0
cc_930 N_A_27_74#_M1037_g N_A_311_119#_c_2034_n 0.0146966f $X=2.93 $Y=0.805
+ $X2=0 $Y2=0
cc_931 N_A_27_74#_c_1196_n N_A_311_119#_c_2034_n 0.0203618f $X=6.525 $Y=0.18
+ $X2=0 $Y2=0
cc_932 N_A_27_74#_c_1203_n N_VGND_M1032_d 0.00210254f $X=0.665 $Y=1.045
+ $X2=-0.19 $Y2=-0.245
cc_933 N_A_27_74#_M1033_g N_VGND_c_2229_n 0.0115341f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_934 N_A_27_74#_c_1194_n N_VGND_c_2229_n 0.0075099f $X=1 $Y=0.18 $X2=0 $Y2=0
cc_935 N_A_27_74#_c_1202_n N_VGND_c_2229_n 0.0164982f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_936 N_A_27_74#_c_1203_n N_VGND_c_2229_n 0.0158226f $X=0.665 $Y=1.045 $X2=0
+ $Y2=0
cc_937 N_A_27_74#_c_1207_n N_VGND_c_2229_n 0.00102653f $X=0.96 $Y=1.465 $X2=0
+ $Y2=0
cc_938 N_A_27_74#_c_1193_n N_VGND_c_2230_n 0.0288848f $X=2.855 $Y=0.18 $X2=0
+ $Y2=0
cc_939 N_A_27_74#_M1037_g N_VGND_c_2230_n 8.09569e-19 $X=2.93 $Y=0.805 $X2=0
+ $Y2=0
cc_940 N_A_27_74#_c_1196_n N_VGND_c_2231_n 0.0257192f $X=6.525 $Y=0.18 $X2=0
+ $Y2=0
cc_941 N_A_27_74#_M1034_g N_VGND_c_2231_n 0.00311462f $X=6.6 $Y=0.835 $X2=0
+ $Y2=0
cc_942 N_A_27_74#_c_1202_n N_VGND_c_2237_n 0.011066f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_943 N_A_27_74#_c_1194_n N_VGND_c_2238_n 0.0338441f $X=1 $Y=0.18 $X2=0 $Y2=0
cc_944 N_A_27_74#_c_1193_n N_VGND_c_2239_n 0.0755745f $X=2.855 $Y=0.18 $X2=0
+ $Y2=0
cc_945 N_A_27_74#_c_1196_n N_VGND_c_2240_n 0.016002f $X=6.525 $Y=0.18 $X2=0
+ $Y2=0
cc_946 N_A_27_74#_c_1193_n N_VGND_c_2252_n 0.0440749f $X=2.855 $Y=0.18 $X2=0
+ $Y2=0
cc_947 N_A_27_74#_c_1194_n N_VGND_c_2252_n 0.00749832f $X=1 $Y=0.18 $X2=0 $Y2=0
cc_948 N_A_27_74#_c_1196_n N_VGND_c_2252_n 0.0907427f $X=6.525 $Y=0.18 $X2=0
+ $Y2=0
cc_949 N_A_27_74#_c_1200_n N_VGND_c_2252_n 0.00370846f $X=2.93 $Y=0.18 $X2=0
+ $Y2=0
cc_950 N_A_27_74#_c_1202_n N_VGND_c_2252_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_951 N_A_27_74#_c_1196_n N_A_867_125#_c_2377_n 0.0187725f $X=6.525 $Y=0.18
+ $X2=0 $Y2=0
cc_952 N_A_27_74#_c_1196_n N_A_867_125#_c_2378_n 0.00418041f $X=6.525 $Y=0.18
+ $X2=0 $Y2=0
cc_953 N_A_1555_410#_c_1389_n N_A_1335_112#_M1008_g 0.00974059f $X=11.29
+ $Y=0.755 $X2=0 $Y2=0
cc_954 N_A_1555_410#_c_1430_n N_A_1335_112#_M1008_g 0.00425977f $X=9.935
+ $Y=0.717 $X2=0 $Y2=0
cc_955 N_A_1555_410#_c_1403_n N_A_1335_112#_c_1606_n 0.015744f $X=10.06 $Y=2.715
+ $X2=0 $Y2=0
cc_956 N_A_1555_410#_c_1404_n N_A_1335_112#_c_1606_n 0.0035506f $X=10.225
+ $Y=2.46 $X2=0 $Y2=0
cc_957 N_A_1555_410#_c_1405_n N_A_1335_112#_c_1606_n 0.00291953f $X=10.225
+ $Y=2.63 $X2=0 $Y2=0
cc_958 N_A_1555_410#_M1018_g N_A_1335_112#_c_1607_n 0.00198618f $X=8.515 $Y=0.9
+ $X2=0 $Y2=0
cc_959 N_A_1555_410#_c_1392_n N_A_1335_112#_c_1611_n 0.00203875f $X=7.865
+ $Y=2.465 $X2=0 $Y2=0
cc_960 N_A_1555_410#_c_1458_n N_A_1335_112#_c_1611_n 0.00609671f $X=8.255
+ $Y=2.715 $X2=0 $Y2=0
cc_961 N_A_1555_410#_c_1401_n N_A_1335_112#_c_1612_n 0.0204961f $X=8.09 $Y=2.215
+ $X2=0 $Y2=0
cc_962 N_A_1555_410#_c_1402_n N_A_1335_112#_c_1612_n 0.00665045f $X=8.09
+ $Y=2.215 $X2=0 $Y2=0
cc_963 N_A_1555_410#_M1018_g N_A_1335_112#_c_1608_n 0.0114225f $X=8.515 $Y=0.9
+ $X2=0 $Y2=0
cc_964 N_A_1555_410#_c_1400_n N_A_1335_112#_c_1608_n 3.02029e-19 $X=8.515
+ $Y=1.81 $X2=0 $Y2=0
cc_965 N_A_1555_410#_M1030_s N_A_1335_112#_c_1615_n 0.0027694f $X=8.59 $Y=1.96
+ $X2=0 $Y2=0
cc_966 N_A_1555_410#_c_1393_n N_A_1335_112#_c_1615_n 0.00718671f $X=8.33 $Y=2.05
+ $X2=0 $Y2=0
cc_967 N_A_1555_410#_c_1400_n N_A_1335_112#_c_1615_n 0.00424677f $X=8.515
+ $Y=1.81 $X2=0 $Y2=0
cc_968 N_A_1555_410#_c_1401_n N_A_1335_112#_c_1615_n 0.0167912f $X=8.09 $Y=2.215
+ $X2=0 $Y2=0
cc_969 N_A_1555_410#_M1030_s N_A_1335_112#_c_1659_n 0.00628628f $X=8.59 $Y=1.96
+ $X2=0 $Y2=0
cc_970 N_A_1555_410#_c_1403_n N_A_1335_112#_c_1659_n 0.0119962f $X=10.06
+ $Y=2.715 $X2=0 $Y2=0
cc_971 N_A_1555_410#_c_1409_n N_A_1335_112#_c_1659_n 0.0639282f $X=8.9 $Y=2.805
+ $X2=0 $Y2=0
cc_972 N_A_1555_410#_c_1401_n N_A_1335_112#_c_1616_n 0.0146656f $X=8.09 $Y=2.215
+ $X2=0 $Y2=0
cc_973 N_A_1555_410#_c_1402_n N_A_1335_112#_c_1616_n 0.0016f $X=8.09 $Y=2.215
+ $X2=0 $Y2=0
cc_974 N_A_1555_410#_c_1408_n N_A_1335_112#_c_1616_n 0.0137507f $X=8.57 $Y=2.805
+ $X2=0 $Y2=0
cc_975 N_A_1555_410#_c_1404_n N_A_1335_112#_c_1609_n 0.00546019f $X=10.225
+ $Y=2.46 $X2=0 $Y2=0
cc_976 N_A_1555_410#_c_1401_n N_A_1335_112#_c_1620_n 0.018468f $X=8.09 $Y=2.215
+ $X2=0 $Y2=0
cc_977 N_A_1555_410#_c_1402_n N_A_1335_112#_c_1620_n 0.00160183f $X=8.09
+ $Y=2.215 $X2=0 $Y2=0
cc_978 N_A_1555_410#_c_1393_n N_A_1335_112#_c_1621_n 0.00209883f $X=8.33 $Y=2.05
+ $X2=0 $Y2=0
cc_979 N_A_1555_410#_M1018_g N_A_1335_112#_c_1621_n 0.00445785f $X=8.515 $Y=0.9
+ $X2=0 $Y2=0
cc_980 N_A_1555_410#_c_1400_n N_A_1335_112#_c_1621_n 0.0136664f $X=8.515 $Y=1.81
+ $X2=0 $Y2=0
cc_981 N_A_1555_410#_c_1395_n N_RESET_B_c_1744_n 0.0247602f $X=11.505 $Y=1.765
+ $X2=-0.19 $Y2=-0.245
cc_982 N_A_1555_410#_c_1386_n N_RESET_B_c_1744_n 0.0236424f $X=12.085 $Y=1.515
+ $X2=-0.19 $Y2=-0.245
cc_983 N_A_1555_410#_c_1405_n N_RESET_B_c_1744_n 0.00386334f $X=10.225 $Y=2.63
+ $X2=-0.19 $Y2=-0.245
cc_984 N_A_1555_410#_c_1406_n N_RESET_B_c_1744_n 0.0183081f $X=11.29 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_985 N_A_1555_410#_c_1407_n N_RESET_B_c_1744_n 0.00840899f $X=11.375 $Y=2.29
+ $X2=-0.19 $Y2=-0.245
cc_986 N_A_1555_410#_c_1390_n N_RESET_B_c_1744_n 0.00530017f $X=11.49 $Y=1.515
+ $X2=-0.19 $Y2=-0.245
cc_987 N_A_1555_410#_c_1383_n N_RESET_B_c_1745_n 0.0148378f $X=11.58 $Y=1.35
+ $X2=0 $Y2=0
cc_988 N_A_1555_410#_c_1389_n N_RESET_B_c_1745_n 0.0132667f $X=11.29 $Y=0.755
+ $X2=0 $Y2=0
cc_989 N_A_1555_410#_c_1391_n N_RESET_B_c_1745_n 0.00530017f $X=11.467 $Y=1.35
+ $X2=0 $Y2=0
cc_990 N_A_1555_410#_c_1386_n N_RESET_B_c_1746_n 6.27139e-19 $X=12.085 $Y=1.515
+ $X2=0 $Y2=0
cc_991 N_A_1555_410#_c_1389_n N_RESET_B_c_1746_n 0.00369733f $X=11.29 $Y=0.755
+ $X2=0 $Y2=0
cc_992 N_A_1555_410#_c_1406_n N_RESET_B_c_1746_n 0.00525533f $X=11.29 $Y=2.375
+ $X2=0 $Y2=0
cc_993 N_A_1555_410#_c_1390_n N_RESET_B_c_1746_n 0.0339135f $X=11.49 $Y=1.515
+ $X2=0 $Y2=0
cc_994 N_A_1555_410#_c_1387_n N_A_2516_368#_c_1780_n 0.0160629f $X=12.935
+ $Y=1.765 $X2=0 $Y2=0
cc_995 N_A_1555_410#_M1025_g N_A_2516_368#_M1006_g 0.0122368f $X=13.015 $Y=0.69
+ $X2=0 $Y2=0
cc_996 N_A_1555_410#_c_1396_n N_A_2516_368#_c_1782_n 0.00720368f $X=11.955
+ $Y=1.765 $X2=0 $Y2=0
cc_997 N_A_1555_410#_c_1385_n N_A_2516_368#_c_1782_n 0.00408594f $X=12.845
+ $Y=1.515 $X2=0 $Y2=0
cc_998 N_A_1555_410#_c_1387_n N_A_2516_368#_c_1782_n 0.00203522f $X=12.935
+ $Y=1.765 $X2=0 $Y2=0
cc_999 N_A_1555_410#_c_1396_n N_A_2516_368#_c_1783_n 0.00121495f $X=11.955
+ $Y=1.765 $X2=0 $Y2=0
cc_1000 N_A_1555_410#_c_1387_n N_A_2516_368#_c_1783_n 0.00933691f $X=12.935
+ $Y=1.765 $X2=0 $Y2=0
cc_1001 N_A_1555_410#_c_1384_n N_A_2516_368#_c_1776_n 0.00156292f $X=12.01
+ $Y=1.35 $X2=0 $Y2=0
cc_1002 N_A_1555_410#_M1025_g N_A_2516_368#_c_1776_n 0.00969293f $X=13.015
+ $Y=0.69 $X2=0 $Y2=0
cc_1003 N_A_1555_410#_c_1387_n N_A_2516_368#_c_1777_n 0.0149276f $X=12.935
+ $Y=1.765 $X2=0 $Y2=0
cc_1004 N_A_1555_410#_M1025_g N_A_2516_368#_c_1777_n 0.0107369f $X=13.015
+ $Y=0.69 $X2=0 $Y2=0
cc_1005 N_A_1555_410#_c_1396_n N_A_2516_368#_c_1784_n 7.76125e-19 $X=11.955
+ $Y=1.765 $X2=0 $Y2=0
cc_1006 N_A_1555_410#_c_1385_n N_A_2516_368#_c_1784_n 0.00894973f $X=12.845
+ $Y=1.515 $X2=0 $Y2=0
cc_1007 N_A_1555_410#_c_1386_n N_A_2516_368#_c_1784_n 0.00128211f $X=12.085
+ $Y=1.515 $X2=0 $Y2=0
cc_1008 N_A_1555_410#_c_1387_n N_A_2516_368#_c_1784_n 0.00716938f $X=12.935
+ $Y=1.765 $X2=0 $Y2=0
cc_1009 N_A_1555_410#_c_1384_n N_A_2516_368#_c_1778_n 0.00130472f $X=12.01
+ $Y=1.35 $X2=0 $Y2=0
cc_1010 N_A_1555_410#_c_1385_n N_A_2516_368#_c_1778_n 0.0176437f $X=12.845
+ $Y=1.515 $X2=0 $Y2=0
cc_1011 N_A_1555_410#_c_1387_n N_A_2516_368#_c_1778_n 0.00158462f $X=12.935
+ $Y=1.765 $X2=0 $Y2=0
cc_1012 N_A_1555_410#_c_1387_n N_A_2516_368#_c_1779_n 0.0103484f $X=12.935
+ $Y=1.765 $X2=0 $Y2=0
cc_1013 N_A_1555_410#_M1025_g N_A_2516_368#_c_1779_n 0.0107158f $X=13.015
+ $Y=0.69 $X2=0 $Y2=0
cc_1014 N_A_1555_410#_c_1401_n N_VPWR_M1004_d 0.00211046f $X=8.09 $Y=2.215 $X2=0
+ $Y2=0
cc_1015 N_A_1555_410#_c_1458_n N_VPWR_M1004_d 0.00398776f $X=8.255 $Y=2.715
+ $X2=0 $Y2=0
cc_1016 N_A_1555_410#_c_1408_n N_VPWR_M1004_d 0.00162375f $X=8.57 $Y=2.805 $X2=0
+ $Y2=0
cc_1017 N_A_1555_410#_c_1403_n N_VPWR_M1030_d 0.00848383f $X=10.06 $Y=2.715
+ $X2=0 $Y2=0
cc_1018 N_A_1555_410#_c_1406_n N_VPWR_M1021_d 0.00956316f $X=11.29 $Y=2.375
+ $X2=0 $Y2=0
cc_1019 N_A_1555_410#_c_1407_n N_VPWR_M1021_d 0.00540847f $X=11.375 $Y=2.29
+ $X2=0 $Y2=0
cc_1020 N_A_1555_410#_c_1395_n N_VPWR_c_1858_n 0.00856666f $X=11.505 $Y=1.765
+ $X2=0 $Y2=0
cc_1021 N_A_1555_410#_c_1396_n N_VPWR_c_1858_n 4.32634e-19 $X=11.955 $Y=1.765
+ $X2=0 $Y2=0
cc_1022 N_A_1555_410#_c_1406_n N_VPWR_c_1858_n 0.0227524f $X=11.29 $Y=2.375
+ $X2=0 $Y2=0
cc_1023 N_A_1555_410#_c_1395_n N_VPWR_c_1859_n 5.66383e-19 $X=11.505 $Y=1.765
+ $X2=0 $Y2=0
cc_1024 N_A_1555_410#_c_1396_n N_VPWR_c_1859_n 0.0149491f $X=11.955 $Y=1.765
+ $X2=0 $Y2=0
cc_1025 N_A_1555_410#_c_1386_n N_VPWR_c_1859_n 0.00893632f $X=12.085 $Y=1.515
+ $X2=0 $Y2=0
cc_1026 N_A_1555_410#_c_1387_n N_VPWR_c_1859_n 0.00394516f $X=12.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1027 N_A_1555_410#_c_1387_n N_VPWR_c_1860_n 0.00879434f $X=12.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1028 N_A_1555_410#_c_1392_n N_VPWR_c_1869_n 0.00478697f $X=7.865 $Y=2.465
+ $X2=0 $Y2=0
cc_1029 N_A_1555_410#_c_1402_n N_VPWR_c_1869_n 9.06413e-19 $X=8.09 $Y=2.215
+ $X2=0 $Y2=0
cc_1030 N_A_1555_410#_c_1458_n N_VPWR_c_1869_n 0.0197767f $X=8.255 $Y=2.715
+ $X2=0 $Y2=0
cc_1031 N_A_1555_410#_c_1408_n N_VPWR_c_1869_n 0.00619165f $X=8.57 $Y=2.805
+ $X2=0 $Y2=0
cc_1032 N_A_1555_410#_c_1409_n N_VPWR_c_1869_n 6.08883e-19 $X=8.9 $Y=2.805 $X2=0
+ $Y2=0
cc_1033 N_A_1555_410#_c_1392_n N_VPWR_c_1870_n 0.00446743f $X=7.865 $Y=2.465
+ $X2=0 $Y2=0
cc_1034 N_A_1555_410#_c_1458_n N_VPWR_c_1870_n 0.00140031f $X=8.255 $Y=2.715
+ $X2=0 $Y2=0
cc_1035 N_A_1555_410#_c_1403_n N_VPWR_c_1872_n 0.00283195f $X=10.06 $Y=2.715
+ $X2=0 $Y2=0
cc_1036 N_A_1555_410#_c_1408_n N_VPWR_c_1872_n 0.00532338f $X=8.57 $Y=2.805
+ $X2=0 $Y2=0
cc_1037 N_A_1555_410#_c_1409_n N_VPWR_c_1872_n 0.013942f $X=8.9 $Y=2.805 $X2=0
+ $Y2=0
cc_1038 N_A_1555_410#_c_1403_n N_VPWR_c_1873_n 0.0256793f $X=10.06 $Y=2.715
+ $X2=0 $Y2=0
cc_1039 N_A_1555_410#_c_1395_n N_VPWR_c_1874_n 0.00413917f $X=11.505 $Y=1.765
+ $X2=0 $Y2=0
cc_1040 N_A_1555_410#_c_1396_n N_VPWR_c_1874_n 0.00413917f $X=11.955 $Y=1.765
+ $X2=0 $Y2=0
cc_1041 N_A_1555_410#_c_1387_n N_VPWR_c_1875_n 0.00481995f $X=12.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1042 N_A_1555_410#_c_1403_n N_VPWR_c_1878_n 0.0244485f $X=10.06 $Y=2.715
+ $X2=0 $Y2=0
cc_1043 N_A_1555_410#_c_1409_n N_VPWR_c_1878_n 6.21521e-19 $X=8.9 $Y=2.805 $X2=0
+ $Y2=0
cc_1044 N_A_1555_410#_c_1392_n N_VPWR_c_1853_n 0.0086167f $X=7.865 $Y=2.465
+ $X2=0 $Y2=0
cc_1045 N_A_1555_410#_c_1395_n N_VPWR_c_1853_n 0.00817726f $X=11.505 $Y=1.765
+ $X2=0 $Y2=0
cc_1046 N_A_1555_410#_c_1396_n N_VPWR_c_1853_n 0.00817726f $X=11.955 $Y=1.765
+ $X2=0 $Y2=0
cc_1047 N_A_1555_410#_c_1387_n N_VPWR_c_1853_n 0.00508379f $X=12.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1048 N_A_1555_410#_c_1402_n N_VPWR_c_1853_n 3.4693e-19 $X=8.09 $Y=2.215 $X2=0
+ $Y2=0
cc_1049 N_A_1555_410#_c_1458_n N_VPWR_c_1853_n 0.00427608f $X=8.255 $Y=2.715
+ $X2=0 $Y2=0
cc_1050 N_A_1555_410#_c_1403_n N_VPWR_c_1853_n 0.0350508f $X=10.06 $Y=2.715
+ $X2=0 $Y2=0
cc_1051 N_A_1555_410#_c_1408_n N_VPWR_c_1853_n 0.00762788f $X=8.57 $Y=2.805
+ $X2=0 $Y2=0
cc_1052 N_A_1555_410#_c_1409_n N_VPWR_c_1853_n 0.0118463f $X=8.9 $Y=2.805 $X2=0
+ $Y2=0
cc_1053 N_A_1555_410#_c_1403_n A_1931_392# 0.0040234f $X=10.06 $Y=2.715
+ $X2=-0.19 $Y2=-0.245
cc_1054 N_A_1555_410#_c_1395_n N_Q_N_c_2157_n 0.00587498f $X=11.505 $Y=1.765
+ $X2=0 $Y2=0
cc_1055 N_A_1555_410#_c_1396_n N_Q_N_c_2157_n 0.00597227f $X=11.955 $Y=1.765
+ $X2=0 $Y2=0
cc_1056 N_A_1555_410#_c_1406_n N_Q_N_c_2157_n 0.0125099f $X=11.29 $Y=2.375 $X2=0
+ $Y2=0
cc_1057 N_A_1555_410#_c_1407_n N_Q_N_c_2157_n 0.0177267f $X=11.375 $Y=2.29 $X2=0
+ $Y2=0
cc_1058 N_A_1555_410#_c_1395_n N_Q_N_c_2155_n 5.50908e-19 $X=11.505 $Y=1.765
+ $X2=0 $Y2=0
cc_1059 N_A_1555_410#_c_1383_n N_Q_N_c_2155_n 0.00120476f $X=11.58 $Y=1.35 $X2=0
+ $Y2=0
cc_1060 N_A_1555_410#_c_1396_n N_Q_N_c_2155_n 0.00297846f $X=11.955 $Y=1.765
+ $X2=0 $Y2=0
cc_1061 N_A_1555_410#_c_1384_n N_Q_N_c_2155_n 0.00401782f $X=12.01 $Y=1.35 $X2=0
+ $Y2=0
cc_1062 N_A_1555_410#_c_1386_n N_Q_N_c_2155_n 0.0243888f $X=12.085 $Y=1.515
+ $X2=0 $Y2=0
cc_1063 N_A_1555_410#_c_1407_n N_Q_N_c_2155_n 0.00697757f $X=11.375 $Y=2.29
+ $X2=0 $Y2=0
cc_1064 N_A_1555_410#_c_1390_n N_Q_N_c_2155_n 0.0237053f $X=11.49 $Y=1.515 $X2=0
+ $Y2=0
cc_1065 N_A_1555_410#_c_1391_n N_Q_N_c_2155_n 0.0061611f $X=11.467 $Y=1.35 $X2=0
+ $Y2=0
cc_1066 N_A_1555_410#_c_1396_n N_Q_N_c_2171_n 0.00917834f $X=11.955 $Y=1.765
+ $X2=0 $Y2=0
cc_1067 N_A_1555_410#_c_1386_n N_Q_N_c_2171_n 0.00531555f $X=12.085 $Y=1.515
+ $X2=0 $Y2=0
cc_1068 N_A_1555_410#_c_1407_n N_Q_N_c_2171_n 0.0117299f $X=11.375 $Y=2.29 $X2=0
+ $Y2=0
cc_1069 N_A_1555_410#_c_1383_n Q_N 0.0124948f $X=11.58 $Y=1.35 $X2=0 $Y2=0
cc_1070 N_A_1555_410#_c_1384_n Q_N 0.00818893f $X=12.01 $Y=1.35 $X2=0 $Y2=0
cc_1071 N_A_1555_410#_c_1383_n Q_N 0.00223139f $X=11.58 $Y=1.35 $X2=0 $Y2=0
cc_1072 N_A_1555_410#_c_1384_n Q_N 0.00218568f $X=12.01 $Y=1.35 $X2=0 $Y2=0
cc_1073 N_A_1555_410#_c_1386_n Q_N 0.00211234f $X=12.085 $Y=1.515 $X2=0 $Y2=0
cc_1074 N_A_1555_410#_c_1390_n Q_N 0.00104314f $X=11.49 $Y=1.515 $X2=0 $Y2=0
cc_1075 N_A_1555_410#_M1025_g N_Q_c_2198_n 2.01998e-19 $X=13.015 $Y=0.69 $X2=0
+ $Y2=0
cc_1076 N_A_1555_410#_c_1389_n N_VGND_M1022_d 0.00794919f $X=11.29 $Y=0.755
+ $X2=0 $Y2=0
cc_1077 N_A_1555_410#_c_1391_n N_VGND_M1022_d 0.00727942f $X=11.467 $Y=1.35
+ $X2=0 $Y2=0
cc_1078 N_A_1555_410#_M1018_g N_VGND_c_2232_n 9.37761e-19 $X=8.515 $Y=0.9 $X2=0
+ $Y2=0
cc_1079 N_A_1555_410#_c_1384_n N_VGND_c_2233_n 0.00784853f $X=12.01 $Y=1.35
+ $X2=0 $Y2=0
cc_1080 N_A_1555_410#_c_1385_n N_VGND_c_2233_n 0.0111024f $X=12.845 $Y=1.515
+ $X2=0 $Y2=0
cc_1081 N_A_1555_410#_M1025_g N_VGND_c_2233_n 0.00412546f $X=13.015 $Y=0.69
+ $X2=0 $Y2=0
cc_1082 N_A_1555_410#_M1025_g N_VGND_c_2234_n 0.00367714f $X=13.015 $Y=0.69
+ $X2=0 $Y2=0
cc_1083 N_A_1555_410#_M1018_g N_VGND_c_2240_n 5.25761e-19 $X=8.515 $Y=0.9 $X2=0
+ $Y2=0
cc_1084 N_A_1555_410#_c_1383_n N_VGND_c_2241_n 0.00466874f $X=11.58 $Y=1.35
+ $X2=0 $Y2=0
cc_1085 N_A_1555_410#_c_1384_n N_VGND_c_2241_n 0.00445217f $X=12.01 $Y=1.35
+ $X2=0 $Y2=0
cc_1086 N_A_1555_410#_M1025_g N_VGND_c_2242_n 0.00461464f $X=13.015 $Y=0.69
+ $X2=0 $Y2=0
cc_1087 N_A_1555_410#_c_1389_n N_VGND_c_2248_n 0.00380543f $X=11.29 $Y=0.755
+ $X2=0 $Y2=0
cc_1088 N_A_1555_410#_c_1383_n N_VGND_c_2249_n 0.00463357f $X=11.58 $Y=1.35
+ $X2=0 $Y2=0
cc_1089 N_A_1555_410#_c_1389_n N_VGND_c_2249_n 0.0621166f $X=11.29 $Y=0.755
+ $X2=0 $Y2=0
cc_1090 N_A_1555_410#_c_1383_n N_VGND_c_2252_n 0.00505379f $X=11.58 $Y=1.35
+ $X2=0 $Y2=0
cc_1091 N_A_1555_410#_c_1384_n N_VGND_c_2252_n 0.00505379f $X=12.01 $Y=1.35
+ $X2=0 $Y2=0
cc_1092 N_A_1555_410#_M1025_g N_VGND_c_2252_n 0.00912712f $X=13.015 $Y=0.69
+ $X2=0 $Y2=0
cc_1093 N_A_1555_410#_c_1389_n N_VGND_c_2252_n 0.0109526f $X=11.29 $Y=0.755
+ $X2=0 $Y2=0
cc_1094 N_A_1555_410#_c_1389_n N_A_1832_74#_M1008_d 0.00776936f $X=11.29
+ $Y=0.755 $X2=0 $Y2=0
cc_1095 N_A_1555_410#_c_1389_n N_A_1832_74#_c_2411_n 0.0231054f $X=11.29
+ $Y=0.755 $X2=0 $Y2=0
cc_1096 N_A_1555_410#_M1019_d N_A_1832_74#_c_2412_n 0.00219516f $X=9.59 $Y=0.37
+ $X2=0 $Y2=0
cc_1097 N_A_1555_410#_c_1389_n N_A_1832_74#_c_2412_n 0.00570513f $X=11.29
+ $Y=0.755 $X2=0 $Y2=0
cc_1098 N_A_1555_410#_c_1430_n N_A_1832_74#_c_2412_n 0.0160573f $X=9.935
+ $Y=0.717 $X2=0 $Y2=0
cc_1099 N_A_1335_112#_c_1606_n N_RESET_B_c_1744_n 0.00455386f $X=10 $Y=1.885
+ $X2=-0.19 $Y2=-0.245
cc_1100 N_A_1335_112#_c_1659_n N_VPWR_M1030_d 0.0168547f $X=9.72 $Y=2.375 $X2=0
+ $Y2=0
cc_1101 N_A_1335_112#_c_1611_n N_VPWR_c_1857_n 0.00959573f $X=7.13 $Y=2.815
+ $X2=0 $Y2=0
cc_1102 N_A_1335_112#_c_1611_n N_VPWR_c_1869_n 3.31509e-19 $X=7.13 $Y=2.815
+ $X2=0 $Y2=0
cc_1103 N_A_1335_112#_c_1611_n N_VPWR_c_1870_n 0.0214821f $X=7.13 $Y=2.815 $X2=0
+ $Y2=0
cc_1104 N_A_1335_112#_c_1606_n N_VPWR_c_1873_n 0.00361118f $X=10 $Y=1.885 $X2=0
+ $Y2=0
cc_1105 N_A_1335_112#_c_1606_n N_VPWR_c_1853_n 0.0056474f $X=10 $Y=1.885 $X2=0
+ $Y2=0
cc_1106 N_A_1335_112#_c_1611_n N_VPWR_c_1853_n 0.0175508f $X=7.13 $Y=2.815 $X2=0
+ $Y2=0
cc_1107 N_A_1335_112#_c_1659_n A_1931_392# 0.0022665f $X=9.72 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_1108 N_A_1335_112#_c_1618_n A_1931_392# 0.00434173f $X=9.805 $Y=2.29
+ $X2=-0.19 $Y2=-0.245
cc_1109 N_A_1335_112#_M1008_g N_VGND_c_2248_n 0.00278271f $X=9.985 $Y=0.74 $X2=0
+ $Y2=0
cc_1110 N_A_1335_112#_M1008_g N_VGND_c_2249_n 0.00113361f $X=9.985 $Y=0.74 $X2=0
+ $Y2=0
cc_1111 N_A_1335_112#_M1008_g N_VGND_c_2252_n 0.00358885f $X=9.985 $Y=0.74 $X2=0
+ $Y2=0
cc_1112 N_A_1335_112#_c_1607_n A_1640_138# 0.00278314f $X=8.105 $Y=0.845
+ $X2=-0.19 $Y2=-0.245
cc_1113 N_A_1335_112#_c_1608_n A_1640_138# 8.25348e-19 $X=8.19 $Y=1.72 $X2=-0.19
+ $Y2=-0.245
cc_1114 N_A_1335_112#_M1008_g N_A_1832_74#_c_2412_n 0.0112967f $X=9.985 $Y=0.74
+ $X2=0 $Y2=0
cc_1115 N_RESET_B_c_1744_n N_VPWR_c_1873_n 0.00314304f $X=10.98 $Y=1.765 $X2=0
+ $Y2=0
cc_1116 N_RESET_B_c_1744_n N_VPWR_c_1853_n 0.00411481f $X=10.98 $Y=1.765 $X2=0
+ $Y2=0
cc_1117 N_RESET_B_c_1745_n N_VGND_c_2249_n 0.00109048f $X=11.04 $Y=1.35 $X2=0
+ $Y2=0
cc_1118 N_A_2516_368#_c_1783_n N_VPWR_c_1859_n 0.0497747f $X=12.71 $Y=2.695
+ $X2=0 $Y2=0
cc_1119 N_A_2516_368#_c_1780_n N_VPWR_c_1860_n 0.00911654f $X=13.455 $Y=1.765
+ $X2=0 $Y2=0
cc_1120 N_A_2516_368#_c_1782_n N_VPWR_c_1860_n 0.0370638f $X=12.71 $Y=1.985
+ $X2=0 $Y2=0
cc_1121 N_A_2516_368#_c_1777_n N_VPWR_c_1860_n 0.0182992f $X=13.53 $Y=1.435
+ $X2=0 $Y2=0
cc_1122 N_A_2516_368#_c_1781_n N_VPWR_c_1862_n 0.0106074f $X=13.905 $Y=1.765
+ $X2=0 $Y2=0
cc_1123 N_A_2516_368#_c_1783_n N_VPWR_c_1875_n 0.0097982f $X=12.71 $Y=2.695
+ $X2=0 $Y2=0
cc_1124 N_A_2516_368#_c_1780_n N_VPWR_c_1876_n 0.00445602f $X=13.455 $Y=1.765
+ $X2=0 $Y2=0
cc_1125 N_A_2516_368#_c_1781_n N_VPWR_c_1876_n 0.00445602f $X=13.905 $Y=1.765
+ $X2=0 $Y2=0
cc_1126 N_A_2516_368#_c_1780_n N_VPWR_c_1853_n 0.00862391f $X=13.455 $Y=1.765
+ $X2=0 $Y2=0
cc_1127 N_A_2516_368#_c_1781_n N_VPWR_c_1853_n 0.0086105f $X=13.905 $Y=1.765
+ $X2=0 $Y2=0
cc_1128 N_A_2516_368#_c_1783_n N_VPWR_c_1853_n 0.0111907f $X=12.71 $Y=2.695
+ $X2=0 $Y2=0
cc_1129 N_A_2516_368#_c_1782_n N_Q_N_c_2155_n 9.27117e-19 $X=12.71 $Y=1.985
+ $X2=0 $Y2=0
cc_1130 N_A_2516_368#_c_1776_n N_Q_N_c_2155_n 2.5156e-19 $X=12.8 $Y=0.515 $X2=0
+ $Y2=0
cc_1131 N_A_2516_368#_c_1784_n N_Q_N_c_2155_n 0.00551167f $X=12.71 $Y=1.82 $X2=0
+ $Y2=0
cc_1132 N_A_2516_368#_c_1778_n N_Q_N_c_2155_n 0.00854201f $X=12.76 $Y=1.435
+ $X2=0 $Y2=0
cc_1133 N_A_2516_368#_c_1782_n N_Q_N_c_2171_n 0.00542337f $X=12.71 $Y=1.985
+ $X2=0 $Y2=0
cc_1134 N_A_2516_368#_M1006_g N_Q_c_2193_n 0.00585678f $X=13.49 $Y=0.74 $X2=0
+ $Y2=0
cc_1135 N_A_2516_368#_M1026_g N_Q_c_2193_n 2.74318e-19 $X=13.92 $Y=0.74 $X2=0
+ $Y2=0
cc_1136 N_A_2516_368#_M1006_g N_Q_c_2194_n 9.98187e-19 $X=13.49 $Y=0.74 $X2=0
+ $Y2=0
cc_1137 N_A_2516_368#_c_1781_n N_Q_c_2194_n 4.02332e-19 $X=13.905 $Y=1.765 $X2=0
+ $Y2=0
cc_1138 N_A_2516_368#_M1026_g N_Q_c_2194_n 0.00716185f $X=13.92 $Y=0.74 $X2=0
+ $Y2=0
cc_1139 N_A_2516_368#_c_1777_n N_Q_c_2194_n 0.0249855f $X=13.53 $Y=1.435 $X2=0
+ $Y2=0
cc_1140 N_A_2516_368#_c_1779_n N_Q_c_2194_n 0.0211802f $X=13.905 $Y=1.517 $X2=0
+ $Y2=0
cc_1141 N_A_2516_368#_c_1780_n N_Q_c_2196_n 0.00325284f $X=13.455 $Y=1.765 $X2=0
+ $Y2=0
cc_1142 N_A_2516_368#_c_1781_n N_Q_c_2196_n 0.0132092f $X=13.905 $Y=1.765 $X2=0
+ $Y2=0
cc_1143 N_A_2516_368#_c_1777_n N_Q_c_2196_n 0.0134719f $X=13.53 $Y=1.435 $X2=0
+ $Y2=0
cc_1144 N_A_2516_368#_c_1784_n N_Q_c_2196_n 0.00122489f $X=12.71 $Y=1.82 $X2=0
+ $Y2=0
cc_1145 N_A_2516_368#_c_1779_n N_Q_c_2196_n 0.00873201f $X=13.905 $Y=1.517 $X2=0
+ $Y2=0
cc_1146 N_A_2516_368#_M1006_g N_Q_c_2198_n 0.00346861f $X=13.49 $Y=0.74 $X2=0
+ $Y2=0
cc_1147 N_A_2516_368#_M1026_g N_Q_c_2198_n 0.0114931f $X=13.92 $Y=0.74 $X2=0
+ $Y2=0
cc_1148 N_A_2516_368#_c_1776_n N_Q_c_2198_n 0.00138446f $X=12.8 $Y=0.515 $X2=0
+ $Y2=0
cc_1149 N_A_2516_368#_c_1777_n N_Q_c_2198_n 0.00948769f $X=13.53 $Y=1.435 $X2=0
+ $Y2=0
cc_1150 N_A_2516_368#_c_1779_n N_Q_c_2198_n 0.00258535f $X=13.905 $Y=1.517 $X2=0
+ $Y2=0
cc_1151 N_A_2516_368#_c_1780_n Q 0.0117465f $X=13.455 $Y=1.765 $X2=0 $Y2=0
cc_1152 N_A_2516_368#_c_1781_n Q 0.0176348f $X=13.905 $Y=1.765 $X2=0 $Y2=0
cc_1153 N_A_2516_368#_c_1776_n N_VGND_c_2233_n 0.0588254f $X=12.8 $Y=0.515 $X2=0
+ $Y2=0
cc_1154 N_A_2516_368#_M1006_g N_VGND_c_2234_n 0.00170242f $X=13.49 $Y=0.74 $X2=0
+ $Y2=0
cc_1155 N_A_2516_368#_c_1776_n N_VGND_c_2234_n 0.00401787f $X=12.8 $Y=0.515
+ $X2=0 $Y2=0
cc_1156 N_A_2516_368#_c_1777_n N_VGND_c_2234_n 0.0193405f $X=13.53 $Y=1.435
+ $X2=0 $Y2=0
cc_1157 N_A_2516_368#_M1006_g N_VGND_c_2236_n 4.37711e-19 $X=13.49 $Y=0.74 $X2=0
+ $Y2=0
cc_1158 N_A_2516_368#_M1026_g N_VGND_c_2236_n 0.00879435f $X=13.92 $Y=0.74 $X2=0
+ $Y2=0
cc_1159 N_A_2516_368#_c_1776_n N_VGND_c_2242_n 0.011066f $X=12.8 $Y=0.515 $X2=0
+ $Y2=0
cc_1160 N_A_2516_368#_M1006_g N_VGND_c_2243_n 0.00434272f $X=13.49 $Y=0.74 $X2=0
+ $Y2=0
cc_1161 N_A_2516_368#_M1026_g N_VGND_c_2243_n 0.00383152f $X=13.92 $Y=0.74 $X2=0
+ $Y2=0
cc_1162 N_A_2516_368#_M1006_g N_VGND_c_2252_n 0.00815946f $X=13.49 $Y=0.74 $X2=0
+ $Y2=0
cc_1163 N_A_2516_368#_M1026_g N_VGND_c_2252_n 0.00386058f $X=13.92 $Y=0.74 $X2=0
+ $Y2=0
cc_1164 N_A_2516_368#_c_1776_n N_VGND_c_2252_n 0.00915947f $X=12.8 $Y=0.515
+ $X2=0 $Y2=0
cc_1165 N_VPWR_c_1858_n N_Q_N_c_2157_n 0.0228252f $X=11.28 $Y=2.805 $X2=0 $Y2=0
cc_1166 N_VPWR_c_1859_n N_Q_N_c_2157_n 0.0514854f $X=12.18 $Y=2.355 $X2=0 $Y2=0
cc_1167 N_VPWR_c_1874_n N_Q_N_c_2157_n 0.00749631f $X=12.015 $Y=3.33 $X2=0 $Y2=0
cc_1168 N_VPWR_c_1853_n N_Q_N_c_2157_n 0.0062048f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1169 N_VPWR_c_1860_n N_Q_c_2196_n 0.00832528f $X=13.23 $Y=1.985 $X2=0 $Y2=0
cc_1170 N_VPWR_c_1860_n Q 0.0697627f $X=13.23 $Y=1.985 $X2=0 $Y2=0
cc_1171 N_VPWR_c_1862_n Q 0.058364f $X=14.13 $Y=2.275 $X2=0 $Y2=0
cc_1172 N_VPWR_c_1876_n Q 0.014552f $X=14.045 $Y=3.33 $X2=0 $Y2=0
cc_1173 N_VPWR_c_1853_n Q 0.0119791f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1174 N_A_311_119#_c_2045_n N_VGND_M1015_d 0.0086414f $X=2.61 $Y=0.925 $X2=0
+ $Y2=0
cc_1175 N_A_311_119#_c_2045_n N_VGND_c_2230_n 0.0311142f $X=2.61 $Y=0.925 $X2=0
+ $Y2=0
cc_1176 N_A_311_119#_c_2027_n N_VGND_c_2230_n 0.0156421f $X=2.695 $Y=0.84 $X2=0
+ $Y2=0
cc_1177 N_A_311_119#_c_2028_n N_VGND_c_2230_n 0.015234f $X=2.78 $Y=0.34 $X2=0
+ $Y2=0
cc_1178 N_A_311_119#_c_2033_n N_VGND_c_2230_n 0.00404325f $X=1.7 $Y=0.79 $X2=0
+ $Y2=0
cc_1179 N_A_311_119#_c_2033_n N_VGND_c_2238_n 0.00559729f $X=1.7 $Y=0.79 $X2=0
+ $Y2=0
cc_1180 N_A_311_119#_c_2028_n N_VGND_c_2239_n 0.0115893f $X=2.78 $Y=0.34 $X2=0
+ $Y2=0
cc_1181 N_A_311_119#_c_2029_n N_VGND_c_2239_n 0.0115893f $X=4.055 $Y=0.435 $X2=0
+ $Y2=0
cc_1182 N_A_311_119#_c_2034_n N_VGND_c_2239_n 0.0835348f $X=3.49 $Y=0.435 $X2=0
+ $Y2=0
cc_1183 N_A_311_119#_c_2045_n N_VGND_c_2252_n 0.0112675f $X=2.61 $Y=0.925 $X2=0
+ $Y2=0
cc_1184 N_A_311_119#_c_2028_n N_VGND_c_2252_n 0.00583135f $X=2.78 $Y=0.34 $X2=0
+ $Y2=0
cc_1185 N_A_311_119#_c_2029_n N_VGND_c_2252_n 0.00583135f $X=4.055 $Y=0.435
+ $X2=0 $Y2=0
cc_1186 N_A_311_119#_c_2033_n N_VGND_c_2252_n 0.00680542f $X=1.7 $Y=0.79 $X2=0
+ $Y2=0
cc_1187 N_A_311_119#_c_2034_n N_VGND_c_2252_n 0.0430568f $X=3.49 $Y=0.435 $X2=0
+ $Y2=0
cc_1188 N_A_311_119#_c_2045_n A_529_119# 0.00287182f $X=2.61 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_1189 N_A_311_119#_c_2027_n A_529_119# 0.00211902f $X=2.695 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_1190 N_A_311_119#_c_2035_n N_A_867_125#_M1035_s 0.00340675f $X=4.35 $Y=1.21
+ $X2=-0.19 $Y2=-0.245
cc_1191 N_A_311_119#_c_2029_n N_A_867_125#_c_2376_n 0.0151648f $X=4.055 $Y=0.435
+ $X2=0 $Y2=0
cc_1192 N_A_311_119#_c_2031_n N_A_867_125#_c_2376_n 0.0251238f $X=4.14 $Y=1.125
+ $X2=0 $Y2=0
cc_1193 N_A_311_119#_c_2035_n N_A_867_125#_c_2376_n 0.00291702f $X=4.35 $Y=1.21
+ $X2=0 $Y2=0
cc_1194 N_A_311_119#_c_2029_n N_A_867_125#_c_2378_n 0.0159286f $X=4.055 $Y=0.435
+ $X2=0 $Y2=0
cc_1195 Q_N N_VGND_c_2233_n 0.0623798f $X=11.675 $Y=0.47 $X2=0 $Y2=0
cc_1196 Q_N N_VGND_c_2241_n 0.0113495f $X=11.675 $Y=0.47 $X2=0 $Y2=0
cc_1197 Q_N N_VGND_c_2249_n 0.00478905f $X=11.675 $Y=0.47 $X2=0 $Y2=0
cc_1198 Q_N N_VGND_c_2252_n 0.0122366f $X=11.675 $Y=0.47 $X2=0 $Y2=0
cc_1199 N_Q_c_2193_n N_VGND_c_2234_n 0.0188572f $X=13.705 $Y=0.515 $X2=0 $Y2=0
cc_1200 N_Q_c_2193_n N_VGND_c_2236_n 0.0131449f $X=13.705 $Y=0.515 $X2=0 $Y2=0
cc_1201 N_Q_c_2198_n N_VGND_c_2236_n 0.0017952f $X=13.95 $Y=0.975 $X2=0 $Y2=0
cc_1202 N_Q_c_2193_n N_VGND_c_2243_n 0.0111905f $X=13.705 $Y=0.515 $X2=0 $Y2=0
cc_1203 N_Q_c_2193_n N_VGND_c_2252_n 0.00931592f $X=13.705 $Y=0.515 $X2=0 $Y2=0
cc_1204 N_Q_c_2198_n N_VGND_c_2252_n 0.00534972f $X=13.95 $Y=0.975 $X2=0 $Y2=0
cc_1205 N_VGND_c_2231_n N_A_867_125#_c_2377_n 0.0150385f $X=5.91 $Y=0.86 $X2=0
+ $Y2=0
cc_1206 N_VGND_c_2239_n N_A_867_125#_c_2377_n 0.063402f $X=5.745 $Y=0 $X2=0
+ $Y2=0
cc_1207 N_VGND_c_2252_n N_A_867_125#_c_2377_n 0.0341454f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1208 N_VGND_c_2239_n N_A_867_125#_c_2378_n 0.0114699f $X=5.745 $Y=0 $X2=0
+ $Y2=0
cc_1209 N_VGND_c_2252_n N_A_867_125#_c_2378_n 0.00590238f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1210 N_VGND_c_2231_n N_A_867_125#_c_2379_n 0.0302085f $X=5.91 $Y=0.86 $X2=0
+ $Y2=0
cc_1211 N_VGND_c_2232_n N_A_1832_74#_c_2410_n 0.010974f $X=8.87 $Y=0.595 $X2=0
+ $Y2=0
cc_1212 N_VGND_c_2248_n N_A_1832_74#_c_2410_n 0.0176346f $X=10.665 $Y=0.207
+ $X2=0 $Y2=0
cc_1213 N_VGND_c_2252_n N_A_1832_74#_c_2410_n 0.00956728f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1214 N_VGND_c_2249_n N_A_1832_74#_c_2411_n 0.0183835f $X=11.45 $Y=0.207 $X2=0
+ $Y2=0
cc_1215 N_VGND_c_2248_n N_A_1832_74#_c_2412_n 0.0675786f $X=10.665 $Y=0.207
+ $X2=0 $Y2=0
cc_1216 N_VGND_c_2252_n N_A_1832_74#_c_2412_n 0.0383916f $X=14.16 $Y=0 $X2=0
+ $Y2=0
