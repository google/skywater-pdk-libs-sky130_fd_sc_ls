* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__buf_4 A VGND VNB VPB VPWR X
M1000 VGND a_86_260# X VNB nshort w=740000u l=150000u
+  ad=1.1063e+12p pd=7.43e+06u as=4.144e+11p ps=4.08e+06u
M1001 a_86_260# A VPWR VPB phighvt w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=1.3202e+12p ps=1.095e+07u
M1002 VPWR a_86_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.72e+11p ps=5.68e+06u
M1003 X a_86_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_86_260# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_86_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_86_260# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_86_260# A VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 X a_86_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_86_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_86_260# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
