* NGSPICE file created from sky130_fd_sc_ls__nor4_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nor4_1 A B C D VGND VNB VPB VPWR Y
M1000 Y A VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=8.7975e+11p ps=6.9e+06u
M1001 Y D a_342_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=4.704e+11p ps=3.08e+06u
M1002 a_228_368# B a_144_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=4.704e+11p pd=3.08e+06u as=3.024e+11p ps=2.78e+06u
M1003 a_342_368# C a_228_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND B Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y C VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND D Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_144_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
.ends

