* File: sky130_fd_sc_ls__and2_1.spice
* Created: Fri Aug 28 13:02:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__and2_1.pex.spice"
.subckt sky130_fd_sc_ls__and2_1  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 A_143_136# N_A_M1002_g N_A_56_136#_M1002_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1376 AS=0.1824 PD=1.14 PS=1.85 NRD=30 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1001_d N_B_M1001_g A_143_136# VNB NSHORT L=0.15 W=0.64
+ AD=0.144093 AS=0.1376 PD=1.08522 PS=1.14 NRD=14.988 NRS=30 M=1 R=4.26667
+ SA=75000.7 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1005 N_X_M1005_d N_A_56_136#_M1005_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.166607 PD=2.05 PS=1.25478 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_56_136#_M1004_d N_A_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.147 AS=0.252 PD=1.19 PS=2.28 NRD=14.0658 NRS=3.5066 M=1 R=5.6 SA=75000.2
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_B_M1000_g N_A_56_136#_M1004_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1704 AS=0.147 PD=1.29 PS=1.19 NRD=22.261 NRS=2.3443 M=1 R=5.6 SA=75000.7
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1003 N_X_M1003_d N_A_56_136#_M1003_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.2272 PD=2.83 PS=1.72 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001 SB=75000.2 A=0.168 P=2.54 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_ls__and2_1.pxi.spice"
*
.ends
*
*
