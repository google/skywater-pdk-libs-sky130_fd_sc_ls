* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 a_89_270# C1 VGND VNB nshort w=640000u l=150000u
+  ad=3.488e+11p pd=3.65e+06u as=5.289e+11p ps=4.33e+06u
M1001 a_264_120# A3 VGND VNB nshort w=640000u l=150000u
+  ad=2.10625e+11p pd=1.96e+06u as=0p ps=0u
M1002 VPWR A2 a_258_392# VPB phighvt w=1e+06u l=150000u
+  ad=9.518e+11p pd=6.08e+06u as=6e+11p ps=5.2e+06u
M1003 VGND a_89_270# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=1.961e+11p ps=2.01e+06u
M1004 a_89_270# A1 a_359_123# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.048e+11p ps=1.92e+06u
M1005 a_258_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_546_392# B1 a_258_392# VPB phighvt w=1e+06u l=150000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1007 a_89_270# C1 a_546_392# VPB phighvt w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1008 a_359_123# A2 a_264_120# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_258_392# A3 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_89_270# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.08e+11p ps=2.79e+06u
M1011 VGND B1 a_89_270# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
