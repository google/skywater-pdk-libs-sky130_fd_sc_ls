* File: sky130_fd_sc_ls__nor3_2.spice
* Created: Fri Aug 28 13:38:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nor3_2.pex.spice"
.subckt sky130_fd_sc_ls__nor3_2  VNB VPB C B A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_C_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.32745 AS=0.2109 PD=1.625 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1008_d N_B_M1008_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.74 AD=0.1295
+ AS=0.32745 PD=1.09 PS=1.625 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_Y_M1008_d VNB NSHORT L=0.15 W=0.74 AD=0.2627
+ AS=0.1295 PD=2.19 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.7 SB=75000.3
+ A=0.111 P=1.78 MULT=1
MM1003 N_A_27_368#_M1003_d N_C_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.2 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1004 N_A_27_368#_M1004_d N_C_M1004_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1002 N_A_27_368#_M1004_d N_B_M1002_g N_A_306_368#_M1002_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.1848 PD=1.42 PS=1.45 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1000 N_A_306_368#_M1002_s N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.1848 AS=0.1792 PD=1.45 PS=1.44 NRD=7.0329 NRS=5.2599 M=1 R=7.46667
+ SA=75001.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1001 N_A_306_368#_M1001_d N_A_M1001_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.1792 PD=1.42 PS=1.44 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1005 N_A_27_368#_M1005_d N_B_M1005_g N_A_306_368#_M1001_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX9_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ls__nor3_2.pxi.spice"
*
.ends
*
*
