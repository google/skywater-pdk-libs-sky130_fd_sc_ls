* File: sky130_fd_sc_ls__or4_1.spice
* Created: Wed Sep  2 11:25:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__or4_1.pex.spice"
.subckt sky130_fd_sc_ls__or4_1  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1002 N_A_44_392#_M1002_d N_D_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.19525 PD=0.83 PS=1.81 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.3
+ SB=75002.5 A=0.0825 P=1.4 MULT=1
MM1001 N_VGND_M1001_d N_C_M1001_g N_A_44_392#_M1002_d VNB NSHORT L=0.15 W=0.55
+ AD=0.1674 AS=0.077 PD=1.165 PS=0.83 NRD=32.724 NRS=0 M=1 R=3.66667 SA=75000.7
+ SB=75002 A=0.0825 P=1.4 MULT=1
MM1004 N_A_44_392#_M1004_d N_B_M1004_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.55
+ AD=0.121 AS=0.1674 PD=0.99 PS=1.165 NRD=17.448 NRS=33.816 M=1 R=3.66667
+ SA=75001.4 SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_44_392#_M1004_d VNB NSHORT L=0.15 W=0.55
+ AD=0.107506 AS=0.121 PD=0.937984 PS=0.99 NRD=17.448 NRS=17.448 M=1 R=3.66667
+ SA=75002 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1006 N_X_M1006_d N_A_44_392#_M1006_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.144644 PD=2.05 PS=1.26202 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 A_133_392# N_D_M1000_g N_A_44_392#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.5 A=0.15 P=2.3 MULT=1
MM1007 A_217_392# N_C_M1007_g A_133_392# VPB PHIGHVT L=0.15 W=1 AD=0.21 AS=0.135
+ PD=1.42 PS=1.27 NRD=30.5153 NRS=15.7403 M=1 R=6.66667 SA=75000.6 SB=75002
+ A=0.15 P=2.3 MULT=1
MM1009 A_331_392# N_B_M1009_g A_217_392# VPB PHIGHVT L=0.15 W=1 AD=0.21 AS=0.21
+ PD=1.42 PS=1.42 NRD=30.5153 NRS=30.5153 M=1 R=6.66667 SA=75001.2 SB=75001.5
+ A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g A_331_392# VPB PHIGHVT L=0.15 W=1 AD=0.269717
+ AS=0.21 PD=1.56604 PS=1.42 NRD=1.9503 NRS=30.5153 M=1 R=6.66667 SA=75001.8
+ SB=75000.9 A=0.15 P=2.3 MULT=1
MM1008 N_X_M1008_d N_A_44_392#_M1008_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.302083 PD=2.83 PS=1.75396 NRD=1.7533 NRS=43.9704 M=1 R=7.46667
+ SA=75002.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ls__or4_1.pxi.spice"
*
.ends
*
*
