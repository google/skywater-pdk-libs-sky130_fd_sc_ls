* File: sky130_fd_sc_ls__xor2_4.pxi.spice
* Created: Fri Aug 28 14:10:21 2020
* 
x_PM_SKY130_FD_SC_LS__XOR2_4%A N_A_c_161_n N_A_M1021_g N_A_M1000_g N_A_c_162_n
+ N_A_M1023_g N_A_M1016_g N_A_c_163_n N_A_M1005_g N_A_M1009_g N_A_c_164_n
+ N_A_M1013_g N_A_M1010_g N_A_M1020_g N_A_c_165_n N_A_M1025_g N_A_c_150_n
+ N_A_c_151_n N_A_c_168_n N_A_M1028_g N_A_M1024_g N_A_c_153_n N_A_c_154_n
+ N_A_c_322_p N_A_c_155_n N_A_c_185_p N_A_c_177_p N_A_c_180_p N_A_c_202_p
+ N_A_c_209_p N_A_c_156_n N_A_c_205_p N_A_c_178_p A A A A N_A_c_158_n
+ N_A_c_159_n N_A_c_160_n PM_SKY130_FD_SC_LS__XOR2_4%A
x_PM_SKY130_FD_SC_LS__XOR2_4%B N_B_c_388_n N_B_M1001_g N_B_M1017_g N_B_c_389_n
+ N_B_M1006_g N_B_M1026_g N_B_c_375_n N_B_c_376_n N_B_M1003_g N_B_c_391_n
+ N_B_M1002_g N_B_c_378_n N_B_c_379_n N_B_M1007_g N_B_c_392_n N_B_M1011_g
+ N_B_c_393_n N_B_M1015_g N_B_M1014_g N_B_c_382_n N_B_M1019_g N_B_c_395_n
+ N_B_M1022_g N_B_c_384_n N_B_c_385_n N_B_c_397_n N_B_c_398_n N_B_c_413_n
+ N_B_c_386_n N_B_c_399_n N_B_c_428_n B B B B B N_B_c_387_n B
+ PM_SKY130_FD_SC_LS__XOR2_4%B
x_PM_SKY130_FD_SC_LS__XOR2_4%A_160_98# N_A_160_98#_M1000_d N_A_160_98#_M1017_d
+ N_A_160_98#_M1001_d N_A_160_98#_c_578_n N_A_160_98#_M1008_g
+ N_A_160_98#_c_587_n N_A_160_98#_M1004_g N_A_160_98#_c_588_n
+ N_A_160_98#_M1012_g N_A_160_98#_c_579_n N_A_160_98#_M1027_g
+ N_A_160_98#_c_589_n N_A_160_98#_M1018_g N_A_160_98#_c_580_n
+ N_A_160_98#_c_581_n N_A_160_98#_c_592_n N_A_160_98#_M1029_g
+ N_A_160_98#_c_582_n N_A_160_98#_c_613_n N_A_160_98#_c_583_n
+ N_A_160_98#_c_621_n N_A_160_98#_c_584_n N_A_160_98#_c_585_n
+ N_A_160_98#_c_624_n N_A_160_98#_c_586_n N_A_160_98#_c_633_n
+ PM_SKY130_FD_SC_LS__XOR2_4%A_160_98#
x_PM_SKY130_FD_SC_LS__XOR2_4%A_36_392# N_A_36_392#_M1021_d N_A_36_392#_M1023_d
+ N_A_36_392#_M1006_s N_A_36_392#_c_718_n N_A_36_392#_c_719_n
+ N_A_36_392#_c_720_n N_A_36_392#_c_734_n N_A_36_392#_c_721_n
+ N_A_36_392#_c_722_n N_A_36_392#_c_723_n PM_SKY130_FD_SC_LS__XOR2_4%A_36_392#
x_PM_SKY130_FD_SC_LS__XOR2_4%VPWR N_VPWR_M1021_s N_VPWR_M1005_s N_VPWR_M1025_s
+ N_VPWR_M1002_d N_VPWR_M1015_d N_VPWR_c_765_n N_VPWR_c_766_n N_VPWR_c_767_n
+ VPWR N_VPWR_c_768_n N_VPWR_c_769_n N_VPWR_c_770_n N_VPWR_c_771_n
+ N_VPWR_c_772_n N_VPWR_c_764_n N_VPWR_c_774_n N_VPWR_c_775_n N_VPWR_c_776_n
+ N_VPWR_c_777_n N_VPWR_c_778_n PM_SKY130_FD_SC_LS__XOR2_4%VPWR
x_PM_SKY130_FD_SC_LS__XOR2_4%A_514_368# N_A_514_368#_M1004_d
+ N_A_514_368#_M1012_d N_A_514_368#_M1029_d N_A_514_368#_M1013_d
+ N_A_514_368#_M1028_d N_A_514_368#_M1011_s N_A_514_368#_M1022_s
+ N_A_514_368#_c_881_n N_A_514_368#_c_882_n N_A_514_368#_c_883_n
+ N_A_514_368#_c_990_p N_A_514_368#_c_884_n N_A_514_368#_c_891_n
+ N_A_514_368#_c_975_p N_A_514_368#_c_885_n N_A_514_368#_c_911_n
+ N_A_514_368#_c_913_n N_A_514_368#_c_886_n N_A_514_368#_c_887_n
+ N_A_514_368#_c_896_n N_A_514_368#_c_888_n N_A_514_368#_c_889_n
+ N_A_514_368#_c_890_n PM_SKY130_FD_SC_LS__XOR2_4%A_514_368#
x_PM_SKY130_FD_SC_LS__XOR2_4%X N_X_M1008_s N_X_M1003_d N_X_M1014_d N_X_M1004_s
+ N_X_M1018_s N_X_c_998_n N_X_c_999_n N_X_c_1017_n N_X_c_1000_n N_X_c_1001_n
+ N_X_c_1034_n N_X_c_1008_n N_X_c_1037_n N_X_c_1040_n N_X_c_1002_n N_X_c_1164_p
+ N_X_c_1003_n N_X_c_1004_n N_X_c_1076_n N_X_c_1005_n N_X_c_1006_n N_X_c_1007_n
+ X N_X_c_1083_n N_X_c_1044_n PM_SKY130_FD_SC_LS__XOR2_4%X
x_PM_SKY130_FD_SC_LS__XOR2_4%VGND N_VGND_M1000_s N_VGND_M1016_s N_VGND_M1026_s
+ N_VGND_M1027_d N_VGND_M1009_d N_VGND_M1020_d N_VGND_c_1170_n N_VGND_c_1171_n
+ N_VGND_c_1172_n N_VGND_c_1173_n N_VGND_c_1174_n N_VGND_c_1175_n
+ N_VGND_c_1176_n N_VGND_c_1177_n N_VGND_c_1178_n N_VGND_c_1179_n VGND
+ N_VGND_c_1180_n N_VGND_c_1181_n N_VGND_c_1182_n N_VGND_c_1183_n
+ N_VGND_c_1184_n N_VGND_c_1185_n N_VGND_c_1186_n N_VGND_c_1187_n
+ PM_SKY130_FD_SC_LS__XOR2_4%VGND
x_PM_SKY130_FD_SC_LS__XOR2_4%A_877_74# N_A_877_74#_M1009_s N_A_877_74#_M1010_s
+ N_A_877_74#_M1024_s N_A_877_74#_M1007_s N_A_877_74#_M1019_s
+ N_A_877_74#_c_1299_n N_A_877_74#_c_1301_n N_A_877_74#_c_1292_n
+ N_A_877_74#_c_1293_n N_A_877_74#_c_1316_n N_A_877_74#_c_1294_n
+ N_A_877_74#_c_1295_n N_A_877_74#_c_1296_n N_A_877_74#_c_1306_n
+ N_A_877_74#_c_1297_n N_A_877_74#_c_1298_n PM_SKY130_FD_SC_LS__XOR2_4%A_877_74#
cc_1 VNB N_A_M1000_g 0.0234074f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.86
cc_2 VNB N_A_M1016_g 0.0225154f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.86
cc_3 VNB N_A_M1009_g 0.0328409f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=0.74
cc_4 VNB N_A_M1010_g 0.025165f $X=-0.19 $Y=-0.245 $X2=5.335 $Y2=0.74
cc_5 VNB N_A_M1020_g 0.025165f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=0.74
cc_6 VNB N_A_c_150_n 0.0398611f $X=-0.19 $Y=-0.245 $X2=6.255 $Y2=1.485
cc_7 VNB N_A_c_151_n 0.0238469f $X=-0.19 $Y=-0.245 $X2=5.855 $Y2=1.485
cc_8 VNB N_A_M1024_g 0.025058f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=0.74
cc_9 VNB N_A_c_153_n 0.0153059f $X=-0.19 $Y=-0.245 $X2=4.605 $Y2=1.35
cc_10 VNB N_A_c_154_n 0.00598948f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.42
cc_11 VNB N_A_c_155_n 0.0125135f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.585
cc_12 VNB N_A_c_156_n 0.00557768f $X=-0.19 $Y=-0.245 $X2=3.85 $Y2=1.35
cc_13 VNB A 0.00199724f $X=-0.19 $Y=-0.245 $X2=5.435 $Y2=1.58
cc_14 VNB N_A_c_158_n 0.0195421f $X=-0.19 $Y=-0.245 $X2=5.225 $Y2=1.515
cc_15 VNB N_A_c_159_n 0.0420802f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=1.652
cc_16 VNB N_A_c_160_n 0.00798232f $X=-0.19 $Y=-0.245 $X2=4.39 $Y2=1.562
cc_17 VNB N_B_M1017_g 0.0256964f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.86
cc_18 VNB N_B_M1026_g 0.0260782f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.86
cc_19 VNB N_B_c_375_n 0.00564747f $X=-0.19 $Y=-0.245 $X2=4.725 $Y2=1.765
cc_20 VNB N_B_c_376_n 0.0179606f $X=-0.19 $Y=-0.245 $X2=4.725 $Y2=2.4
cc_21 VNB N_B_M1003_g 0.00619066f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=0.74
cc_22 VNB N_B_c_378_n 0.0283688f $X=-0.19 $Y=-0.245 $X2=5.315 $Y2=2.4
cc_23 VNB N_B_c_379_n 0.0115262f $X=-0.19 $Y=-0.245 $X2=5.335 $Y2=1.35
cc_24 VNB N_B_M1007_g 0.00656268f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=1.35
cc_25 VNB N_B_M1014_g 0.0230909f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=1.765
cc_26 VNB N_B_c_382_n 0.067871f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=2.4
cc_27 VNB N_B_M1019_g 0.0260971f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=0.74
cc_28 VNB N_B_c_384_n 0.00100736f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.42
cc_29 VNB N_B_c_385_n 0.0378918f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=0.665
cc_30 VNB N_B_c_386_n 4.22572e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_B_c_387_n 0.00498375f $X=-0.19 $Y=-0.245 $X2=5.45 $Y2=1.515
cc_32 VNB N_A_160_98#_c_578_n 0.020942f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=2.46
cc_33 VNB N_A_160_98#_c_579_n 0.020159f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=0.74
cc_34 VNB N_A_160_98#_c_580_n 0.0110058f $X=-0.19 $Y=-0.245 $X2=5.335 $Y2=1.35
cc_35 VNB N_A_160_98#_c_581_n 0.0692353f $X=-0.19 $Y=-0.245 $X2=5.335 $Y2=0.74
cc_36 VNB N_A_160_98#_c_582_n 0.009127f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=0.74
cc_37 VNB N_A_160_98#_c_583_n 0.00258679f $X=-0.19 $Y=-0.245 $X2=6.255 $Y2=1.485
cc_38 VNB N_A_160_98#_c_584_n 0.00234522f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=0.74
cc_39 VNB N_A_160_98#_c_585_n 0.00241736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_160_98#_c_586_n 0.00188856f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.585
cc_41 VNB N_VPWR_c_764_n 0.362705f $X=-0.19 $Y=-0.245 $X2=2.87 $Y2=0.685
cc_42 VNB N_X_c_998_n 0.00435724f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=1.35
cc_43 VNB N_X_c_999_n 0.00276895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_X_c_1000_n 0.0209692f $X=-0.19 $Y=-0.245 $X2=5.315 $Y2=2.4
cc_45 VNB N_X_c_1001_n 0.00207986f $X=-0.19 $Y=-0.245 $X2=5.335 $Y2=1.35
cc_46 VNB N_X_c_1002_n 0.0025951f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=2.4
cc_47 VNB N_X_c_1003_n 0.0112366f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=2.4
cc_48 VNB N_X_c_1004_n 0.0222851f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=0.74
cc_49 VNB N_X_c_1005_n 0.00345724f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.42
cc_50 VNB N_X_c_1006_n 0.00253527f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.585
cc_51 VNB N_X_c_1007_n 0.00124931f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.585
cc_52 VNB N_VGND_c_1170_n 0.01004f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=0.74
cc_53 VNB N_VGND_c_1171_n 0.0567336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1172_n 0.015878f $X=-0.19 $Y=-0.245 $X2=5.335 $Y2=1.35
cc_55 VNB N_VGND_c_1173_n 0.015091f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=1.35
cc_56 VNB N_VGND_c_1174_n 0.00790705f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=1.765
cc_57 VNB N_VGND_c_1175_n 0.0075298f $X=-0.19 $Y=-0.245 $X2=5.855 $Y2=1.485
cc_58 VNB N_VGND_c_1176_n 0.0218315f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=2.4
cc_59 VNB N_VGND_c_1177_n 0.0260634f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=2.4
cc_60 VNB N_VGND_c_1178_n 0.026797f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=1.485
cc_61 VNB N_VGND_c_1179_n 0.00795087f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=1.35
cc_62 VNB N_VGND_c_1180_n 0.0216203f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.585
cc_63 VNB N_VGND_c_1181_n 0.0202269f $X=-0.19 $Y=-0.245 $X2=3.04 $Y2=1.105
cc_64 VNB N_VGND_c_1182_n 0.0178371f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=0.675
cc_65 VNB N_VGND_c_1183_n 0.0576436f $X=-0.19 $Y=-0.245 $X2=5.11 $Y2=1.515
cc_66 VNB N_VGND_c_1184_n 0.471044f $X=-0.19 $Y=-0.245 $X2=5.11 $Y2=1.515
cc_67 VNB N_VGND_c_1185_n 0.00631222f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.42
cc_68 VNB N_VGND_c_1186_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=5.45 $Y2=1.557
cc_69 VNB N_VGND_c_1187_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=1.557
cc_70 VNB N_A_877_74#_c_1292_n 6.9777e-19 $X=-0.19 $Y=-0.245 $X2=5.315 $Y2=2.4
cc_71 VNB N_A_877_74#_c_1293_n 0.00163372f $X=-0.19 $Y=-0.245 $X2=5.335 $Y2=1.35
cc_72 VNB N_A_877_74#_c_1294_n 0.011697f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=0.74
cc_73 VNB N_A_877_74#_c_1295_n 0.0164799f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=2.4
cc_74 VNB N_A_877_74#_c_1296_n 0.00217595f $X=-0.19 $Y=-0.245 $X2=5.855
+ $Y2=1.485
cc_75 VNB N_A_877_74#_c_1297_n 0.00239138f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=1.35
cc_76 VNB N_A_877_74#_c_1298_n 0.00220733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VPB N_A_c_161_n 0.0205706f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=1.885
cc_78 VPB N_A_c_162_n 0.0153074f $X=-0.19 $Y=1.66 $X2=1.05 $Y2=1.885
cc_79 VPB N_A_c_163_n 0.0162726f $X=-0.19 $Y=1.66 $X2=4.725 $Y2=1.765
cc_80 VPB N_A_c_164_n 0.0164879f $X=-0.19 $Y=1.66 $X2=5.315 $Y2=1.765
cc_81 VPB N_A_c_165_n 0.0161133f $X=-0.19 $Y=1.66 $X2=5.765 $Y2=1.765
cc_82 VPB N_A_c_150_n 0.00606658f $X=-0.19 $Y=1.66 $X2=6.255 $Y2=1.485
cc_83 VPB N_A_c_151_n 0.0198301f $X=-0.19 $Y=1.66 $X2=5.855 $Y2=1.485
cc_84 VPB N_A_c_168_n 0.0167871f $X=-0.19 $Y=1.66 $X2=6.345 $Y2=1.765
cc_85 VPB N_A_c_153_n 0.00678804f $X=-0.19 $Y=1.66 $X2=4.605 $Y2=1.35
cc_86 VPB N_A_c_155_n 0.00422592f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=1.585
cc_87 VPB A 0.00936437f $X=-0.19 $Y=1.66 $X2=5.435 $Y2=1.58
cc_88 VPB N_A_c_158_n 0.0123696f $X=-0.19 $Y=1.66 $X2=5.225 $Y2=1.515
cc_89 VPB N_A_c_159_n 0.0409148f $X=-0.19 $Y=1.66 $X2=1.05 $Y2=1.652
cc_90 VPB N_A_c_160_n 0.0035835f $X=-0.19 $Y=1.66 $X2=4.39 $Y2=1.562
cc_91 VPB N_B_c_388_n 0.0145789f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=1.885
cc_92 VPB N_B_c_389_n 0.0169964f $X=-0.19 $Y=1.66 $X2=1.05 $Y2=1.885
cc_93 VPB N_B_c_376_n 6.28632e-19 $X=-0.19 $Y=1.66 $X2=4.725 $Y2=2.4
cc_94 VPB N_B_c_391_n 0.0202035f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_B_c_392_n 0.0155127f $X=-0.19 $Y=1.66 $X2=5.765 $Y2=0.74
cc_96 VPB N_B_c_393_n 0.0155109f $X=-0.19 $Y=1.66 $X2=5.765 $Y2=1.765
cc_97 VPB N_B_c_382_n 0.0332062f $X=-0.19 $Y=1.66 $X2=6.345 $Y2=2.4
cc_98 VPB N_B_c_395_n 0.0192217f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_B_c_385_n 0.0515999f $X=-0.19 $Y=1.66 $X2=1.275 $Y2=0.665
cc_100 VPB N_B_c_397_n 0.00968953f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=1.585
cc_101 VPB N_B_c_398_n 0.00163083f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.585
cc_102 VPB N_B_c_399_n 6.26324e-19 $X=-0.19 $Y=1.66 $X2=2.87 $Y2=0.685
cc_103 VPB N_B_c_387_n 0.0148779f $X=-0.19 $Y=1.66 $X2=5.45 $Y2=1.515
cc_104 VPB N_A_160_98#_c_587_n 0.0173997f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=0.86
cc_105 VPB N_A_160_98#_c_588_n 0.0147723f $X=-0.19 $Y=1.66 $X2=4.725 $Y2=2.4
cc_106 VPB N_A_160_98#_c_589_n 0.0147695f $X=-0.19 $Y=1.66 $X2=5.315 $Y2=1.765
cc_107 VPB N_A_160_98#_c_580_n 0.00800349f $X=-0.19 $Y=1.66 $X2=5.335 $Y2=1.35
cc_108 VPB N_A_160_98#_c_581_n 0.0395614f $X=-0.19 $Y=1.66 $X2=5.335 $Y2=0.74
cc_109 VPB N_A_160_98#_c_592_n 0.0147737f $X=-0.19 $Y=1.66 $X2=5.335 $Y2=0.74
cc_110 VPB N_A_160_98#_c_582_n 0.00528852f $X=-0.19 $Y=1.66 $X2=5.765 $Y2=0.74
cc_111 VPB N_A_160_98#_c_583_n 0.00107328f $X=-0.19 $Y=1.66 $X2=6.255 $Y2=1.485
cc_112 VPB N_A_160_98#_c_585_n 0.00170979f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_36_392#_c_718_n 0.0365351f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=0.86
cc_114 VPB N_A_36_392#_c_719_n 0.0090713f $X=-0.19 $Y=1.66 $X2=4.725 $Y2=2.4
cc_115 VPB N_A_36_392#_c_720_n 0.014517f $X=-0.19 $Y=1.66 $X2=4.725 $Y2=2.4
cc_116 VPB N_A_36_392#_c_721_n 0.00682979f $X=-0.19 $Y=1.66 $X2=5.315 $Y2=2.4
cc_117 VPB N_A_36_392#_c_722_n 0.00171072f $X=-0.19 $Y=1.66 $X2=5.335 $Y2=1.35
cc_118 VPB N_A_36_392#_c_723_n 0.00672394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_765_n 0.00847f $X=-0.19 $Y=1.66 $X2=4.745 $Y2=0.74
cc_120 VPB N_VPWR_c_766_n 0.00512608f $X=-0.19 $Y=1.66 $X2=5.315 $Y2=2.4
cc_121 VPB N_VPWR_c_767_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_768_n 0.0908858f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_769_n 0.018101f $X=-0.19 $Y=1.66 $X2=6.345 $Y2=2.4
cc_124 VPB N_VPWR_c_770_n 0.0175244f $X=-0.19 $Y=1.66 $X2=4.82 $Y2=1.515
cc_125 VPB N_VPWR_c_771_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.42
cc_126 VPB N_VPWR_c_772_n 0.0197879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_764_n 0.102501f $X=-0.19 $Y=1.66 $X2=2.87 $Y2=0.685
cc_128 VPB N_VPWR_c_774_n 0.0263173f $X=-0.19 $Y=1.66 $X2=2.955 $Y2=1.02
cc_129 VPB N_VPWR_c_775_n 0.0141241f $X=-0.19 $Y=1.66 $X2=3.85 $Y2=1.19
cc_130 VPB N_VPWR_c_776_n 0.0138912f $X=-0.19 $Y=1.66 $X2=5.435 $Y2=1.58
cc_131 VPB N_VPWR_c_777_n 0.00460249f $X=-0.19 $Y=1.66 $X2=5.11 $Y2=1.515
cc_132 VPB N_VPWR_c_778_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.652
cc_133 VPB N_A_514_368#_c_881_n 0.00662236f $X=-0.19 $Y=1.66 $X2=5.315 $Y2=2.4
cc_134 VPB N_A_514_368#_c_882_n 0.0030474f $X=-0.19 $Y=1.66 $X2=5.335 $Y2=0.74
cc_135 VPB N_A_514_368#_c_883_n 0.00377007f $X=-0.19 $Y=1.66 $X2=5.335 $Y2=0.74
cc_136 VPB N_A_514_368#_c_884_n 0.00328226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_514_368#_c_885_n 0.00179305f $X=-0.19 $Y=1.66 $X2=6.345 $Y2=2.4
cc_138 VPB N_A_514_368#_c_886_n 0.00121438f $X=-0.19 $Y=1.66 $X2=6.345 $Y2=1.35
cc_139 VPB N_A_514_368#_c_887_n 0.00190506f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.75
cc_140 VPB N_A_514_368#_c_888_n 0.002547f $X=-0.19 $Y=1.66 $X2=2.87 $Y2=0.685
cc_141 VPB N_A_514_368#_c_889_n 0.00257417f $X=-0.19 $Y=1.66 $X2=3.85 $Y2=1.19
cc_142 VPB N_A_514_368#_c_890_n 0.0309665f $X=-0.19 $Y=1.66 $X2=1.275 $Y2=0.675
cc_143 VPB N_X_c_1008_n 0.00692367f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_X_c_1004_n 0.00836399f $X=-0.19 $Y=1.66 $X2=6.355 $Y2=0.74
cc_145 N_A_c_162_n N_B_c_388_n 0.00830807f $X=1.05 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_146 N_A_M1016_g N_B_M1017_g 0.0289814f $X=1.155 $Y=0.86 $X2=0 $Y2=0
cc_147 N_A_c_177_p N_B_M1017_g 0.0124999f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_148 N_A_c_178_p N_B_M1017_g 5.1812e-19 $X=1.445 $Y=0.675 $X2=0 $Y2=0
cc_149 N_A_c_177_p N_B_M1026_g 0.0125312f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_150 N_A_c_180_p N_B_M1026_g 9.06409e-19 $X=2.955 $Y=1.02 $X2=0 $Y2=0
cc_151 N_A_M1024_g N_B_c_375_n 0.00858677f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_c_150_n N_B_c_376_n 0.0196758f $X=6.255 $Y=1.485 $X2=0 $Y2=0
cc_153 N_A_c_168_n N_B_c_391_n 0.026502f $X=6.345 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A_M1024_g N_B_c_379_n 0.024894f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_c_185_p N_B_c_385_n 0.00117645f $X=0.945 $Y=1.585 $X2=0 $Y2=0
cc_156 N_A_c_159_n N_B_c_385_n 0.02171f $X=1.05 $Y=1.652 $X2=0 $Y2=0
cc_157 N_A_c_163_n N_B_c_413_n 0.0113493f $X=4.725 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A_c_164_n N_B_c_413_n 0.011363f $X=5.315 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A_c_165_n N_B_c_413_n 0.0133065f $X=5.765 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A_c_151_n N_B_c_413_n 0.0011792f $X=5.855 $Y=1.485 $X2=0 $Y2=0
cc_161 N_A_c_168_n N_B_c_413_n 6.68492e-19 $X=6.345 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A_c_153_n N_B_c_413_n 0.0020905f $X=4.605 $Y=1.35 $X2=0 $Y2=0
cc_163 A N_B_c_413_n 0.0880524f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A_c_160_n N_B_c_413_n 0.0363523f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_165 N_A_c_165_n N_B_c_386_n 4.43582e-19 $X=5.765 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A_c_150_n N_B_c_386_n 0.00998843f $X=6.255 $Y=1.485 $X2=0 $Y2=0
cc_167 N_A_c_151_n N_B_c_386_n 0.00732481f $X=5.855 $Y=1.485 $X2=0 $Y2=0
cc_168 A N_B_c_386_n 0.031682f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_169 N_A_c_164_n N_B_c_399_n 8.14491e-19 $X=5.315 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A_c_165_n N_B_c_399_n 0.00460047f $X=5.765 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A_c_168_n N_B_c_399_n 0.00310756f $X=6.345 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A_c_202_p N_B_c_428_n 0.00146532f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_173 N_A_c_150_n N_B_c_387_n 0.0308523f $X=6.255 $Y=1.485 $X2=0 $Y2=0
cc_174 N_A_c_168_n N_B_c_387_n 0.00269426f $X=6.345 $Y=1.765 $X2=0 $Y2=0
cc_175 N_A_c_205_p N_A_160_98#_M1000_d 0.00439657f $X=1.275 $Y=0.675 $X2=-0.19
+ $Y2=-0.245
cc_176 N_A_c_177_p N_A_160_98#_M1017_d 0.00782857f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_177 N_A_c_177_p N_A_160_98#_c_578_n 0.0115801f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_178 N_A_c_180_p N_A_160_98#_c_578_n 0.00775701f $X=2.955 $Y=1.02 $X2=0 $Y2=0
cc_179 N_A_c_209_p N_A_160_98#_c_578_n 0.00681965f $X=3.04 $Y=1.105 $X2=0 $Y2=0
cc_180 N_A_c_180_p N_A_160_98#_c_579_n 0.00271318f $X=2.955 $Y=1.02 $X2=0 $Y2=0
cc_181 N_A_c_202_p N_A_160_98#_c_579_n 0.0140111f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_182 N_A_c_156_n N_A_160_98#_c_579_n 0.00585519f $X=3.85 $Y=1.35 $X2=0 $Y2=0
cc_183 N_A_c_160_n N_A_160_98#_c_589_n 3.10764e-19 $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_184 N_A_c_160_n N_A_160_98#_c_580_n 0.0138757f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_185 N_A_c_177_p N_A_160_98#_c_581_n 0.00181746f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_186 N_A_c_202_p N_A_160_98#_c_581_n 0.0113772f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_187 N_A_c_160_n N_A_160_98#_c_581_n 0.0151457f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_188 N_A_c_163_n N_A_160_98#_c_592_n 0.0424336f $X=4.725 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A_c_160_n N_A_160_98#_c_592_n 0.0024566f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_190 N_A_c_153_n N_A_160_98#_c_582_n 0.0123305f $X=4.605 $Y=1.35 $X2=0 $Y2=0
cc_191 N_A_c_160_n N_A_160_98#_c_582_n 0.010912f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_192 N_A_M1016_g N_A_160_98#_c_613_n 0.0139847f $X=1.155 $Y=0.86 $X2=0 $Y2=0
cc_193 N_A_c_185_p N_A_160_98#_c_613_n 2.60315e-19 $X=0.945 $Y=1.585 $X2=0 $Y2=0
cc_194 N_A_c_205_p N_A_160_98#_c_613_n 0.00795398f $X=1.275 $Y=0.675 $X2=0 $Y2=0
cc_195 N_A_c_178_p N_A_160_98#_c_613_n 0.0204402f $X=1.445 $Y=0.675 $X2=0 $Y2=0
cc_196 N_A_c_162_n N_A_160_98#_c_583_n 4.29131e-19 $X=1.05 $Y=1.885 $X2=0 $Y2=0
cc_197 N_A_M1016_g N_A_160_98#_c_583_n 0.00431001f $X=1.155 $Y=0.86 $X2=0 $Y2=0
cc_198 N_A_c_185_p N_A_160_98#_c_583_n 0.0118099f $X=0.945 $Y=1.585 $X2=0 $Y2=0
cc_199 N_A_c_159_n N_A_160_98#_c_583_n 0.00171544f $X=1.05 $Y=1.652 $X2=0 $Y2=0
cc_200 N_A_c_177_p N_A_160_98#_c_621_n 0.053955f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_201 N_A_c_180_p N_A_160_98#_c_621_n 0.00628036f $X=2.955 $Y=1.02 $X2=0 $Y2=0
cc_202 N_A_c_209_p N_A_160_98#_c_621_n 0.0148586f $X=3.04 $Y=1.105 $X2=0 $Y2=0
cc_203 N_A_c_177_p N_A_160_98#_c_624_n 0.00371196f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_204 N_A_c_202_p N_A_160_98#_c_624_n 0.0385816f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_205 N_A_c_209_p N_A_160_98#_c_624_n 0.0111271f $X=3.04 $Y=1.105 $X2=0 $Y2=0
cc_206 N_A_c_160_n N_A_160_98#_c_624_n 0.0213902f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_207 N_A_M1016_g N_A_160_98#_c_586_n 0.00279462f $X=1.155 $Y=0.86 $X2=0 $Y2=0
cc_208 N_A_c_154_n N_A_160_98#_c_586_n 0.0118907f $X=0.6 $Y=1.42 $X2=0 $Y2=0
cc_209 N_A_c_185_p N_A_160_98#_c_586_n 0.0196847f $X=0.945 $Y=1.585 $X2=0 $Y2=0
cc_210 N_A_c_205_p N_A_160_98#_c_586_n 0.0144338f $X=1.275 $Y=0.675 $X2=0 $Y2=0
cc_211 N_A_c_159_n N_A_160_98#_c_586_n 0.00236202f $X=1.05 $Y=1.652 $X2=0 $Y2=0
cc_212 N_A_c_177_p N_A_160_98#_c_633_n 0.0149765f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_213 N_A_c_161_n N_A_36_392#_c_718_n 0.0110352f $X=0.55 $Y=1.885 $X2=0 $Y2=0
cc_214 N_A_c_162_n N_A_36_392#_c_718_n 7.07825e-19 $X=1.05 $Y=1.885 $X2=0 $Y2=0
cc_215 N_A_c_161_n N_A_36_392#_c_719_n 0.0122751f $X=0.55 $Y=1.885 $X2=0 $Y2=0
cc_216 N_A_c_162_n N_A_36_392#_c_719_n 0.0136119f $X=1.05 $Y=1.885 $X2=0 $Y2=0
cc_217 N_A_c_155_n N_A_36_392#_c_719_n 0.0149347f $X=0.685 $Y=1.585 $X2=0 $Y2=0
cc_218 N_A_c_185_p N_A_36_392#_c_719_n 0.0313645f $X=0.945 $Y=1.585 $X2=0 $Y2=0
cc_219 N_A_c_159_n N_A_36_392#_c_719_n 0.0125714f $X=1.05 $Y=1.652 $X2=0 $Y2=0
cc_220 N_A_c_161_n N_A_36_392#_c_720_n 0.00123848f $X=0.55 $Y=1.885 $X2=0 $Y2=0
cc_221 N_A_c_155_n N_A_36_392#_c_720_n 0.00416948f $X=0.685 $Y=1.585 $X2=0 $Y2=0
cc_222 N_A_c_159_n N_A_36_392#_c_720_n 5.99033e-19 $X=1.05 $Y=1.652 $X2=0 $Y2=0
cc_223 N_A_c_161_n N_A_36_392#_c_734_n 5.95972e-19 $X=0.55 $Y=1.885 $X2=0 $Y2=0
cc_224 N_A_c_162_n N_A_36_392#_c_734_n 0.00927516f $X=1.05 $Y=1.885 $X2=0 $Y2=0
cc_225 N_A_c_162_n N_A_36_392#_c_722_n 0.00312124f $X=1.05 $Y=1.885 $X2=0 $Y2=0
cc_226 N_A_c_161_n N_VPWR_c_765_n 0.0054463f $X=0.55 $Y=1.885 $X2=0 $Y2=0
cc_227 N_A_c_162_n N_VPWR_c_765_n 0.00508297f $X=1.05 $Y=1.885 $X2=0 $Y2=0
cc_228 N_A_c_168_n N_VPWR_c_766_n 3.91613e-19 $X=6.345 $Y=1.765 $X2=0 $Y2=0
cc_229 N_A_c_162_n N_VPWR_c_768_n 0.0044313f $X=1.05 $Y=1.885 $X2=0 $Y2=0
cc_230 N_A_c_163_n N_VPWR_c_768_n 0.00312499f $X=4.725 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A_c_164_n N_VPWR_c_769_n 0.00312629f $X=5.315 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A_c_165_n N_VPWR_c_769_n 0.00361464f $X=5.765 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A_c_168_n N_VPWR_c_770_n 0.00314961f $X=6.345 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A_c_161_n N_VPWR_c_764_n 0.00861685f $X=0.55 $Y=1.885 $X2=0 $Y2=0
cc_235 N_A_c_162_n N_VPWR_c_764_n 0.00853234f $X=1.05 $Y=1.885 $X2=0 $Y2=0
cc_236 N_A_c_163_n N_VPWR_c_764_n 0.00386659f $X=4.725 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A_c_164_n N_VPWR_c_764_n 0.00388054f $X=5.315 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A_c_165_n N_VPWR_c_764_n 0.00560771f $X=5.765 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A_c_168_n N_VPWR_c_764_n 0.003911f $X=6.345 $Y=1.765 $X2=0 $Y2=0
cc_240 N_A_c_161_n N_VPWR_c_774_n 0.00445602f $X=0.55 $Y=1.885 $X2=0 $Y2=0
cc_241 N_A_c_163_n N_VPWR_c_775_n 0.00148242f $X=4.725 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A_c_164_n N_VPWR_c_775_n 0.00333649f $X=5.315 $Y=1.765 $X2=0 $Y2=0
cc_243 N_A_c_165_n N_VPWR_c_776_n 0.00334336f $X=5.765 $Y=1.765 $X2=0 $Y2=0
cc_244 N_A_c_168_n N_VPWR_c_776_n 0.00192155f $X=6.345 $Y=1.765 $X2=0 $Y2=0
cc_245 N_A_c_165_n N_A_514_368#_c_891_n 0.00828871f $X=5.765 $Y=1.765 $X2=0
+ $Y2=0
cc_246 N_A_c_168_n N_A_514_368#_c_891_n 0.0110022f $X=6.345 $Y=1.765 $X2=0 $Y2=0
cc_247 N_A_c_168_n N_A_514_368#_c_885_n 0.00346639f $X=6.345 $Y=1.765 $X2=0
+ $Y2=0
cc_248 N_A_c_163_n N_A_514_368#_c_887_n 0.00650778f $X=4.725 $Y=1.765 $X2=0
+ $Y2=0
cc_249 N_A_c_164_n N_A_514_368#_c_887_n 8.60548e-19 $X=5.315 $Y=1.765 $X2=0
+ $Y2=0
cc_250 N_A_c_163_n N_A_514_368#_c_896_n 0.00971339f $X=4.725 $Y=1.765 $X2=0
+ $Y2=0
cc_251 N_A_c_164_n N_A_514_368#_c_896_n 0.00916701f $X=5.315 $Y=1.765 $X2=0
+ $Y2=0
cc_252 N_A_c_163_n N_A_514_368#_c_888_n 7.59211e-19 $X=4.725 $Y=1.765 $X2=0
+ $Y2=0
cc_253 N_A_c_164_n N_A_514_368#_c_888_n 0.00429318f $X=5.315 $Y=1.765 $X2=0
+ $Y2=0
cc_254 N_A_c_165_n N_A_514_368#_c_888_n 0.00426546f $X=5.765 $Y=1.765 $X2=0
+ $Y2=0
cc_255 N_A_c_168_n N_A_514_368#_c_888_n 7.63182e-19 $X=6.345 $Y=1.765 $X2=0
+ $Y2=0
cc_256 N_A_c_177_p N_X_M1008_s 0.00223669f $X=2.87 $Y=0.685 $X2=-0.19 $Y2=-0.245
cc_257 N_A_c_180_p N_X_M1008_s 0.00327917f $X=2.955 $Y=1.02 $X2=-0.19 $Y2=-0.245
cc_258 N_A_c_202_p N_X_M1008_s 0.0144824f $X=3.765 $Y=1.105 $X2=-0.19 $Y2=-0.245
cc_259 N_A_c_209_p N_X_M1008_s 3.64502e-19 $X=3.04 $Y=1.105 $X2=-0.19 $Y2=-0.245
cc_260 N_A_c_202_p N_X_c_998_n 0.0250503f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_261 N_A_c_160_n N_X_c_998_n 0.00617915f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_262 N_A_M1009_g N_X_c_999_n 0.00402271f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_c_163_n N_X_c_1017_n 0.0113487f $X=4.725 $Y=1.765 $X2=0 $Y2=0
cc_264 N_A_c_164_n N_X_c_1017_n 0.0114141f $X=5.315 $Y=1.765 $X2=0 $Y2=0
cc_265 N_A_c_165_n N_X_c_1017_n 0.0113061f $X=5.765 $Y=1.765 $X2=0 $Y2=0
cc_266 N_A_c_150_n N_X_c_1017_n 9.97318e-19 $X=6.255 $Y=1.485 $X2=0 $Y2=0
cc_267 N_A_c_168_n N_X_c_1017_n 0.00546153f $X=6.345 $Y=1.765 $X2=0 $Y2=0
cc_268 N_A_M1009_g N_X_c_1000_n 0.0131565f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_M1010_g N_X_c_1000_n 0.0112941f $X=5.335 $Y=0.74 $X2=0 $Y2=0
cc_270 N_A_M1020_g N_X_c_1000_n 0.0150594f $X=5.765 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A_c_150_n N_X_c_1000_n 0.00494416f $X=6.255 $Y=1.485 $X2=0 $Y2=0
cc_272 N_A_c_151_n N_X_c_1000_n 0.00224206f $X=5.855 $Y=1.485 $X2=0 $Y2=0
cc_273 N_A_M1024_g N_X_c_1000_n 0.0112465f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A_c_153_n N_X_c_1000_n 0.00155242f $X=4.605 $Y=1.35 $X2=0 $Y2=0
cc_275 A N_X_c_1000_n 0.0950924f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_276 N_A_c_158_n N_X_c_1000_n 0.00582934f $X=5.225 $Y=1.515 $X2=0 $Y2=0
cc_277 N_A_c_160_n N_X_c_1000_n 0.00930879f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_278 N_A_c_202_p N_X_c_1001_n 0.0144259f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_279 N_A_c_160_n N_X_c_1001_n 0.0150081f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_280 N_A_c_165_n N_X_c_1034_n 0.00307027f $X=5.765 $Y=1.765 $X2=0 $Y2=0
cc_281 N_A_c_168_n N_X_c_1034_n 0.00468176f $X=6.345 $Y=1.765 $X2=0 $Y2=0
cc_282 N_A_c_168_n N_X_c_1008_n 0.00773372f $X=6.345 $Y=1.765 $X2=0 $Y2=0
cc_283 N_A_c_165_n N_X_c_1037_n 6.5518e-19 $X=5.765 $Y=1.765 $X2=0 $Y2=0
cc_284 N_A_c_150_n N_X_c_1037_n 4.83713e-19 $X=6.255 $Y=1.485 $X2=0 $Y2=0
cc_285 N_A_c_168_n N_X_c_1037_n 0.0030306f $X=6.345 $Y=1.765 $X2=0 $Y2=0
cc_286 N_A_M1024_g N_X_c_1040_n 7.61432e-19 $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A_c_177_p N_X_c_1005_n 0.0144777f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_288 N_A_c_180_p N_X_c_1005_n 0.00607737f $X=2.955 $Y=1.02 $X2=0 $Y2=0
cc_289 N_A_c_202_p N_X_c_1005_n 0.0208829f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_290 N_A_c_163_n N_X_c_1044_n 7.64699e-19 $X=4.725 $Y=1.765 $X2=0 $Y2=0
cc_291 N_A_c_154_n N_VGND_M1000_s 0.00510428f $X=0.6 $Y=1.42 $X2=-0.19
+ $Y2=-0.245
cc_292 N_A_c_322_p N_VGND_M1000_s 0.00321586f $X=0.685 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_293 N_A_c_177_p N_VGND_M1016_s 0.00394843f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_294 N_A_c_178_p N_VGND_M1016_s 0.00392577f $X=1.445 $Y=0.675 $X2=0 $Y2=0
cc_295 N_A_c_177_p N_VGND_M1026_s 0.00765915f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_296 N_A_c_202_p N_VGND_M1027_d 0.00594424f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_297 N_A_c_156_n N_VGND_M1027_d 0.0021153f $X=3.85 $Y=1.35 $X2=0 $Y2=0
cc_298 N_A_M1000_g N_VGND_c_1171_n 0.0103672f $X=0.725 $Y=0.86 $X2=0 $Y2=0
cc_299 N_A_c_154_n N_VGND_c_1171_n 0.0374154f $X=0.6 $Y=1.42 $X2=0 $Y2=0
cc_300 N_A_c_322_p N_VGND_c_1171_n 0.0141996f $X=0.685 $Y=0.665 $X2=0 $Y2=0
cc_301 N_A_c_177_p N_VGND_c_1172_n 0.0247182f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_302 N_A_M1009_g N_VGND_c_1173_n 0.00348294f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_303 N_A_M1009_g N_VGND_c_1174_n 0.00416335f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_304 N_A_M1010_g N_VGND_c_1174_n 0.00418252f $X=5.335 $Y=0.74 $X2=0 $Y2=0
cc_305 N_A_M1020_g N_VGND_c_1175_n 0.00418252f $X=5.765 $Y=0.74 $X2=0 $Y2=0
cc_306 N_A_M1024_g N_VGND_c_1175_n 0.00231005f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A_M1016_g N_VGND_c_1176_n 0.0014541f $X=1.155 $Y=0.86 $X2=0 $Y2=0
cc_308 N_A_c_177_p N_VGND_c_1176_n 0.0114916f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_309 N_A_c_178_p N_VGND_c_1176_n 0.0119842f $X=1.445 $Y=0.675 $X2=0 $Y2=0
cc_310 N_A_M1000_g N_VGND_c_1177_n 0.00374701f $X=0.725 $Y=0.86 $X2=0 $Y2=0
cc_311 N_A_M1016_g N_VGND_c_1177_n 0.00374721f $X=1.155 $Y=0.86 $X2=0 $Y2=0
cc_312 N_A_c_322_p N_VGND_c_1177_n 0.00306302f $X=0.685 $Y=0.665 $X2=0 $Y2=0
cc_313 N_A_c_205_p N_VGND_c_1177_n 0.0101323f $X=1.275 $Y=0.675 $X2=0 $Y2=0
cc_314 N_A_c_177_p N_VGND_c_1178_n 0.00464991f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_315 N_A_c_177_p N_VGND_c_1180_n 0.0129334f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_316 N_A_M1009_g N_VGND_c_1181_n 0.00324657f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A_M1010_g N_VGND_c_1182_n 0.00323547f $X=5.335 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A_M1020_g N_VGND_c_1182_n 0.00323547f $X=5.765 $Y=0.74 $X2=0 $Y2=0
cc_319 N_A_M1024_g N_VGND_c_1183_n 0.00321293f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A_M1000_g N_VGND_c_1184_n 0.00508379f $X=0.725 $Y=0.86 $X2=0 $Y2=0
cc_321 N_A_M1016_g N_VGND_c_1184_n 0.00508379f $X=1.155 $Y=0.86 $X2=0 $Y2=0
cc_322 N_A_M1009_g N_VGND_c_1184_n 0.00416139f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_323 N_A_M1010_g N_VGND_c_1184_n 0.00412104f $X=5.335 $Y=0.74 $X2=0 $Y2=0
cc_324 N_A_M1020_g N_VGND_c_1184_n 0.00412104f $X=5.765 $Y=0.74 $X2=0 $Y2=0
cc_325 N_A_M1024_g N_VGND_c_1184_n 0.0041125f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_326 N_A_c_322_p N_VGND_c_1184_n 0.00533032f $X=0.685 $Y=0.665 $X2=0 $Y2=0
cc_327 N_A_c_177_p N_VGND_c_1184_n 0.0344715f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_328 N_A_c_205_p N_VGND_c_1184_n 0.0176507f $X=1.275 $Y=0.675 $X2=0 $Y2=0
cc_329 N_A_c_178_p N_VGND_c_1184_n 7.98341e-19 $X=1.445 $Y=0.675 $X2=0 $Y2=0
cc_330 N_A_M1020_g N_A_877_74#_c_1299_n 0.00927675f $X=5.765 $Y=0.74 $X2=0 $Y2=0
cc_331 N_A_M1024_g N_A_877_74#_c_1299_n 0.00927675f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_332 N_A_M1020_g N_A_877_74#_c_1301_n 7.8287e-19 $X=5.765 $Y=0.74 $X2=0 $Y2=0
cc_333 N_A_M1024_g N_A_877_74#_c_1301_n 0.00539834f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_334 N_A_M1024_g N_A_877_74#_c_1293_n 0.0039285f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_335 N_A_M1009_g N_A_877_74#_c_1296_n 0.00838898f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_336 N_A_M1010_g N_A_877_74#_c_1296_n 7.98198e-19 $X=5.335 $Y=0.74 $X2=0 $Y2=0
cc_337 N_A_M1009_g N_A_877_74#_c_1306_n 0.00927675f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_338 N_A_M1010_g N_A_877_74#_c_1306_n 0.00927675f $X=5.335 $Y=0.74 $X2=0 $Y2=0
cc_339 N_A_M1009_g N_A_877_74#_c_1297_n 7.98516e-19 $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_340 N_A_M1010_g N_A_877_74#_c_1297_n 0.00763599f $X=5.335 $Y=0.74 $X2=0 $Y2=0
cc_341 N_A_M1020_g N_A_877_74#_c_1297_n 0.00763599f $X=5.765 $Y=0.74 $X2=0 $Y2=0
cc_342 N_A_M1024_g N_A_877_74#_c_1297_n 7.98516e-19 $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_343 N_B_M1026_g N_A_160_98#_c_578_n 0.0239678f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_344 N_B_c_384_n N_A_160_98#_c_587_n 5.46419e-19 $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_345 N_B_c_385_n N_A_160_98#_c_587_n 0.00225337f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_346 N_B_c_397_n N_A_160_98#_c_587_n 0.0167551f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_347 N_B_c_397_n N_A_160_98#_c_588_n 0.00984894f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_348 N_B_c_413_n N_A_160_98#_c_589_n 0.0109565f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_349 N_B_c_428_n N_A_160_98#_c_589_n 0.00246188f $X=3.57 $Y=1.935 $X2=0 $Y2=0
cc_350 N_B_c_413_n N_A_160_98#_c_580_n 0.00192852f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_351 N_B_M1026_g N_A_160_98#_c_581_n 0.0193036f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_352 N_B_c_384_n N_A_160_98#_c_581_n 7.08336e-19 $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_353 N_B_c_385_n N_A_160_98#_c_581_n 0.0025678f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_354 N_B_c_397_n N_A_160_98#_c_581_n 0.00985098f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_355 N_B_c_413_n N_A_160_98#_c_581_n 0.00188169f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_356 N_B_c_428_n N_A_160_98#_c_581_n 0.00473887f $X=3.57 $Y=1.935 $X2=0 $Y2=0
cc_357 N_B_c_413_n N_A_160_98#_c_592_n 0.0106242f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_358 N_B_c_385_n N_A_160_98#_c_613_n 0.00498833f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_359 N_B_c_388_n N_A_160_98#_c_583_n 0.0104911f $X=1.5 $Y=1.885 $X2=0 $Y2=0
cc_360 N_B_M1017_g N_A_160_98#_c_583_n 0.0104353f $X=1.745 $Y=0.86 $X2=0 $Y2=0
cc_361 N_B_c_389_n N_A_160_98#_c_583_n 0.00664878f $X=1.95 $Y=1.885 $X2=0 $Y2=0
cc_362 N_B_M1026_g N_A_160_98#_c_583_n 0.00149841f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_363 N_B_c_384_n N_A_160_98#_c_583_n 0.0229329f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_364 N_B_c_385_n N_A_160_98#_c_583_n 0.0287848f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_365 N_B_c_398_n N_A_160_98#_c_583_n 0.00966187f $X=2.36 $Y=1.935 $X2=0 $Y2=0
cc_366 N_B_M1017_g N_A_160_98#_c_621_n 6.52662e-19 $X=1.745 $Y=0.86 $X2=0 $Y2=0
cc_367 N_B_M1026_g N_A_160_98#_c_621_n 0.0117669f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_368 N_B_c_384_n N_A_160_98#_c_621_n 0.0158037f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_369 N_B_c_385_n N_A_160_98#_c_621_n 0.0052093f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_370 N_B_c_397_n N_A_160_98#_c_621_n 0.00402169f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_371 N_B_M1026_g N_A_160_98#_c_584_n 0.0037313f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_372 N_B_M1026_g N_A_160_98#_c_585_n 0.0044251f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_373 N_B_c_384_n N_A_160_98#_c_585_n 0.01771f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_374 N_B_c_397_n N_A_160_98#_c_585_n 0.0136221f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_375 N_B_c_397_n N_A_160_98#_c_624_n 0.0495782f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_376 N_B_c_428_n N_A_160_98#_c_624_n 0.00752433f $X=3.57 $Y=1.935 $X2=0 $Y2=0
cc_377 N_B_M1017_g N_A_160_98#_c_633_n 0.0093952f $X=1.745 $Y=0.86 $X2=0 $Y2=0
cc_378 N_B_c_398_n N_A_36_392#_M1006_s 0.00239688f $X=2.36 $Y=1.935 $X2=0 $Y2=0
cc_379 N_B_c_388_n N_A_36_392#_c_719_n 9.21122e-19 $X=1.5 $Y=1.885 $X2=0 $Y2=0
cc_380 N_B_c_388_n N_A_36_392#_c_721_n 0.0128006f $X=1.5 $Y=1.885 $X2=0 $Y2=0
cc_381 N_B_c_389_n N_A_36_392#_c_721_n 0.0134708f $X=1.95 $Y=1.885 $X2=0 $Y2=0
cc_382 N_B_c_388_n N_A_36_392#_c_723_n 6.49809e-19 $X=1.5 $Y=1.885 $X2=0 $Y2=0
cc_383 N_B_c_389_n N_A_36_392#_c_723_n 0.0107987f $X=1.95 $Y=1.885 $X2=0 $Y2=0
cc_384 N_B_c_385_n N_A_36_392#_c_723_n 0.00146311f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_385 N_B_c_398_n N_A_36_392#_c_723_n 0.0229474f $X=2.36 $Y=1.935 $X2=0 $Y2=0
cc_386 N_B_c_413_n N_VPWR_M1005_s 0.00704523f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_387 N_B_c_413_n N_VPWR_M1025_s 0.00243402f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_388 N_B_c_399_n N_VPWR_M1025_s 0.00133155f $X=5.89 $Y=1.945 $X2=0 $Y2=0
cc_389 N_B_c_391_n N_VPWR_c_766_n 0.00729564f $X=6.795 $Y=1.765 $X2=0 $Y2=0
cc_390 N_B_c_392_n N_VPWR_c_766_n 0.00409001f $X=7.245 $Y=1.765 $X2=0 $Y2=0
cc_391 N_B_c_393_n N_VPWR_c_767_n 0.00379374f $X=7.695 $Y=1.765 $X2=0 $Y2=0
cc_392 N_B_c_395_n N_VPWR_c_767_n 0.00379374f $X=8.145 $Y=1.765 $X2=0 $Y2=0
cc_393 N_B_c_388_n N_VPWR_c_768_n 0.00278271f $X=1.5 $Y=1.885 $X2=0 $Y2=0
cc_394 N_B_c_389_n N_VPWR_c_768_n 0.00278257f $X=1.95 $Y=1.885 $X2=0 $Y2=0
cc_395 N_B_c_391_n N_VPWR_c_770_n 0.00413917f $X=6.795 $Y=1.765 $X2=0 $Y2=0
cc_396 N_B_c_392_n N_VPWR_c_771_n 0.00445602f $X=7.245 $Y=1.765 $X2=0 $Y2=0
cc_397 N_B_c_393_n N_VPWR_c_771_n 0.00445602f $X=7.695 $Y=1.765 $X2=0 $Y2=0
cc_398 N_B_c_395_n N_VPWR_c_772_n 0.00445602f $X=8.145 $Y=1.765 $X2=0 $Y2=0
cc_399 N_B_c_388_n N_VPWR_c_764_n 0.00353907f $X=1.5 $Y=1.885 $X2=0 $Y2=0
cc_400 N_B_c_389_n N_VPWR_c_764_n 0.00358623f $X=1.95 $Y=1.885 $X2=0 $Y2=0
cc_401 N_B_c_391_n N_VPWR_c_764_n 0.0081781f $X=6.795 $Y=1.765 $X2=0 $Y2=0
cc_402 N_B_c_392_n N_VPWR_c_764_n 0.00857589f $X=7.245 $Y=1.765 $X2=0 $Y2=0
cc_403 N_B_c_393_n N_VPWR_c_764_n 0.00857589f $X=7.695 $Y=1.765 $X2=0 $Y2=0
cc_404 N_B_c_395_n N_VPWR_c_764_n 0.0086105f $X=8.145 $Y=1.765 $X2=0 $Y2=0
cc_405 N_B_c_397_n N_A_514_368#_M1004_d 0.00539645f $X=3.485 $Y=1.935 $X2=-0.19
+ $Y2=-0.245
cc_406 N_B_c_413_n N_A_514_368#_M1012_d 0.00128952f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_407 N_B_c_428_n N_A_514_368#_M1012_d 0.00467648f $X=3.57 $Y=1.935 $X2=0 $Y2=0
cc_408 N_B_c_413_n N_A_514_368#_M1029_d 0.00396407f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_409 N_B_c_413_n N_A_514_368#_M1013_d 0.00359524f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_410 N_B_c_389_n N_A_514_368#_c_881_n 0.0012003f $X=1.95 $Y=1.885 $X2=0 $Y2=0
cc_411 N_B_c_397_n N_A_514_368#_c_881_n 0.0202824f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_412 N_B_c_389_n N_A_514_368#_c_883_n 5.76545e-19 $X=1.95 $Y=1.885 $X2=0 $Y2=0
cc_413 N_B_c_391_n N_A_514_368#_c_885_n 0.00145414f $X=6.795 $Y=1.765 $X2=0
+ $Y2=0
cc_414 N_B_c_391_n N_A_514_368#_c_911_n 0.0124723f $X=6.795 $Y=1.765 $X2=0 $Y2=0
cc_415 N_B_c_392_n N_A_514_368#_c_911_n 0.0117449f $X=7.245 $Y=1.765 $X2=0 $Y2=0
cc_416 N_B_c_393_n N_A_514_368#_c_913_n 0.011796f $X=7.695 $Y=1.765 $X2=0 $Y2=0
cc_417 N_B_c_395_n N_A_514_368#_c_913_n 0.011796f $X=8.145 $Y=1.765 $X2=0 $Y2=0
cc_418 N_B_c_391_n N_A_514_368#_c_889_n 5.87784e-19 $X=6.795 $Y=1.765 $X2=0
+ $Y2=0
cc_419 N_B_c_392_n N_A_514_368#_c_889_n 0.00750751f $X=7.245 $Y=1.765 $X2=0
+ $Y2=0
cc_420 N_B_c_393_n N_A_514_368#_c_889_n 0.00730551f $X=7.695 $Y=1.765 $X2=0
+ $Y2=0
cc_421 N_B_c_395_n N_A_514_368#_c_889_n 5.64076e-19 $X=8.145 $Y=1.765 $X2=0
+ $Y2=0
cc_422 N_B_c_393_n N_A_514_368#_c_890_n 5.64076e-19 $X=7.695 $Y=1.765 $X2=0
+ $Y2=0
cc_423 N_B_c_395_n N_A_514_368#_c_890_n 0.00745145f $X=8.145 $Y=1.765 $X2=0
+ $Y2=0
cc_424 N_B_c_397_n N_X_M1004_s 0.00353387f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_425 N_B_c_413_n N_X_M1018_s 0.00362444f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_426 N_B_c_413_n N_X_c_1017_n 0.00892623f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_427 N_B_c_387_n N_X_c_1017_n 0.00618698f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_428 N_B_M1003_g N_X_c_1000_n 0.00895879f $X=6.785 $Y=0.74 $X2=0 $Y2=0
cc_429 N_B_c_386_n N_X_c_1000_n 0.010549f $X=5.89 $Y=1.78 $X2=0 $Y2=0
cc_430 N_B_c_387_n N_X_c_1000_n 0.065983f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_431 N_B_c_391_n N_X_c_1034_n 7.72218e-19 $X=6.795 $Y=1.765 $X2=0 $Y2=0
cc_432 N_B_c_391_n N_X_c_1008_n 0.0106815f $X=6.795 $Y=1.765 $X2=0 $Y2=0
cc_433 N_B_c_392_n N_X_c_1008_n 0.0107319f $X=7.245 $Y=1.765 $X2=0 $Y2=0
cc_434 N_B_c_393_n N_X_c_1008_n 0.0107319f $X=7.695 $Y=1.765 $X2=0 $Y2=0
cc_435 N_B_c_382_n N_X_c_1008_n 0.00262918f $X=8.145 $Y=1.35 $X2=0 $Y2=0
cc_436 N_B_c_395_n N_X_c_1008_n 0.0136266f $X=8.145 $Y=1.765 $X2=0 $Y2=0
cc_437 N_B_c_387_n N_X_c_1008_n 0.126413f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_438 N_B_c_413_n N_X_c_1037_n 0.0148765f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_439 N_B_c_387_n N_X_c_1037_n 0.011938f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_440 N_B_M1003_g N_X_c_1040_n 0.00659181f $X=6.785 $Y=0.74 $X2=0 $Y2=0
cc_441 N_B_c_378_n N_X_c_1040_n 5.72926e-19 $X=7.14 $Y=0.22 $X2=0 $Y2=0
cc_442 N_B_M1007_g N_X_c_1040_n 0.00674159f $X=7.215 $Y=0.74 $X2=0 $Y2=0
cc_443 N_B_M1014_g N_X_c_1040_n 7.30686e-19 $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_444 N_B_M1007_g N_X_c_1002_n 0.0093986f $X=7.215 $Y=0.74 $X2=0 $Y2=0
cc_445 N_B_M1014_g N_X_c_1002_n 0.0124803f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_446 N_B_c_382_n N_X_c_1002_n 0.00816204f $X=8.145 $Y=1.35 $X2=0 $Y2=0
cc_447 N_B_c_387_n N_X_c_1002_n 0.0510605f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_448 N_B_c_382_n N_X_c_1003_n 5.79778e-19 $X=8.145 $Y=1.35 $X2=0 $Y2=0
cc_449 N_B_M1019_g N_X_c_1003_n 0.0151483f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_450 N_B_c_387_n N_X_c_1003_n 0.0111136f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_451 N_B_c_382_n N_X_c_1004_n 0.0112809f $X=8.145 $Y=1.35 $X2=0 $Y2=0
cc_452 N_B_M1019_g N_X_c_1004_n 0.00614193f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_453 N_B_c_395_n N_X_c_1004_n 0.00646353f $X=8.145 $Y=1.765 $X2=0 $Y2=0
cc_454 N_B_c_387_n N_X_c_1004_n 0.034159f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_455 N_B_c_397_n N_X_c_1076_n 0.0168755f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_456 N_B_c_375_n N_X_c_1006_n 8.06164e-19 $X=6.795 $Y=1.275 $X2=0 $Y2=0
cc_457 N_B_M1003_g N_X_c_1006_n 0.00277633f $X=6.785 $Y=0.74 $X2=0 $Y2=0
cc_458 N_B_M1007_g N_X_c_1006_n 0.00269795f $X=7.215 $Y=0.74 $X2=0 $Y2=0
cc_459 N_B_c_387_n N_X_c_1006_n 0.0289344f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_460 N_B_c_382_n N_X_c_1007_n 0.00231547f $X=8.145 $Y=1.35 $X2=0 $Y2=0
cc_461 N_B_c_387_n N_X_c_1007_n 0.0144276f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_462 N_B_c_397_n N_X_c_1083_n 0.00641807f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_463 N_B_c_413_n N_X_c_1083_n 0.116551f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_464 N_B_c_428_n N_X_c_1083_n 0.0110991f $X=3.57 $Y=1.935 $X2=0 $Y2=0
cc_465 N_B_M1026_g N_VGND_c_1172_n 0.00203574f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_466 N_B_c_379_n N_VGND_c_1175_n 0.00170967f $X=6.86 $Y=0.22 $X2=0 $Y2=0
cc_467 N_B_M1017_g N_VGND_c_1176_n 0.0014541f $X=1.745 $Y=0.86 $X2=0 $Y2=0
cc_468 N_B_M1017_g N_VGND_c_1180_n 0.00376411f $X=1.745 $Y=0.86 $X2=0 $Y2=0
cc_469 N_B_M1026_g N_VGND_c_1180_n 0.00376411f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_470 N_B_c_379_n N_VGND_c_1183_n 0.0124522f $X=6.86 $Y=0.22 $X2=0 $Y2=0
cc_471 N_B_M1014_g N_VGND_c_1183_n 0.00278247f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_472 N_B_M1019_g N_VGND_c_1183_n 0.00278247f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_473 N_B_M1017_g N_VGND_c_1184_n 0.00508379f $X=1.745 $Y=0.86 $X2=0 $Y2=0
cc_474 N_B_M1026_g N_VGND_c_1184_n 0.00508379f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_475 N_B_c_378_n N_VGND_c_1184_n 0.0121953f $X=7.14 $Y=0.22 $X2=0 $Y2=0
cc_476 N_B_c_379_n N_VGND_c_1184_n 0.00536641f $X=6.86 $Y=0.22 $X2=0 $Y2=0
cc_477 N_B_M1014_g N_VGND_c_1184_n 0.00354085f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_478 N_B_M1019_g N_VGND_c_1184_n 0.00357084f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_479 N_B_M1003_g N_A_877_74#_c_1292_n 0.00852441f $X=6.785 $Y=0.74 $X2=0 $Y2=0
cc_480 N_B_c_378_n N_A_877_74#_c_1292_n 0.00709642f $X=7.14 $Y=0.22 $X2=0 $Y2=0
cc_481 N_B_c_379_n N_A_877_74#_c_1292_n 0.00216415f $X=6.86 $Y=0.22 $X2=0 $Y2=0
cc_482 N_B_M1007_g N_A_877_74#_c_1292_n 0.0088595f $X=7.215 $Y=0.74 $X2=0 $Y2=0
cc_483 N_B_M1014_g N_A_877_74#_c_1316_n 0.00646522f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_484 N_B_M1019_g N_A_877_74#_c_1316_n 5.7278e-19 $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_485 N_B_M1014_g N_A_877_74#_c_1294_n 0.00792642f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_486 N_B_M1019_g N_A_877_74#_c_1294_n 0.0118796f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_487 N_B_M1014_g N_A_877_74#_c_1295_n 5.7278e-19 $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_488 N_B_M1019_g N_A_877_74#_c_1295_n 0.00690717f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_489 N_B_M1014_g N_A_877_74#_c_1298_n 0.00294698f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_490 N_A_160_98#_c_583_n N_A_36_392#_c_719_n 0.0122194f $X=1.725 $Y=2.105
+ $X2=0 $Y2=0
cc_491 N_A_160_98#_c_583_n N_A_36_392#_c_734_n 0.0423287f $X=1.725 $Y=2.105
+ $X2=0 $Y2=0
cc_492 N_A_160_98#_M1001_d N_A_36_392#_c_721_n 0.00222494f $X=1.575 $Y=1.96
+ $X2=0 $Y2=0
cc_493 N_A_160_98#_c_587_n N_A_36_392#_c_721_n 5.7057e-19 $X=2.925 $Y=1.765
+ $X2=0 $Y2=0
cc_494 N_A_160_98#_c_583_n N_A_36_392#_c_721_n 0.0144323f $X=1.725 $Y=2.105
+ $X2=0 $Y2=0
cc_495 N_A_160_98#_c_583_n N_A_36_392#_c_723_n 0.0365429f $X=1.725 $Y=2.105
+ $X2=0 $Y2=0
cc_496 N_A_160_98#_c_587_n N_VPWR_c_768_n 0.00278271f $X=2.925 $Y=1.765 $X2=0
+ $Y2=0
cc_497 N_A_160_98#_c_588_n N_VPWR_c_768_n 0.00278271f $X=3.375 $Y=1.765 $X2=0
+ $Y2=0
cc_498 N_A_160_98#_c_589_n N_VPWR_c_768_n 0.00278271f $X=3.825 $Y=1.765 $X2=0
+ $Y2=0
cc_499 N_A_160_98#_c_592_n N_VPWR_c_768_n 0.00278271f $X=4.275 $Y=1.765 $X2=0
+ $Y2=0
cc_500 N_A_160_98#_c_587_n N_VPWR_c_764_n 0.00358624f $X=2.925 $Y=1.765 $X2=0
+ $Y2=0
cc_501 N_A_160_98#_c_588_n N_VPWR_c_764_n 0.00353823f $X=3.375 $Y=1.765 $X2=0
+ $Y2=0
cc_502 N_A_160_98#_c_589_n N_VPWR_c_764_n 0.00353823f $X=3.825 $Y=1.765 $X2=0
+ $Y2=0
cc_503 N_A_160_98#_c_592_n N_VPWR_c_764_n 0.00353907f $X=4.275 $Y=1.765 $X2=0
+ $Y2=0
cc_504 N_A_160_98#_c_587_n N_A_514_368#_c_881_n 0.00679598f $X=2.925 $Y=1.765
+ $X2=0 $Y2=0
cc_505 N_A_160_98#_c_587_n N_A_514_368#_c_882_n 0.0137046f $X=2.925 $Y=1.765
+ $X2=0 $Y2=0
cc_506 N_A_160_98#_c_588_n N_A_514_368#_c_882_n 0.00999576f $X=3.375 $Y=1.765
+ $X2=0 $Y2=0
cc_507 N_A_160_98#_c_589_n N_A_514_368#_c_884_n 0.00995895f $X=3.825 $Y=1.765
+ $X2=0 $Y2=0
cc_508 N_A_160_98#_c_592_n N_A_514_368#_c_884_n 0.00918039f $X=4.275 $Y=1.765
+ $X2=0 $Y2=0
cc_509 N_A_160_98#_c_592_n N_A_514_368#_c_887_n 2.20491e-19 $X=4.275 $Y=1.765
+ $X2=0 $Y2=0
cc_510 N_A_160_98#_c_579_n N_X_c_998_n 0.0108146f $X=3.59 $Y=1.35 $X2=0 $Y2=0
cc_511 N_A_160_98#_c_580_n N_X_c_998_n 5.72677e-19 $X=4.185 $Y=1.605 $X2=0 $Y2=0
cc_512 N_A_160_98#_c_579_n N_X_c_999_n 0.00409433f $X=3.59 $Y=1.35 $X2=0 $Y2=0
cc_513 N_A_160_98#_c_592_n N_X_c_1017_n 0.00916137f $X=4.275 $Y=1.765 $X2=0
+ $Y2=0
cc_514 N_A_160_98#_c_582_n N_X_c_1000_n 4.06994e-19 $X=4.275 $Y=1.605 $X2=0
+ $Y2=0
cc_515 N_A_160_98#_c_579_n N_X_c_1001_n 0.00102704f $X=3.59 $Y=1.35 $X2=0 $Y2=0
cc_516 N_A_160_98#_c_580_n N_X_c_1001_n 8.51159e-19 $X=4.185 $Y=1.605 $X2=0
+ $Y2=0
cc_517 N_A_160_98#_c_587_n N_X_c_1076_n 0.00622519f $X=2.925 $Y=1.765 $X2=0
+ $Y2=0
cc_518 N_A_160_98#_c_588_n N_X_c_1076_n 0.00688021f $X=3.375 $Y=1.765 $X2=0
+ $Y2=0
cc_519 N_A_160_98#_c_589_n N_X_c_1076_n 0.00102753f $X=3.825 $Y=1.765 $X2=0
+ $Y2=0
cc_520 N_A_160_98#_c_578_n N_X_c_1005_n 0.00391079f $X=2.875 $Y=1.35 $X2=0 $Y2=0
cc_521 N_A_160_98#_c_579_n N_X_c_1005_n 0.00967015f $X=3.59 $Y=1.35 $X2=0 $Y2=0
cc_522 N_A_160_98#_c_588_n N_X_c_1083_n 0.0107397f $X=3.375 $Y=1.765 $X2=0 $Y2=0
cc_523 N_A_160_98#_c_589_n N_X_c_1083_n 0.00921244f $X=3.825 $Y=1.765 $X2=0
+ $Y2=0
cc_524 N_A_160_98#_c_581_n N_X_c_1083_n 2.25987e-19 $X=3.915 $Y=1.605 $X2=0
+ $Y2=0
cc_525 N_A_160_98#_c_588_n N_X_c_1044_n 4.92205e-19 $X=3.375 $Y=1.765 $X2=0
+ $Y2=0
cc_526 N_A_160_98#_c_589_n N_X_c_1044_n 0.00548579f $X=3.825 $Y=1.765 $X2=0
+ $Y2=0
cc_527 N_A_160_98#_c_592_n N_X_c_1044_n 0.00553331f $X=4.275 $Y=1.765 $X2=0
+ $Y2=0
cc_528 N_A_160_98#_c_613_n N_VGND_M1016_s 0.0113915f $X=1.56 $Y=1.065 $X2=0
+ $Y2=0
cc_529 N_A_160_98#_c_583_n N_VGND_M1016_s 4.81637e-19 $X=1.725 $Y=2.105 $X2=0
+ $Y2=0
cc_530 N_A_160_98#_c_633_n N_VGND_M1016_s 5.87954e-19 $X=1.685 $Y=1.065 $X2=0
+ $Y2=0
cc_531 N_A_160_98#_c_621_n N_VGND_M1026_s 0.00947801f $X=2.53 $Y=1.065 $X2=0
+ $Y2=0
cc_532 N_A_160_98#_c_584_n N_VGND_M1026_s 8.87448e-19 $X=2.615 $Y=1.36 $X2=0
+ $Y2=0
cc_533 N_A_160_98#_c_578_n N_VGND_c_1172_n 0.00203574f $X=2.875 $Y=1.35 $X2=0
+ $Y2=0
cc_534 N_A_160_98#_c_579_n N_VGND_c_1173_n 0.00559625f $X=3.59 $Y=1.35 $X2=0
+ $Y2=0
cc_535 N_A_160_98#_c_578_n N_VGND_c_1178_n 0.00376367f $X=2.875 $Y=1.35 $X2=0
+ $Y2=0
cc_536 N_A_160_98#_c_579_n N_VGND_c_1178_n 0.00380789f $X=3.59 $Y=1.35 $X2=0
+ $Y2=0
cc_537 N_A_160_98#_c_578_n N_VGND_c_1184_n 0.00508379f $X=2.875 $Y=1.35 $X2=0
+ $Y2=0
cc_538 N_A_160_98#_c_579_n N_VGND_c_1184_n 0.00508379f $X=3.59 $Y=1.35 $X2=0
+ $Y2=0
cc_539 N_A_36_392#_c_719_n N_VPWR_M1021_s 0.00275645f $X=1.11 $Y=2.005 $X2=-0.19
+ $Y2=1.66
cc_540 N_A_36_392#_c_718_n N_VPWR_c_765_n 0.0483063f $X=0.325 $Y=2.105 $X2=0
+ $Y2=0
cc_541 N_A_36_392#_c_719_n N_VPWR_c_765_n 0.0184684f $X=1.11 $Y=2.005 $X2=0
+ $Y2=0
cc_542 N_A_36_392#_c_722_n N_VPWR_c_765_n 0.0117278f $X=1.36 $Y=2.99 $X2=0 $Y2=0
cc_543 N_A_36_392#_c_721_n N_VPWR_c_768_n 0.0645908f $X=2.01 $Y=2.99 $X2=0 $Y2=0
cc_544 N_A_36_392#_c_722_n N_VPWR_c_768_n 0.017869f $X=1.36 $Y=2.99 $X2=0 $Y2=0
cc_545 N_A_36_392#_c_718_n N_VPWR_c_764_n 0.0120466f $X=0.325 $Y=2.105 $X2=0
+ $Y2=0
cc_546 N_A_36_392#_c_721_n N_VPWR_c_764_n 0.0358952f $X=2.01 $Y=2.99 $X2=0 $Y2=0
cc_547 N_A_36_392#_c_722_n N_VPWR_c_764_n 0.00965079f $X=1.36 $Y=2.99 $X2=0
+ $Y2=0
cc_548 N_A_36_392#_c_718_n N_VPWR_c_774_n 0.0145938f $X=0.325 $Y=2.105 $X2=0
+ $Y2=0
cc_549 N_A_36_392#_c_723_n N_A_514_368#_c_881_n 0.0528784f $X=2.175 $Y=2.355
+ $X2=0 $Y2=0
cc_550 N_A_36_392#_c_721_n N_A_514_368#_c_883_n 0.0144477f $X=2.01 $Y=2.99 $X2=0
+ $Y2=0
cc_551 N_A_36_392#_c_720_n N_VGND_c_1171_n 0.00657381f $X=0.49 $Y=2.005 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_768_n N_A_514_368#_c_882_n 0.0460938f $X=4.855 $Y=3.33 $X2=0
+ $Y2=0
cc_553 N_VPWR_c_764_n N_A_514_368#_c_882_n 0.0260732f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_554 N_VPWR_c_768_n N_A_514_368#_c_883_n 0.0179217f $X=4.855 $Y=3.33 $X2=0
+ $Y2=0
cc_555 N_VPWR_c_764_n N_A_514_368#_c_883_n 0.00971942f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_768_n N_A_514_368#_c_884_n 0.0461229f $X=4.855 $Y=3.33 $X2=0
+ $Y2=0
cc_557 N_VPWR_c_764_n N_A_514_368#_c_884_n 0.0260772f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_558 N_VPWR_M1025_s N_A_514_368#_c_891_n 0.00716177f $X=5.84 $Y=1.84 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_769_n N_A_514_368#_c_891_n 0.00241722f $X=5.89 $Y=3.33 $X2=0
+ $Y2=0
cc_560 N_VPWR_c_770_n N_A_514_368#_c_891_n 0.00395989f $X=6.855 $Y=3.33 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_764_n N_A_514_368#_c_891_n 0.0115059f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_562 N_VPWR_c_776_n N_A_514_368#_c_891_n 0.0238912f $X=6.055 $Y=3.05 $X2=0
+ $Y2=0
cc_563 N_VPWR_c_766_n N_A_514_368#_c_885_n 0.02367f $X=7.02 $Y=2.805 $X2=0 $Y2=0
cc_564 N_VPWR_c_770_n N_A_514_368#_c_885_n 0.00759366f $X=6.855 $Y=3.33 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_764_n N_A_514_368#_c_885_n 0.00628181f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_776_n N_A_514_368#_c_885_n 8.74655e-19 $X=6.055 $Y=3.05 $X2=0
+ $Y2=0
cc_567 N_VPWR_M1002_d N_A_514_368#_c_911_n 0.00420698f $X=6.87 $Y=1.84 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_766_n N_A_514_368#_c_911_n 0.0154248f $X=7.02 $Y=2.805 $X2=0
+ $Y2=0
cc_569 N_VPWR_M1015_d N_A_514_368#_c_913_n 0.00428955f $X=7.77 $Y=1.84 $X2=0
+ $Y2=0
cc_570 N_VPWR_c_767_n N_A_514_368#_c_913_n 0.0136682f $X=7.92 $Y=2.805 $X2=0
+ $Y2=0
cc_571 N_VPWR_c_768_n N_A_514_368#_c_886_n 0.0118207f $X=4.855 $Y=3.33 $X2=0
+ $Y2=0
cc_572 N_VPWR_c_764_n N_A_514_368#_c_886_n 0.00654074f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_573 N_VPWR_c_768_n N_A_514_368#_c_887_n 0.0171913f $X=4.855 $Y=3.33 $X2=0
+ $Y2=0
cc_574 N_VPWR_c_764_n N_A_514_368#_c_887_n 0.00947661f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_575 N_VPWR_c_775_n N_A_514_368#_c_887_n 0.00784976f $X=5.02 $Y=3.05 $X2=0
+ $Y2=0
cc_576 N_VPWR_M1005_s N_A_514_368#_c_896_n 0.00747361f $X=4.8 $Y=1.84 $X2=0
+ $Y2=0
cc_577 N_VPWR_c_768_n N_A_514_368#_c_896_n 0.00352633f $X=4.855 $Y=3.33 $X2=0
+ $Y2=0
cc_578 N_VPWR_c_769_n N_A_514_368#_c_896_n 0.00351825f $X=5.89 $Y=3.33 $X2=0
+ $Y2=0
cc_579 N_VPWR_c_764_n N_A_514_368#_c_896_n 0.0122633f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_580 N_VPWR_c_775_n N_A_514_368#_c_896_n 0.0241887f $X=5.02 $Y=3.05 $X2=0
+ $Y2=0
cc_581 N_VPWR_c_769_n N_A_514_368#_c_888_n 0.0139149f $X=5.89 $Y=3.33 $X2=0
+ $Y2=0
cc_582 N_VPWR_c_764_n N_A_514_368#_c_888_n 0.0117794f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_583 N_VPWR_c_775_n N_A_514_368#_c_888_n 0.00102355f $X=5.02 $Y=3.05 $X2=0
+ $Y2=0
cc_584 N_VPWR_c_776_n N_A_514_368#_c_888_n 0.00104431f $X=6.055 $Y=3.05 $X2=0
+ $Y2=0
cc_585 N_VPWR_c_766_n N_A_514_368#_c_889_n 0.0234974f $X=7.02 $Y=2.805 $X2=0
+ $Y2=0
cc_586 N_VPWR_c_767_n N_A_514_368#_c_889_n 0.0228252f $X=7.92 $Y=2.805 $X2=0
+ $Y2=0
cc_587 N_VPWR_c_771_n N_A_514_368#_c_889_n 0.0145674f $X=7.835 $Y=3.33 $X2=0
+ $Y2=0
cc_588 N_VPWR_c_764_n N_A_514_368#_c_889_n 0.0119851f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_589 N_VPWR_c_767_n N_A_514_368#_c_890_n 0.0228252f $X=7.92 $Y=2.805 $X2=0
+ $Y2=0
cc_590 N_VPWR_c_772_n N_A_514_368#_c_890_n 0.0146094f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_591 N_VPWR_c_764_n N_A_514_368#_c_890_n 0.0120527f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_592 N_VPWR_M1005_s N_X_c_1017_n 0.00739825f $X=4.8 $Y=1.84 $X2=0 $Y2=0
cc_593 N_VPWR_M1025_s N_X_c_1017_n 0.00752668f $X=5.84 $Y=1.84 $X2=0 $Y2=0
cc_594 N_VPWR_M1025_s N_X_c_1034_n 0.00210547f $X=5.84 $Y=1.84 $X2=0 $Y2=0
cc_595 N_VPWR_M1002_d N_X_c_1008_n 0.00396407f $X=6.87 $Y=1.84 $X2=0 $Y2=0
cc_596 N_VPWR_M1015_d N_X_c_1008_n 0.00359847f $X=7.77 $Y=1.84 $X2=0 $Y2=0
cc_597 N_VPWR_M1025_s N_X_c_1037_n 0.00221099f $X=5.84 $Y=1.84 $X2=0 $Y2=0
cc_598 N_A_514_368#_c_882_n N_X_M1004_s 0.00197722f $X=3.515 $Y=2.99 $X2=0 $Y2=0
cc_599 N_A_514_368#_c_884_n N_X_M1018_s 0.00198204f $X=4.415 $Y=2.99 $X2=0 $Y2=0
cc_600 N_A_514_368#_M1029_d N_X_c_1017_n 0.00400018f $X=4.35 $Y=1.84 $X2=0 $Y2=0
cc_601 N_A_514_368#_M1013_d N_X_c_1017_n 0.00379665f $X=5.39 $Y=1.84 $X2=0 $Y2=0
cc_602 N_A_514_368#_c_884_n N_X_c_1017_n 0.00441078f $X=4.415 $Y=2.99 $X2=0
+ $Y2=0
cc_603 N_A_514_368#_c_891_n N_X_c_1017_n 0.00874461f $X=6.485 $Y=2.71 $X2=0
+ $Y2=0
cc_604 N_A_514_368#_c_975_p N_X_c_1017_n 0.0144215f $X=6.57 $Y=2.46 $X2=0 $Y2=0
cc_605 N_A_514_368#_c_887_n N_X_c_1017_n 0.0149196f $X=4.54 $Y=2.71 $X2=0 $Y2=0
cc_606 N_A_514_368#_c_896_n N_X_c_1017_n 0.0858075f $X=5.375 $Y=2.802 $X2=0
+ $Y2=0
cc_607 N_A_514_368#_M1028_d N_X_c_1008_n 0.00401969f $X=6.42 $Y=1.84 $X2=0 $Y2=0
cc_608 N_A_514_368#_M1011_s N_X_c_1008_n 0.00359365f $X=7.32 $Y=1.84 $X2=0 $Y2=0
cc_609 N_A_514_368#_M1022_s N_X_c_1008_n 0.0132967f $X=8.22 $Y=1.84 $X2=0 $Y2=0
cc_610 N_A_514_368#_c_891_n N_X_c_1008_n 0.00316891f $X=6.485 $Y=2.71 $X2=0
+ $Y2=0
cc_611 N_A_514_368#_c_975_p N_X_c_1008_n 0.0138475f $X=6.57 $Y=2.46 $X2=0 $Y2=0
cc_612 N_A_514_368#_c_911_n N_X_c_1008_n 0.0333042f $X=7.305 $Y=2.375 $X2=0
+ $Y2=0
cc_613 N_A_514_368#_c_913_n N_X_c_1008_n 0.0317427f $X=8.205 $Y=2.375 $X2=0
+ $Y2=0
cc_614 N_A_514_368#_c_889_n N_X_c_1008_n 0.0173542f $X=7.47 $Y=2.455 $X2=0 $Y2=0
cc_615 N_A_514_368#_c_890_n N_X_c_1008_n 0.0209985f $X=8.37 $Y=2.455 $X2=0 $Y2=0
cc_616 N_A_514_368#_M1022_s N_X_c_1004_n 0.00601094f $X=8.22 $Y=1.84 $X2=0 $Y2=0
cc_617 N_A_514_368#_c_881_n N_X_c_1076_n 0.0365429f $X=2.7 $Y=2.355 $X2=0 $Y2=0
cc_618 N_A_514_368#_c_882_n N_X_c_1076_n 0.0158076f $X=3.515 $Y=2.99 $X2=0 $Y2=0
cc_619 N_A_514_368#_c_990_p N_X_c_1076_n 0.00716505f $X=3.6 $Y=2.8 $X2=0 $Y2=0
cc_620 N_A_514_368#_M1012_d N_X_c_1083_n 0.00386063f $X=3.45 $Y=1.84 $X2=0 $Y2=0
cc_621 N_A_514_368#_c_882_n N_X_c_1083_n 0.00440848f $X=3.515 $Y=2.99 $X2=0
+ $Y2=0
cc_622 N_A_514_368#_c_990_p N_X_c_1083_n 0.0132204f $X=3.6 $Y=2.8 $X2=0 $Y2=0
cc_623 N_A_514_368#_c_884_n N_X_c_1083_n 0.00439308f $X=4.415 $Y=2.99 $X2=0
+ $Y2=0
cc_624 N_A_514_368#_c_990_p N_X_c_1044_n 0.00713066f $X=3.6 $Y=2.8 $X2=0 $Y2=0
cc_625 N_A_514_368#_c_884_n N_X_c_1044_n 0.0157037f $X=4.415 $Y=2.99 $X2=0 $Y2=0
cc_626 N_A_514_368#_c_887_n N_X_c_1044_n 0.00734009f $X=4.54 $Y=2.71 $X2=0 $Y2=0
cc_627 N_X_c_998_n N_VGND_M1027_d 0.011365f $X=4.105 $Y=0.765 $X2=0 $Y2=0
cc_628 N_X_c_999_n N_VGND_M1027_d 0.00238572f $X=4.19 $Y=1.01 $X2=0 $Y2=0
cc_629 N_X_c_1001_n N_VGND_M1027_d 0.00189155f $X=4.275 $Y=1.095 $X2=0 $Y2=0
cc_630 N_X_c_1000_n N_VGND_M1009_d 0.00391227f $X=6.835 $Y=1.095 $X2=0 $Y2=0
cc_631 N_X_c_1000_n N_VGND_M1020_d 0.00391227f $X=6.835 $Y=1.095 $X2=0 $Y2=0
cc_632 N_X_c_998_n N_VGND_c_1173_n 0.0320467f $X=4.105 $Y=0.765 $X2=0 $Y2=0
cc_633 N_X_c_1005_n N_VGND_c_1173_n 0.00221964f $X=3.375 $Y=0.66 $X2=0 $Y2=0
cc_634 N_X_c_998_n N_VGND_c_1178_n 0.0023127f $X=4.105 $Y=0.765 $X2=0 $Y2=0
cc_635 N_X_c_1005_n N_VGND_c_1178_n 0.00937878f $X=3.375 $Y=0.66 $X2=0 $Y2=0
cc_636 N_X_c_998_n N_VGND_c_1181_n 0.00251932f $X=4.105 $Y=0.765 $X2=0 $Y2=0
cc_637 N_X_c_998_n N_VGND_c_1184_n 0.0106811f $X=4.105 $Y=0.765 $X2=0 $Y2=0
cc_638 N_X_c_1005_n N_VGND_c_1184_n 0.0109286f $X=3.375 $Y=0.66 $X2=0 $Y2=0
cc_639 N_X_c_1000_n N_A_877_74#_M1009_s 0.00463994f $X=6.835 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_640 N_X_c_1000_n N_A_877_74#_M1010_s 0.00176891f $X=6.835 $Y=1.095 $X2=0
+ $Y2=0
cc_641 N_X_c_1000_n N_A_877_74#_M1024_s 0.00176461f $X=6.835 $Y=1.095 $X2=0
+ $Y2=0
cc_642 N_X_c_1002_n N_A_877_74#_M1007_s 0.00250873f $X=7.845 $Y=1.095 $X2=0
+ $Y2=0
cc_643 N_X_c_1003_n N_A_877_74#_M1019_s 0.00757941f $X=8.335 $Y=1.095 $X2=0
+ $Y2=0
cc_644 N_X_c_1000_n N_A_877_74#_c_1301_n 0.0151804f $X=6.835 $Y=1.095 $X2=0
+ $Y2=0
cc_645 N_X_M1003_d N_A_877_74#_c_1292_n 0.00176461f $X=6.86 $Y=0.37 $X2=0 $Y2=0
cc_646 N_X_c_1000_n N_A_877_74#_c_1292_n 0.00304353f $X=6.835 $Y=1.095 $X2=0
+ $Y2=0
cc_647 N_X_c_1040_n N_A_877_74#_c_1292_n 0.0157964f $X=7 $Y=0.76 $X2=0 $Y2=0
cc_648 N_X_c_1002_n N_A_877_74#_c_1292_n 0.00304353f $X=7.845 $Y=1.095 $X2=0
+ $Y2=0
cc_649 N_X_c_1002_n N_A_877_74#_c_1316_n 0.020731f $X=7.845 $Y=1.095 $X2=0 $Y2=0
cc_650 N_X_M1014_d N_A_877_74#_c_1294_n 0.00176461f $X=7.79 $Y=0.37 $X2=0 $Y2=0
cc_651 N_X_c_1002_n N_A_877_74#_c_1294_n 0.00304353f $X=7.845 $Y=1.095 $X2=0
+ $Y2=0
cc_652 N_X_c_1164_p N_A_877_74#_c_1294_n 0.0124895f $X=7.93 $Y=0.805 $X2=0 $Y2=0
cc_653 N_X_c_1003_n N_A_877_74#_c_1294_n 0.00304353f $X=8.335 $Y=1.095 $X2=0
+ $Y2=0
cc_654 N_X_c_1003_n N_A_877_74#_c_1295_n 0.0215474f $X=8.335 $Y=1.095 $X2=0
+ $Y2=0
cc_655 N_X_c_998_n N_A_877_74#_c_1296_n 0.0147083f $X=4.105 $Y=0.765 $X2=0 $Y2=0
cc_656 N_X_c_1000_n N_A_877_74#_c_1296_n 0.0150829f $X=6.835 $Y=1.095 $X2=0
+ $Y2=0
cc_657 N_X_c_1000_n N_A_877_74#_c_1306_n 0.0978095f $X=6.835 $Y=1.095 $X2=0
+ $Y2=0
cc_658 N_VGND_M1020_d N_A_877_74#_c_1299_n 0.00726893f $X=5.84 $Y=0.37 $X2=0
+ $Y2=0
cc_659 N_VGND_c_1175_n N_A_877_74#_c_1299_n 0.0251188f $X=6.06 $Y=0.335 $X2=0
+ $Y2=0
cc_660 N_VGND_c_1182_n N_A_877_74#_c_1299_n 0.00236055f $X=5.895 $Y=0 $X2=0
+ $Y2=0
cc_661 N_VGND_c_1183_n N_A_877_74#_c_1299_n 0.00236055f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_662 N_VGND_c_1184_n N_A_877_74#_c_1299_n 0.0102106f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_663 N_VGND_c_1183_n N_A_877_74#_c_1292_n 0.0420053f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_664 N_VGND_c_1184_n N_A_877_74#_c_1292_n 0.022853f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_665 N_VGND_c_1175_n N_A_877_74#_c_1293_n 0.0114117f $X=6.06 $Y=0.335 $X2=0
+ $Y2=0
cc_666 N_VGND_c_1183_n N_A_877_74#_c_1293_n 0.0176331f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_667 N_VGND_c_1184_n N_A_877_74#_c_1293_n 0.00956698f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_668 N_VGND_c_1183_n N_A_877_74#_c_1294_n 0.0566663f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_669 N_VGND_c_1184_n N_A_877_74#_c_1294_n 0.0314476f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_670 N_VGND_c_1173_n N_A_877_74#_c_1296_n 0.00853811f $X=3.925 $Y=0.345 $X2=0
+ $Y2=0
cc_671 N_VGND_c_1174_n N_A_877_74#_c_1296_n 0.00591149f $X=5.04 $Y=0.335 $X2=0
+ $Y2=0
cc_672 N_VGND_c_1181_n N_A_877_74#_c_1296_n 0.0107387f $X=4.875 $Y=0 $X2=0 $Y2=0
cc_673 N_VGND_c_1184_n N_A_877_74#_c_1296_n 0.00894442f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_674 N_VGND_M1009_d N_A_877_74#_c_1306_n 0.00726893f $X=4.82 $Y=0.37 $X2=0
+ $Y2=0
cc_675 N_VGND_c_1174_n N_A_877_74#_c_1306_n 0.0251188f $X=5.04 $Y=0.335 $X2=0
+ $Y2=0
cc_676 N_VGND_c_1181_n N_A_877_74#_c_1306_n 0.00236055f $X=4.875 $Y=0 $X2=0
+ $Y2=0
cc_677 N_VGND_c_1182_n N_A_877_74#_c_1306_n 0.00236055f $X=5.895 $Y=0 $X2=0
+ $Y2=0
cc_678 N_VGND_c_1184_n N_A_877_74#_c_1306_n 0.0102106f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_679 N_VGND_c_1174_n N_A_877_74#_c_1297_n 0.0060913f $X=5.04 $Y=0.335 $X2=0
+ $Y2=0
cc_680 N_VGND_c_1175_n N_A_877_74#_c_1297_n 0.0060913f $X=6.06 $Y=0.335 $X2=0
+ $Y2=0
cc_681 N_VGND_c_1182_n N_A_877_74#_c_1297_n 0.0141766f $X=5.895 $Y=0 $X2=0 $Y2=0
cc_682 N_VGND_c_1184_n N_A_877_74#_c_1297_n 0.0118057f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_683 N_VGND_c_1183_n N_A_877_74#_c_1298_n 0.0233048f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_684 N_VGND_c_1184_n N_A_877_74#_c_1298_n 0.0126653f $X=8.4 $Y=0 $X2=0 $Y2=0
