* File: sky130_fd_sc_ls__o21bai_1.pex.spice
* Created: Wed Sep  2 11:18:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O21BAI_1%B1_N 3 5 7 8 12
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.4
+ $Y=1.615 $X2=0.4 $Y2=1.615
r33 8 12 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.24 $Y=1.615 $X2=0.4
+ $Y2=1.615
r34 5 11 87.63 $w=2.63e-07 $l=4.77389e-07 $layer=POLY_cond $X=0.525 $Y=2.045
+ $X2=0.425 $Y2=1.615
r35 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.525 $Y=2.045
+ $X2=0.525 $Y2=2.54
r36 1 11 39.0634 $w=2.63e-07 $l=1.94808e-07 $layer=POLY_cond $X=0.49 $Y=1.45
+ $X2=0.425 $Y2=1.615
r37 1 3 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=0.49 $Y=1.45 $X2=0.49
+ $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__O21BAI_1%A_27_74# 1 2 7 10 11 13 16 18 21 25 27 28
+ 29 30 31 32 37
r78 36 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.97 $Y=1.465 $X2=0.97
+ $Y2=1.375
r79 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.465 $X2=0.97 $Y2=1.465
r80 31 35 8.96496 $w=3.09e-07 $l=2.13014e-07 $layer=LI1_cond $X=0.83 $Y=1.63
+ $X2=0.94 $Y2=1.465
r81 31 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.83 $Y=1.63 $X2=0.83
+ $Y2=1.95
r82 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.745 $Y=2.035
+ $X2=0.83 $Y2=1.95
r83 29 30 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.745 $Y=2.035
+ $X2=0.465 $Y2=2.035
r84 27 35 10.6602 $w=3.09e-07 $l=3.5433e-07 $layer=LI1_cond $X=0.745 $Y=1.195
+ $X2=0.94 $Y2=1.465
r85 27 28 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.745 $Y=1.195
+ $X2=0.36 $Y2=1.195
r86 23 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.3 $Y=2.12
+ $X2=0.465 $Y2=2.035
r87 23 25 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.3 $Y=2.12 $X2=0.3
+ $Y2=2.265
r88 19 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.235 $Y=1.11
+ $X2=0.36 $Y2=1.195
r89 19 21 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=0.235 $Y=1.11
+ $X2=0.235 $Y2=0.645
r90 14 18 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.465 $Y=1.3
+ $X2=1.45 $Y2=1.375
r91 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.465 $Y=1.3
+ $X2=1.465 $Y2=0.74
r92 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.45 $Y=1.765
+ $X2=1.45 $Y2=2.4
r93 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.45 $Y=1.675 $X2=1.45
+ $Y2=1.765
r94 9 18 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.45 $Y=1.45
+ $X2=1.45 $Y2=1.375
r95 9 10 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=1.45 $Y=1.45
+ $X2=1.45 $Y2=1.675
r96 8 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.135 $Y=1.375
+ $X2=0.97 $Y2=1.375
r97 7 18 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.36 $Y=1.375 $X2=1.45
+ $Y2=1.375
r98 7 8 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.36 $Y=1.375
+ $X2=1.135 $Y2=1.375
r99 2 25 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.155
+ $Y=2.12 $X2=0.3 $Y2=2.265
r100 1 21 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.275 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__O21BAI_1%A2 1 3 6 8 9 10 11 22
r40 20 22 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.16 $Y=1.63
+ $X2=2.16 $Y2=1.665
r41 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.915
+ $Y=1.465 $X2=1.915 $Y2=1.465
r42 10 11 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=2.405
+ $X2=2.16 $Y2=2.775
r43 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=2.035
+ $X2=2.16 $Y2=2.405
r44 8 20 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.16 $Y=1.465
+ $X2=2.16 $Y2=1.63
r45 8 19 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.16 $Y=1.465
+ $X2=1.915 $Y2=1.465
r46 8 9 17.2866 $w=2.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.16 $Y=1.69 $X2=2.16
+ $Y2=2.035
r47 8 22 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2.16 $Y=1.69 $X2=2.16
+ $Y2=1.665
r48 4 18 38.6549 $w=2.86e-07 $l=1.79374e-07 $layer=POLY_cond $X=1.945 $Y=1.3
+ $X2=1.915 $Y2=1.465
r49 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.945 $Y=1.3 $X2=1.945
+ $Y2=0.74
r50 1 18 61.4066 $w=2.86e-07 $l=3.07409e-07 $layer=POLY_cond $X=1.9 $Y=1.765
+ $X2=1.915 $Y2=1.465
r51 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.9 $Y=1.765 $X2=1.9
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O21BAI_1%A1 1 3 6 8 12
r24 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.465 $X2=2.61 $Y2=1.465
r25 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.61 $Y=1.665 $X2=2.61
+ $Y2=1.465
r26 4 11 39.5078 $w=3.96e-07 $l=2.26892e-07 $layer=POLY_cond $X=2.385 $Y=1.3
+ $X2=2.532 $Y2=1.465
r27 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.385 $Y=1.3 $X2=2.385
+ $Y2=0.74
r28 1 11 55.9396 $w=3.96e-07 $l=3.68239e-07 $layer=POLY_cond $X=2.38 $Y=1.765
+ $X2=2.532 $Y2=1.465
r29 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.38 $Y=1.765
+ $X2=2.38 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O21BAI_1%VPWR 1 2 9 11 13 17 19 24 30 34
r33 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r35 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 25 30 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=0.97 $Y2=3.33
r38 25 27 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 24 33 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.52 $Y=3.33 $X2=2.7
+ $Y2=3.33
r40 24 27 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.52 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 22 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r42 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 19 30 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.97 $Y2=3.33
r44 19 21 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 17 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 17 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 13 16 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=2.645 $Y=2.115
+ $X2=2.645 $Y2=2.815
r48 11 33 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=2.645 $Y=3.245
+ $X2=2.7 $Y2=3.33
r49 11 16 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.645 $Y=3.245
+ $X2=2.645 $Y2=2.815
r50 7 30 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.97 $Y=3.245 $X2=0.97
+ $Y2=3.33
r51 7 9 14.103 $w=6.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.97 $Y=3.245 $X2=0.97
+ $Y2=2.455
r52 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.455
+ $Y=1.84 $X2=2.605 $Y2=2.815
r53 2 13 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.455
+ $Y=1.84 $X2=2.605 $Y2=2.115
r54 1 9 150 $w=1.7e-07 $l=6.87386e-07 $layer=licon1_PDIFF $count=4 $X=0.6
+ $Y=2.12 $X2=1.14 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__O21BAI_1%Y 1 2 9 13 14 15 16 23 32
r44 23 34 1.42082 $w=3.63e-07 $l=4.5e-08 $layer=LI1_cond $X=1.657 $Y=2.035
+ $X2=1.657 $Y2=1.99
r45 15 16 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.657 $Y=2.405
+ $X2=1.657 $Y2=2.775
r46 14 34 1.66283 $w=5.33e-07 $l=2e-08 $layer=LI1_cond $X=1.572 $Y=1.97
+ $X2=1.572 $Y2=1.99
r47 14 32 9.40076 $w=5.33e-07 $l=1.5e-07 $layer=LI1_cond $X=1.572 $Y=1.97
+ $X2=1.572 $Y2=1.82
r48 14 15 11.0508 $w=3.63e-07 $l=3.5e-07 $layer=LI1_cond $X=1.657 $Y=2.055
+ $X2=1.657 $Y2=2.405
r49 14 23 0.631476 $w=3.63e-07 $l=2e-08 $layer=LI1_cond $X=1.657 $Y=2.055
+ $X2=1.657 $Y2=2.035
r50 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.39 $Y=1.13 $X2=1.39
+ $Y2=1.82
r51 7 13 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=1.28 $Y=0.935
+ $X2=1.28 $Y2=1.13
r52 7 9 12.4109 $w=3.88e-07 $l=4.2e-07 $layer=LI1_cond $X=1.28 $Y=0.935 $X2=1.28
+ $Y2=0.515
r53 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.84 $X2=1.675 $Y2=1.985
r54 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.84 $X2=1.675 $Y2=2.815
r55 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.11
+ $Y=0.37 $X2=1.25 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O21BAI_1%VGND 1 2 9 13 15 17 22 29 30 33 36
r38 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r39 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r41 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 27 36 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.165
+ $Y2=0
r43 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.64
+ $Y2=0
r44 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r45 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r46 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.87 $Y=0 $X2=0.705
+ $Y2=0
r47 23 25 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.87 $Y=0 $X2=1.68
+ $Y2=0
r48 22 36 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.995 $Y=0 $X2=2.165
+ $Y2=0
r49 22 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=0 $X2=1.68
+ $Y2=0
r50 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r51 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r52 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.54 $Y=0 $X2=0.705
+ $Y2=0
r53 17 19 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.54 $Y=0 $X2=0.24
+ $Y2=0
r54 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r55 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r56 11 36 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0
r57 11 13 14.575 $w=3.38e-07 $l=4.3e-07 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0.515
r58 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r59 7 9 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.645
r60 2 13 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=2.02
+ $Y=0.37 $X2=2.165 $Y2=0.515
r61 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.37 $X2=0.705 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__O21BAI_1%A_308_74# 1 2 9 11 12 15
r26 13 15 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.64 $Y=0.96
+ $X2=2.64 $Y2=0.515
r27 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.515 $Y=1.045
+ $X2=2.64 $Y2=0.96
r28 11 12 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.515 $Y=1.045
+ $X2=1.815 $Y2=1.045
r29 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.73 $Y=0.96
+ $X2=1.815 $Y2=1.045
r30 7 9 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.73 $Y=0.96 $X2=1.73
+ $Y2=0.515
r31 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.46
+ $Y=0.37 $X2=2.6 $Y2=0.515
r32 1 9 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=1.54 $Y=0.37
+ $X2=1.73 $Y2=0.515
.ends

