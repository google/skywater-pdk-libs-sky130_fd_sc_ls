* NGSPICE file created from sky130_fd_sc_ls__a222o_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a222o_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR X
M1000 X a_32_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=9.082e+11p ps=5.52e+06u
M1001 VGND A2 a_651_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1002 a_27_390# B1 a_337_390# VPB phighvt w=1e+06u l=150000u
+  ad=9.4e+11p pd=7.88e+06u as=7.4e+11p ps=5.48e+06u
M1003 a_337_390# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=8.154e+11p ps=5.8e+06u
M1004 a_651_74# A1 a_32_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=6.848e+11p ps=4.7e+06u
M1005 X a_32_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1006 a_119_74# C1 a_32_74# VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1007 a_386_74# B2 VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1008 a_32_74# B1 a_386_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_32_74# C1 a_27_390# VPB phighvt w=1e+06u l=150000u
+  ad=4.55e+11p pd=2.91e+06u as=0p ps=0u
M1010 VPWR A2 a_337_390# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_390# C2 a_32_74# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_337_390# B2 a_27_390# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND C2 a_119_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

