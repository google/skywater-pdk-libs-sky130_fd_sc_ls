* File: sky130_fd_sc_ls__o311a_1.pex.spice
* Created: Fri Aug 28 13:51:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O311A_1%C1 2 3 5 8 10 17
r30 16 17 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=0.525 $Y=1.305
+ $X2=0.58 $Y2=1.305
r31 13 16 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=0.27 $Y=1.305
+ $X2=0.525 $Y2=1.305
r32 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.305 $X2=0.27 $Y2=1.305
r33 6 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.14
+ $X2=0.58 $Y2=1.305
r34 6 8 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.58 $Y=1.14 $X2=0.58
+ $Y2=0.69
r35 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.525 $Y=1.86
+ $X2=0.525 $Y2=2.435
r36 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.525 $Y=1.77 $X2=0.525
+ $Y2=1.86
r37 1 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.47
+ $X2=0.525 $Y2=1.305
r38 1 2 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=0.525 $Y=1.47 $X2=0.525
+ $Y2=1.77
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_1%B1 3 6 7 9 10 13
r39 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.305
+ $X2=1.06 $Y2=1.47
r40 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.305
+ $X2=1.06 $Y2=1.14
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=1.305 $X2=1.06 $Y2=1.305
r42 10 14 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.2 $Y=1.305
+ $X2=1.06 $Y2=1.305
r43 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.075 $Y=1.86
+ $X2=1.075 $Y2=2.435
r44 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.075 $Y=1.77 $X2=1.075
+ $Y2=1.86
r45 6 16 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=1.075 $Y=1.77 $X2=1.075
+ $Y2=1.47
r46 3 15 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.97 $Y=0.69 $X2=0.97
+ $Y2=1.14
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_1%A2 3 5 7 9 10 11 14 17 20 28
c69 14 0 1.74145e-20 $X=2.68 $Y=1.61
c70 3 0 1.12678e-19 $X=1.51 $Y=0.69
r71 20 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.6 $Y=1.305
+ $X2=1.6 $Y2=1.14
r72 17 28 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.6 $Y=1.305 $X2=1.72
+ $Y2=1.305
r73 17 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.305 $X2=1.6 $Y2=1.305
r74 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.61 $X2=2.68 $Y2=1.61
r75 12 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.68 $Y=2.32 $X2=2.68
+ $Y2=1.61
r76 10 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.515 $Y=2.405
+ $X2=2.68 $Y2=2.32
r77 10 11 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.515 $Y=2.405
+ $X2=1.805 $Y2=2.405
r78 9 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.72 $Y=2.32
+ $X2=1.805 $Y2=2.405
r79 8 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=1.47 $X2=1.72
+ $Y2=1.305
r80 8 9 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.72 $Y=1.47 $X2=1.72
+ $Y2=2.32
r81 5 15 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.605 $Y=1.86
+ $X2=2.68 $Y2=1.61
r82 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.605 $Y=1.86
+ $X2=2.605 $Y2=2.435
r83 3 22 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.51 $Y=0.69 $X2=1.51
+ $Y2=1.14
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_1%A3 1 3 4 5 7 10 11 12 13 18 20
c45 18 0 1.74145e-20 $X=2.14 $Y=1.285
c46 11 0 1.12678e-19 $X=2.16 $Y=1.295
r47 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.285
+ $X2=2.14 $Y2=1.45
r48 18 20 52.3316 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=2.14 $Y=1.285 $X2=2.14
+ $Y2=1.085
r49 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.14 $Y=1.665
+ $X2=2.14 $Y2=2.035
r50 11 12 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.14 $Y=1.285
+ $X2=2.14 $Y2=1.665
r51 11 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.285 $X2=2.14 $Y2=1.285
r52 10 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.23 $Y=0.69
+ $X2=2.23 $Y2=1.085
r53 7 21 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=2.05 $Y=1.71 $X2=2.05
+ $Y2=1.45
r54 4 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.975 $Y=1.785
+ $X2=2.05 $Y2=1.71
r55 4 5 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.975 $Y=1.785
+ $X2=1.6 $Y2=1.785
r56 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.525 $Y=1.86
+ $X2=1.6 $Y2=1.785
r57 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.525 $Y=1.86
+ $X2=1.525 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_1%A1 2 3 5 8 9 12 13 14
c42 14 0 1.54042e-19 $X=3.22 $Y=1.12
c43 12 0 1.3462e-19 $X=3.22 $Y=1.285
r44 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.285
+ $X2=3.22 $Y2=1.45
r45 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.285
+ $X2=3.22 $Y2=1.12
r46 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.22
+ $Y=1.285 $X2=3.22 $Y2=1.285
r47 9 13 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=3.12 $Y=1.285 $X2=3.22
+ $Y2=1.285
r48 8 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.31 $Y=0.69 $X2=3.31
+ $Y2=1.12
r49 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.175 $Y=1.86
+ $X2=3.175 $Y2=2.435
r50 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.175 $Y=1.77 $X2=3.175
+ $Y2=1.86
r51 2 15 124.387 $w=1.8e-07 $l=3.2e-07 $layer=POLY_cond $X=3.175 $Y=1.77
+ $X2=3.175 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_1%A_31_387# 1 2 3 10 12 15 19 25 28 29 30 32
+ 34 35 38 39 40 46 51
c123 51 0 1.25197e-19 $X=3.76 $Y=1.515
r124 51 54 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=3.745 $Y=1.515
+ $X2=3.745 $Y2=1.705
r125 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.76
+ $Y=1.515 $X2=3.76 $Y2=1.515
r126 39 54 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.595 $Y=1.705
+ $X2=3.745 $Y2=1.705
r127 39 40 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.595 $Y=1.705
+ $X2=3.185 $Y2=1.705
r128 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.1 $Y=1.79
+ $X2=3.185 $Y2=1.705
r129 37 38 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=3.1 $Y=1.79
+ $X2=3.1 $Y2=2.785
r130 36 49 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.87
+ $X2=1.3 $Y2=2.87
r131 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.015 $Y=2.87
+ $X2=3.1 $Y2=2.785
r132 35 36 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=3.015 $Y=2.87
+ $X2=1.465 $Y2=2.87
r133 32 49 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=2.785 $X2=1.3
+ $Y2=2.87
r134 32 34 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.3 $Y=2.785
+ $X2=1.3 $Y2=2.08
r135 31 34 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=1.3 $Y=1.81 $X2=1.3
+ $Y2=2.08
r136 30 43 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=1.725
+ $X2=0.665 $Y2=1.725
r137 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.135 $Y=1.725
+ $X2=1.3 $Y2=1.81
r138 29 30 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.135 $Y=1.725
+ $X2=0.75 $Y2=1.725
r139 28 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=1.64
+ $X2=0.665 $Y2=1.725
r140 27 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=0.97
+ $X2=0.665 $Y2=0.885
r141 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.665 $Y=0.97
+ $X2=0.665 $Y2=1.64
r142 23 46 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.365 $Y=0.885
+ $X2=0.665 $Y2=0.885
r143 23 25 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.365 $Y=0.8
+ $X2=0.365 $Y2=0.515
r144 19 21 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.3 $Y=2.08 $X2=0.3
+ $Y2=2.79
r145 17 43 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.3 $Y=1.725
+ $X2=0.665 $Y2=1.725
r146 17 19 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=0.3 $Y=1.81 $X2=0.3
+ $Y2=2.08
r147 13 52 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.82 $Y=1.35
+ $X2=3.76 $Y2=1.515
r148 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.82 $Y=1.35
+ $X2=3.82 $Y2=0.74
r149 10 52 52.2586 $w=2.99e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.795 $Y=1.765
+ $X2=3.76 $Y2=1.515
r150 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.795 $Y=1.765
+ $X2=3.795 $Y2=2.4
r151 3 49 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.15
+ $Y=1.935 $X2=1.3 $Y2=2.79
r152 3 34 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.15
+ $Y=1.935 $X2=1.3 $Y2=2.08
r153 2 21 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.935 $X2=0.3 $Y2=2.79
r154 2 19 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.935 $X2=0.3 $Y2=2.08
r155 1 25 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.22
+ $Y=0.37 $X2=0.365 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_1%VPWR 1 2 9 15 19 21 26 36 37 40 43
r41 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r42 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 37 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r44 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r45 34 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=3.52 $Y2=3.33
r46 34 36 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=4.08 $Y2=3.33
r47 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r48 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 30 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 29 32 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 27 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=0.8 $Y2=3.33
r53 27 29 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 26 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.52 $Y2=3.33
r55 26 32 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 24 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 21 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.8 $Y2=3.33
r59 21 23 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 19 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 19 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r62 15 18 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.52 $Y=2.125
+ $X2=3.52 $Y2=2.815
r63 13 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.52 $Y=3.245
+ $X2=3.52 $Y2=3.33
r64 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.52 $Y=3.245
+ $X2=3.52 $Y2=2.815
r65 9 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.8 $Y=2.11 $X2=0.8
+ $Y2=2.79
r66 7 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=3.245 $X2=0.8
+ $Y2=3.33
r67 7 12 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.8 $Y=3.245 $X2=0.8
+ $Y2=2.79
r68 2 18 400 $w=1.7e-07 $l=1.00598e-06 $layer=licon1_PDIFF $count=1 $X=3.25
+ $Y=1.935 $X2=3.52 $Y2=2.815
r69 2 15 400 $w=1.7e-07 $l=3.5242e-07 $layer=licon1_PDIFF $count=1 $X=3.25
+ $Y=1.935 $X2=3.52 $Y2=2.125
r70 1 12 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.935 $X2=0.8 $Y2=2.79
r71 1 9 400 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.935 $X2=0.8 $Y2=2.11
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_1%X 1 2 9 14 15 16 17 28
c24 17 0 9.42383e-21 $X=3.995 $Y=0.84
c25 16 0 1.54042e-19 $X=4.08 $Y=0.555
r26 21 28 0.726197 $w=3.63e-07 $l=2.3e-08 $layer=LI1_cond $X=4.052 $Y=0.948
+ $X2=4.052 $Y2=0.925
r27 17 30 8.08227 $w=3.63e-07 $l=1.51e-07 $layer=LI1_cond $X=4.052 $Y=0.979
+ $X2=4.052 $Y2=1.13
r28 17 21 0.978787 $w=3.63e-07 $l=3.1e-08 $layer=LI1_cond $X=4.052 $Y=0.979
+ $X2=4.052 $Y2=0.948
r29 17 28 0.978787 $w=3.63e-07 $l=3.1e-08 $layer=LI1_cond $X=4.052 $Y=0.894
+ $X2=4.052 $Y2=0.925
r30 16 17 11.9665 $w=3.63e-07 $l=3.79e-07 $layer=LI1_cond $X=4.052 $Y=0.515
+ $X2=4.052 $Y2=0.894
r31 15 30 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.15 $Y=1.96
+ $X2=4.15 $Y2=1.13
r32 14 15 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=4.045 $Y=2.125
+ $X2=4.045 $Y2=1.96
r33 7 14 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=4.045 $Y=2.15
+ $X2=4.045 $Y2=2.125
r34 7 9 20.1678 $w=3.78e-07 $l=6.65e-07 $layer=LI1_cond $X=4.045 $Y=2.15
+ $X2=4.045 $Y2=2.815
r35 2 14 400 $w=1.7e-07 $l=3.52101e-07 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=1.84 $X2=4.02 $Y2=2.125
r36 2 9 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=1.84 $X2=4.02 $Y2=2.815
r37 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.895
+ $Y=0.37 $X2=4.035 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_1%A_209_74# 1 2 7 9 13
r19 11 16 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=0.445
+ $X2=1.225 $Y2=0.445
r20 11 13 56.7491 $w=3.28e-07 $l=1.625e-06 $layer=LI1_cond $X=1.39 $Y=0.445
+ $X2=3.015 $Y2=0.445
r21 7 16 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=0.61
+ $X2=1.225 $Y2=0.445
r22 7 9 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.225 $Y=0.61
+ $X2=1.225 $Y2=0.855
r23 2 13 91 $w=1.7e-07 $l=7.83677e-07 $layer=licon1_NDIFF $count=2 $X=2.305
+ $Y=0.37 $X2=3.015 $Y2=0.525
r24 1 16 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=0.37 $X2=1.225 $Y2=0.515
r25 1 9 182 $w=1.7e-07 $l=5.67913e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=0.37 $X2=1.225 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LS__O311A_1%VGND 1 2 7 14 15 17 27 28 31
r47 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r48 28 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r49 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r50 25 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.69 $Y=0 $X2=3.525
+ $Y2=0
r51 25 27 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.69 $Y=0 $X2=4.08
+ $Y2=0
r52 24 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r53 23 24 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r54 19 23 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.12
+ $Y2=0
r55 19 20 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r56 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.36 $Y=0 $X2=3.525
+ $Y2=0
r57 17 23 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.36 $Y=0 $X2=3.12
+ $Y2=0
r58 15 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r59 15 20 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=0.24
+ $Y2=0
r60 12 14 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.525 $Y=0.78
+ $X2=3.525 $Y2=0.515
r61 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=0.085
+ $X2=3.525 $Y2=0
r62 11 14 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.525 $Y=0.085
+ $X2=3.525 $Y2=0.515
r63 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.36 $Y=0.865
+ $X2=3.525 $Y2=0.78
r64 7 9 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=3.36 $Y=0.865
+ $X2=1.87 $Y2=0.865
r65 2 14 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.385
+ $Y=0.37 $X2=3.525 $Y2=0.515
r66 1 9 182 $w=1.7e-07 $l=6.21369e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.37 $X2=1.87 $Y2=0.865
.ends

