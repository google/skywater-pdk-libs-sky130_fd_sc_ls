* File: sky130_fd_sc_ls__inv_4.spice
* Created: Fri Aug 28 13:28:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__inv_4.pex.spice"
.subckt sky130_fd_sc_ls__inv_4  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.74 AD=0.2331
+ AS=0.1184 PD=2.11 PS=1.06 NRD=4.86 NRS=6.48 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.74 AD=0.1221
+ AS=0.1184 PD=1.07 PS=1.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7 SB=75001.1
+ A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1003_d N_A_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.74 AD=0.1221
+ AS=0.1036 PD=1.07 PS=1.02 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75001.2 SB=75000.6
+ A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.74 AD=0.2109
+ AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75001.6 A=0.168 P=2.54 MULT=1
MM1002 N_Y_M1000_d N_A_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.7
+ SB=75001.1 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.1
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1006_d N_A_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.12 AD=0.168
+ AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.6
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_ls__inv_4.pxi.spice"
*
.ends
*
*
