* File: sky130_fd_sc_ls__o221ai_4.pxi.spice
* Created: Fri Aug 28 13:48:16 2020
* 
x_PM_SKY130_FD_SC_LS__O221AI_4%C1 N_C1_M1000_g N_C1_c_148_n N_C1_M1002_g
+ N_C1_M1021_g N_C1_c_149_n N_C1_M1023_g N_C1_M1038_g N_C1_c_150_n N_C1_M1024_g
+ N_C1_M1039_g N_C1_c_151_n N_C1_M1032_g C1 C1 C1 N_C1_c_146_n N_C1_c_147_n
+ PM_SKY130_FD_SC_LS__O221AI_4%C1
x_PM_SKY130_FD_SC_LS__O221AI_4%B1 N_B1_c_231_n N_B1_M1001_g N_B1_M1008_g
+ N_B1_c_232_n N_B1_M1012_g N_B1_c_224_n N_B1_M1009_g N_B1_c_233_n N_B1_M1014_g
+ N_B1_c_225_n N_B1_M1030_g N_B1_M1035_g N_B1_c_227_n N_B1_M1016_g N_B1_c_235_n
+ N_B1_c_236_n N_B1_c_228_n B1 N_B1_c_229_n N_B1_c_230_n
+ PM_SKY130_FD_SC_LS__O221AI_4%B1
x_PM_SKY130_FD_SC_LS__O221AI_4%B2 N_B2_c_351_n N_B2_M1006_g N_B2_c_345_n
+ N_B2_M1003_g N_B2_c_352_n N_B2_M1010_g N_B2_c_346_n N_B2_M1015_g N_B2_c_353_n
+ N_B2_M1026_g N_B2_c_347_n N_B2_M1017_g N_B2_c_354_n N_B2_M1036_g N_B2_c_348_n
+ N_B2_M1028_g B2 B2 N_B2_c_350_n PM_SKY130_FD_SC_LS__O221AI_4%B2
x_PM_SKY130_FD_SC_LS__O221AI_4%A1 N_A1_M1005_g N_A1_c_429_n N_A1_M1019_g
+ N_A1_M1029_g N_A1_c_439_n N_A1_M1020_g N_A1_c_440_n N_A1_M1025_g N_A1_M1031_g
+ N_A1_c_441_n N_A1_M1033_g N_A1_M1034_g N_A1_c_433_n A1 A1 A1 A1 N_A1_c_435_n
+ N_A1_c_436_n A1 N_A1_c_437_n PM_SKY130_FD_SC_LS__O221AI_4%A1
x_PM_SKY130_FD_SC_LS__O221AI_4%A2 N_A2_M1004_g N_A2_c_549_n N_A2_M1007_g
+ N_A2_M1011_g N_A2_c_550_n N_A2_M1013_g N_A2_c_551_n N_A2_M1027_g N_A2_M1018_g
+ N_A2_M1022_g N_A2_c_552_n N_A2_M1037_g A2 A2 A2 N_A2_c_548_n
+ PM_SKY130_FD_SC_LS__O221AI_4%A2
x_PM_SKY130_FD_SC_LS__O221AI_4%VPWR N_VPWR_M1002_s N_VPWR_M1023_s N_VPWR_M1032_s
+ N_VPWR_M1012_s N_VPWR_M1016_s N_VPWR_M1020_s N_VPWR_M1033_s N_VPWR_c_631_n
+ N_VPWR_c_632_n N_VPWR_c_633_n N_VPWR_c_634_n N_VPWR_c_635_n N_VPWR_c_636_n
+ N_VPWR_c_637_n N_VPWR_c_638_n N_VPWR_c_639_n VPWR N_VPWR_c_640_n
+ N_VPWR_c_641_n N_VPWR_c_642_n N_VPWR_c_643_n N_VPWR_c_644_n N_VPWR_c_645_n
+ N_VPWR_c_646_n N_VPWR_c_647_n N_VPWR_c_648_n N_VPWR_c_649_n N_VPWR_c_650_n
+ N_VPWR_c_630_n PM_SKY130_FD_SC_LS__O221AI_4%VPWR
x_PM_SKY130_FD_SC_LS__O221AI_4%Y N_Y_M1000_d N_Y_M1038_d N_Y_M1002_d N_Y_M1024_d
+ N_Y_M1006_d N_Y_M1026_d N_Y_M1007_d N_Y_M1027_d N_Y_c_769_n N_Y_c_772_n
+ N_Y_c_765_n N_Y_c_761_n N_Y_c_762_n N_Y_c_787_n N_Y_c_791_n N_Y_c_766_n
+ N_Y_c_795_n N_Y_c_824_n N_Y_c_815_n N_Y_c_816_n N_Y_c_817_n N_Y_c_836_n
+ N_Y_c_763_n N_Y_c_767_n N_Y_c_764_n N_Y_c_821_n N_Y_c_822_n N_Y_c_840_n Y
+ PM_SKY130_FD_SC_LS__O221AI_4%Y
x_PM_SKY130_FD_SC_LS__O221AI_4%A_508_368# N_A_508_368#_M1001_d
+ N_A_508_368#_M1014_d N_A_508_368#_M1010_s N_A_508_368#_M1036_s
+ N_A_508_368#_c_914_n N_A_508_368#_c_916_n N_A_508_368#_c_917_n
+ N_A_508_368#_c_905_n N_A_508_368#_c_906_n N_A_508_368#_c_931_n
+ N_A_508_368#_c_907_n N_A_508_368#_c_921_n N_A_508_368#_c_908_n
+ N_A_508_368#_c_909_n PM_SKY130_FD_SC_LS__O221AI_4%A_508_368#
x_PM_SKY130_FD_SC_LS__O221AI_4%A_1288_368# N_A_1288_368#_M1019_d
+ N_A_1288_368#_M1013_s N_A_1288_368#_M1037_s N_A_1288_368#_M1025_d
+ N_A_1288_368#_c_972_n N_A_1288_368#_c_1018_n N_A_1288_368#_c_973_n
+ N_A_1288_368#_c_978_n N_A_1288_368#_c_1001_n N_A_1288_368#_c_979_n
+ N_A_1288_368#_c_983_n N_A_1288_368#_c_974_n N_A_1288_368#_c_975_n
+ N_A_1288_368#_c_976_n PM_SKY130_FD_SC_LS__O221AI_4%A_1288_368#
x_PM_SKY130_FD_SC_LS__O221AI_4%A_27_84# N_A_27_84#_M1000_s N_A_27_84#_M1021_s
+ N_A_27_84#_M1039_s N_A_27_84#_M1008_d N_A_27_84#_M1030_d N_A_27_84#_M1015_s
+ N_A_27_84#_M1028_s N_A_27_84#_c_1027_n N_A_27_84#_c_1028_n N_A_27_84#_c_1029_n
+ N_A_27_84#_c_1078_n N_A_27_84#_c_1030_n N_A_27_84#_c_1031_n
+ N_A_27_84#_c_1032_n N_A_27_84#_c_1033_n N_A_27_84#_c_1034_n
+ N_A_27_84#_c_1035_n N_A_27_84#_c_1036_n N_A_27_84#_c_1037_n
+ N_A_27_84#_c_1061_n N_A_27_84#_c_1067_n PM_SKY130_FD_SC_LS__O221AI_4%A_27_84#
x_PM_SKY130_FD_SC_LS__O221AI_4%A_483_74# N_A_483_74#_M1008_s N_A_483_74#_M1009_s
+ N_A_483_74#_M1003_d N_A_483_74#_M1017_d N_A_483_74#_M1035_s
+ N_A_483_74#_M1004_s N_A_483_74#_M1018_s N_A_483_74#_M1029_d
+ N_A_483_74#_M1034_d N_A_483_74#_c_1107_n N_A_483_74#_c_1108_n
+ N_A_483_74#_c_1129_n N_A_483_74#_c_1109_n N_A_483_74#_c_1134_n
+ N_A_483_74#_c_1110_n N_A_483_74#_c_1135_n N_A_483_74#_c_1111_n
+ N_A_483_74#_c_1112_n N_A_483_74#_c_1113_n N_A_483_74#_c_1114_n
+ N_A_483_74#_c_1147_n N_A_483_74#_c_1148_n N_A_483_74#_c_1149_n
+ PM_SKY130_FD_SC_LS__O221AI_4%A_483_74#
x_PM_SKY130_FD_SC_LS__O221AI_4%VGND N_VGND_M1005_s N_VGND_M1011_d N_VGND_M1022_d
+ N_VGND_M1031_s N_VGND_c_1217_n N_VGND_c_1218_n N_VGND_c_1219_n N_VGND_c_1220_n
+ VGND N_VGND_c_1221_n N_VGND_c_1222_n N_VGND_c_1223_n N_VGND_c_1224_n
+ N_VGND_c_1225_n N_VGND_c_1226_n N_VGND_c_1227_n N_VGND_c_1228_n
+ N_VGND_c_1229_n N_VGND_c_1230_n PM_SKY130_FD_SC_LS__O221AI_4%VGND
cc_1 VNB N_C1_M1000_g 0.0263359f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.79
cc_2 VNB N_C1_M1021_g 0.0191476f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.79
cc_3 VNB N_C1_M1038_g 0.0191247f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.79
cc_4 VNB N_C1_M1039_g 0.0256157f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.79
cc_5 VNB N_C1_c_146_n 0.0167416f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=1.515
cc_6 VNB N_C1_c_147_n 0.0831605f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.557
cc_7 VNB N_B1_M1008_g 0.0308588f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_8 VNB N_B1_c_224_n 0.0146162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_c_225_n 0.0147307f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.79
cc_10 VNB N_B1_M1035_g 0.0257119f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.35
cc_11 VNB N_B1_c_227_n 0.0250039f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.79
cc_12 VNB N_B1_c_228_n 0.0037594f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.557
cc_13 VNB N_B1_c_229_n 0.0859413f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=1.557
cc_14 VNB N_B1_c_230_n 0.00725477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B2_c_345_n 0.0169363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B2_c_346_n 0.0166753f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.79
cc_17 VNB N_B2_c_347_n 0.0166979f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.79
cc_18 VNB N_B2_c_348_n 0.017373f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.35
cc_19 VNB B2 0.00745009f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=1.765
cc_20 VNB N_B2_c_350_n 0.106656f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.557
cc_21 VNB N_A1_M1005_g 0.021903f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.79
cc_22 VNB N_A1_c_429_n 0.0327799f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_23 VNB N_A1_M1029_g 0.0196218f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.79
cc_24 VNB N_A1_M1031_g 0.0192941f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.4
cc_25 VNB N_A1_M1034_g 0.0262473f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=2.4
cc_26 VNB N_A1_c_433_n 0.0104553f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_27 VNB A1 0.0222352f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.515
cc_28 VNB N_A1_c_435_n 0.0841437f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_29 VNB N_A1_c_436_n 0.0147594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A1_c_437_n 0.0016599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A2_M1004_g 0.0238876f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.79
cc_32 VNB N_A2_M1011_g 0.0227944f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.79
cc_33 VNB N_A2_M1018_g 0.0233499f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.4
cc_34 VNB N_A2_M1022_g 0.0216231f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.79
cc_35 VNB N_A2_c_548_n 0.0691851f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.557
cc_36 VNB N_VPWR_c_630_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_761_n 0.00225436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_762_n 0.00229834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_763_n 0.00421298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_764_n 0.00159633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_84#_c_1027_n 0.0307564f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.79
cc_42 VNB N_A_27_84#_c_1028_n 0.00475623f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=1.765
cc_43 VNB N_A_27_84#_c_1029_n 0.00958293f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=2.4
cc_44 VNB N_A_27_84#_c_1030_n 0.00952739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_27_84#_c_1031_n 0.00400018f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.557
cc_46 VNB N_A_27_84#_c_1032_n 0.0199341f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.515
cc_47 VNB N_A_27_84#_c_1033_n 0.00690962f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.515
cc_48 VNB N_A_27_84#_c_1034_n 0.00225825f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.557
cc_49 VNB N_A_27_84#_c_1035_n 0.00136506f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=1.557
cc_50 VNB N_A_27_84#_c_1036_n 0.00138842f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_51 VNB N_A_27_84#_c_1037_n 0.00348266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_483_74#_c_1107_n 0.00940936f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=2.4
cc_53 VNB N_A_483_74#_c_1108_n 0.0127258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_483_74#_c_1109_n 0.00206045f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=1.557
cc_55 VNB N_A_483_74#_c_1110_n 0.00206045f $X=-0.19 $Y=-0.245 $X2=1.965
+ $Y2=1.557
cc_56 VNB N_A_483_74#_c_1111_n 0.00252795f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.565
cc_57 VNB N_A_483_74#_c_1112_n 0.0075506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_483_74#_c_1113_n 0.0233055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_483_74#_c_1114_n 0.0026414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1217_n 0.00886652f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.35
cc_61 VNB N_VGND_c_1218_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=1.765
cc_62 VNB N_VGND_c_1219_n 0.00269659f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.79
cc_63 VNB N_VGND_c_1220_n 0.00333063f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=2.4
cc_64 VNB N_VGND_c_1221_n 0.156139f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_65 VNB N_VGND_c_1222_n 0.0156795f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.557
cc_66 VNB N_VGND_c_1223_n 0.0156795f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.557
cc_67 VNB N_VGND_c_1224_n 0.0161665f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=1.557
cc_68 VNB N_VGND_c_1225_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1226_n 0.523727f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.565
cc_70 VNB N_VGND_c_1227_n 0.00632082f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=1.565
cc_71 VNB N_VGND_c_1228_n 0.00613127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1229_n 0.00619876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1230_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VPB N_C1_c_148_n 0.0179801f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_75 VPB N_C1_c_149_n 0.0161326f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_76 VPB N_C1_c_150_n 0.0164961f $X=-0.19 $Y=1.66 $X2=1.49 $Y2=1.765
cc_77 VPB N_C1_c_151_n 0.015772f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=1.765
cc_78 VPB N_C1_c_146_n 0.016388f $X=-0.19 $Y=1.66 $X2=1.24 $Y2=1.515
cc_79 VPB N_C1_c_147_n 0.0525347f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.557
cc_80 VPB N_B1_c_231_n 0.0162628f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_81 VPB N_B1_c_232_n 0.0156617f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.35
cc_82 VPB N_B1_c_233_n 0.0152989f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_83 VPB N_B1_c_227_n 0.0265995f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=0.79
cc_84 VPB N_B1_c_235_n 7.91081e-19 $X=-0.19 $Y=1.66 $X2=1.965 $Y2=2.4
cc_85 VPB N_B1_c_236_n 0.0089811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_B1_c_228_n 6.14949e-19 $X=-0.19 $Y=1.66 $X2=0.9 $Y2=1.557
cc_87 VPB N_B1_c_229_n 0.0367217f $X=-0.19 $Y=1.66 $X2=1.49 $Y2=1.557
cc_88 VPB N_B1_c_230_n 0.00273218f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_B2_c_351_n 0.014134f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_90 VPB N_B2_c_352_n 0.0141056f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_91 VPB N_B2_c_353_n 0.0144819f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_92 VPB N_B2_c_354_n 0.0148849f $X=-0.19 $Y=1.66 $X2=1.49 $Y2=1.765
cc_93 VPB N_B2_c_350_n 0.0321965f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.557
cc_94 VPB N_A1_c_429_n 0.0240392f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_95 VPB N_A1_c_439_n 0.015274f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_96 VPB N_A1_c_440_n 0.0155127f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.35
cc_97 VPB N_A1_c_441_n 0.0179811f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.35
cc_98 VPB A1 0.0171479f $X=-0.19 $Y=1.66 $X2=0.9 $Y2=1.515
cc_99 VPB N_A1_c_435_n 0.0183525f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_100 VPB N_A1_c_437_n 0.00354333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A2_c_549_n 0.0152692f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_102 VPB N_A2_c_550_n 0.014664f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_103 VPB N_A2_c_551_n 0.014664f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.35
cc_104 VPB N_A2_c_552_n 0.0148403f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=1.765
cc_105 VPB A2 0.00800933f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_106 VPB N_A2_c_548_n 0.0466434f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.557
cc_107 VPB N_VPWR_c_631_n 0.0106521f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.35
cc_108 VPB N_VPWR_c_632_n 0.0498694f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=0.79
cc_109 VPB N_VPWR_c_633_n 0.00898683f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_110 VPB N_VPWR_c_634_n 0.00522246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_635_n 0.00858913f $X=-0.19 $Y=1.66 $X2=0.9 $Y2=1.515
cc_112 VPB N_VPWR_c_636_n 0.00886214f $X=-0.19 $Y=1.66 $X2=1.24 $Y2=1.557
cc_113 VPB N_VPWR_c_637_n 0.00571271f $X=-0.19 $Y=1.66 $X2=1.49 $Y2=1.557
cc_114 VPB N_VPWR_c_638_n 0.0107598f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=1.557
cc_115 VPB N_VPWR_c_639_n 0.0495498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_640_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_641_n 0.0178889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_642_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_643_n 0.0599386f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_644_n 0.0580909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_645_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_646_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_647_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_648_n 0.00631813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_649_n 0.00631418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_650_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_630_n 0.0973853f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_Y_c_765_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_129 VPB N_Y_c_766_n 0.00254397f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.557
cc_130 VPB N_Y_c_767_n 0.0012522f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_Y_c_764_n 0.00174733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_508_368#_c_905_n 0.00213603f $X=-0.19 $Y=1.66 $X2=1.49 $Y2=1.765
cc_133 VPB N_A_508_368#_c_906_n 0.00218418f $X=-0.19 $Y=1.66 $X2=1.49 $Y2=2.4
cc_134 VPB N_A_508_368#_c_907_n 0.00502022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_508_368#_c_908_n 0.00256678f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_508_368#_c_909_n 0.00218418f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_137 VPB N_A_1288_368#_c_972_n 0.0028338f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_138 VPB N_A_1288_368#_c_973_n 0.00523584f $X=-0.19 $Y=1.66 $X2=1.49 $Y2=1.765
cc_139 VPB N_A_1288_368#_c_974_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_140 VPB N_A_1288_368#_c_975_n 0.00230866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_1288_368#_c_976_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 N_C1_c_151_n N_B1_c_231_n 0.0306963f $X=1.965 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_143 N_C1_c_147_n N_B1_c_235_n 0.00207454f $X=1.785 $Y=1.557 $X2=0 $Y2=0
cc_144 N_C1_c_147_n N_B1_c_229_n 0.0146531f $X=1.785 $Y=1.557 $X2=0 $Y2=0
cc_145 N_C1_c_148_n N_VPWR_c_632_n 0.00831454f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_146 N_C1_c_146_n N_VPWR_c_632_n 0.0211447f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_147 N_C1_c_149_n N_VPWR_c_633_n 0.0072254f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_148 N_C1_c_150_n N_VPWR_c_633_n 0.00198511f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_149 N_C1_c_150_n N_VPWR_c_634_n 5.03202e-19 $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_150 N_C1_c_151_n N_VPWR_c_634_n 0.01009f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_151 N_C1_c_148_n N_VPWR_c_640_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_152 N_C1_c_149_n N_VPWR_c_640_n 0.00445602f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_153 N_C1_c_150_n N_VPWR_c_641_n 0.00461464f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_154 N_C1_c_151_n N_VPWR_c_641_n 0.00413917f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_155 N_C1_c_148_n N_VPWR_c_630_n 0.00861084f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_156 N_C1_c_149_n N_VPWR_c_630_n 0.00857676f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_157 N_C1_c_150_n N_VPWR_c_630_n 0.00908937f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_158 N_C1_c_151_n N_VPWR_c_630_n 0.00817962f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_159 N_C1_M1000_g N_Y_c_769_n 0.00473639f $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_160 N_C1_M1021_g N_Y_c_769_n 0.00575058f $X=0.925 $Y=0.79 $X2=0 $Y2=0
cc_161 N_C1_M1038_g N_Y_c_769_n 5.36571e-19 $X=1.355 $Y=0.79 $X2=0 $Y2=0
cc_162 N_C1_c_148_n N_Y_c_772_n 0.00203651f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_163 N_C1_c_149_n N_Y_c_772_n 4.27055e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_164 N_C1_c_146_n N_Y_c_772_n 0.0237598f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_165 N_C1_c_147_n N_Y_c_772_n 0.00144162f $X=1.785 $Y=1.557 $X2=0 $Y2=0
cc_166 N_C1_c_148_n N_Y_c_765_n 0.00960826f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_167 N_C1_c_149_n N_Y_c_765_n 0.0102182f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_168 N_C1_c_150_n N_Y_c_765_n 8.49006e-19 $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_169 N_C1_M1021_g N_Y_c_761_n 0.00900535f $X=0.925 $Y=0.79 $X2=0 $Y2=0
cc_170 N_C1_M1038_g N_Y_c_761_n 0.00900535f $X=1.355 $Y=0.79 $X2=0 $Y2=0
cc_171 N_C1_c_146_n N_Y_c_761_n 0.039654f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_172 N_C1_c_147_n N_Y_c_761_n 0.00224206f $X=1.785 $Y=1.557 $X2=0 $Y2=0
cc_173 N_C1_M1000_g N_Y_c_762_n 0.0023927f $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_174 N_C1_M1021_g N_Y_c_762_n 9.58661e-19 $X=0.925 $Y=0.79 $X2=0 $Y2=0
cc_175 N_C1_c_146_n N_Y_c_762_n 0.0277843f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_176 N_C1_c_147_n N_Y_c_762_n 0.00231547f $X=1.785 $Y=1.557 $X2=0 $Y2=0
cc_177 N_C1_c_149_n N_Y_c_787_n 0.0123851f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_178 N_C1_c_150_n N_Y_c_787_n 0.0180303f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_179 N_C1_c_146_n N_Y_c_787_n 0.0359083f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_180 N_C1_c_147_n N_Y_c_787_n 0.0017661f $X=1.785 $Y=1.557 $X2=0 $Y2=0
cc_181 N_C1_M1021_g N_Y_c_791_n 5.3642e-19 $X=0.925 $Y=0.79 $X2=0 $Y2=0
cc_182 N_C1_M1038_g N_Y_c_791_n 0.00575058f $X=1.355 $Y=0.79 $X2=0 $Y2=0
cc_183 N_C1_M1039_g N_Y_c_791_n 0.0051579f $X=1.785 $Y=0.79 $X2=0 $Y2=0
cc_184 N_C1_c_150_n N_Y_c_766_n 4.35278e-19 $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_185 N_C1_c_151_n N_Y_c_795_n 0.017258f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_186 N_C1_c_147_n N_Y_c_795_n 0.00100117f $X=1.785 $Y=1.557 $X2=0 $Y2=0
cc_187 N_C1_M1038_g N_Y_c_763_n 0.00181594f $X=1.355 $Y=0.79 $X2=0 $Y2=0
cc_188 N_C1_M1039_g N_Y_c_763_n 0.0021587f $X=1.785 $Y=0.79 $X2=0 $Y2=0
cc_189 N_C1_c_147_n N_Y_c_763_n 0.00257107f $X=1.785 $Y=1.557 $X2=0 $Y2=0
cc_190 N_C1_c_151_n N_Y_c_767_n 0.0109139f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_191 N_C1_c_147_n N_Y_c_767_n 0.00394873f $X=1.785 $Y=1.557 $X2=0 $Y2=0
cc_192 N_C1_M1038_g N_Y_c_764_n 0.00360365f $X=1.355 $Y=0.79 $X2=0 $Y2=0
cc_193 N_C1_c_150_n N_Y_c_764_n 0.0016873f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_194 N_C1_M1039_g N_Y_c_764_n 0.00809756f $X=1.785 $Y=0.79 $X2=0 $Y2=0
cc_195 N_C1_c_151_n N_Y_c_764_n 0.00117811f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_196 N_C1_c_146_n N_Y_c_764_n 0.0327181f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_197 N_C1_c_147_n N_Y_c_764_n 0.0246374f $X=1.785 $Y=1.557 $X2=0 $Y2=0
cc_198 N_C1_M1000_g N_A_27_84#_c_1027_n 0.00160853f $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_199 N_C1_c_146_n N_A_27_84#_c_1027_n 0.0224519f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_200 N_C1_M1000_g N_A_27_84#_c_1028_n 0.0141481f $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_201 N_C1_M1021_g N_A_27_84#_c_1028_n 0.0109808f $X=0.925 $Y=0.79 $X2=0 $Y2=0
cc_202 N_C1_M1038_g N_A_27_84#_c_1030_n 0.0109808f $X=1.355 $Y=0.79 $X2=0 $Y2=0
cc_203 N_C1_M1039_g N_A_27_84#_c_1030_n 0.0138423f $X=1.785 $Y=0.79 $X2=0 $Y2=0
cc_204 N_C1_M1039_g N_A_27_84#_c_1033_n 0.00141527f $X=1.785 $Y=0.79 $X2=0 $Y2=0
cc_205 N_C1_c_147_n N_A_27_84#_c_1033_n 0.00552595f $X=1.785 $Y=1.557 $X2=0
+ $Y2=0
cc_206 N_C1_M1039_g N_A_483_74#_c_1107_n 3.01901e-19 $X=1.785 $Y=0.79 $X2=0
+ $Y2=0
cc_207 N_C1_M1000_g N_VGND_c_1221_n 8.76084e-19 $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_208 N_C1_M1021_g N_VGND_c_1221_n 8.76084e-19 $X=0.925 $Y=0.79 $X2=0 $Y2=0
cc_209 N_C1_M1038_g N_VGND_c_1221_n 8.76084e-19 $X=1.355 $Y=0.79 $X2=0 $Y2=0
cc_210 N_C1_M1039_g N_VGND_c_1221_n 8.76084e-19 $X=1.785 $Y=0.79 $X2=0 $Y2=0
cc_211 N_B1_c_233_n N_B2_c_351_n 0.0278406f $X=3.465 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_212 N_B1_c_236_n N_B2_c_351_n 0.00647572f $X=5.405 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_213 N_B1_c_225_n N_B2_c_345_n 0.0179023f $X=3.635 $Y=1.185 $X2=0 $Y2=0
cc_214 N_B1_c_236_n N_B2_c_352_n 0.00651007f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_215 N_B1_c_236_n N_B2_c_353_n 0.00665306f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_216 N_B1_c_227_n N_B2_c_354_n 0.0328731f $X=5.815 $Y=1.765 $X2=0 $Y2=0
cc_217 N_B1_c_236_n N_B2_c_354_n 0.00581493f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_218 N_B1_c_230_n N_B2_c_354_n 5.02425e-19 $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_219 N_B1_M1035_g N_B2_c_348_n 0.0347442f $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_220 N_B1_M1035_g B2 5.14568e-19 $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_221 N_B1_c_236_n B2 0.0747366f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_222 N_B1_c_228_n B2 0.00532239f $X=3.555 $Y=1.615 $X2=0 $Y2=0
cc_223 N_B1_c_229_n B2 8.13044e-19 $X=3.465 $Y=1.475 $X2=0 $Y2=0
cc_224 N_B1_c_230_n B2 0.0132957f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_225 N_B1_c_227_n N_B2_c_350_n 0.0198148f $X=5.815 $Y=1.765 $X2=0 $Y2=0
cc_226 N_B1_c_236_n N_B2_c_350_n 0.0460917f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_227 N_B1_c_228_n N_B2_c_350_n 0.00219506f $X=3.555 $Y=1.615 $X2=0 $Y2=0
cc_228 N_B1_c_229_n N_B2_c_350_n 0.0335472f $X=3.465 $Y=1.475 $X2=0 $Y2=0
cc_229 N_B1_c_230_n N_B2_c_350_n 0.0131362f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_230 N_B1_M1035_g N_A1_M1005_g 0.0237178f $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_231 N_B1_c_227_n N_A1_c_429_n 0.0564297f $X=5.815 $Y=1.765 $X2=0 $Y2=0
cc_232 N_B1_c_230_n N_A1_c_429_n 0.00569369f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_233 N_B1_M1035_g N_A1_c_433_n 5.32822e-19 $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_234 N_B1_c_227_n N_A1_c_433_n 8.36735e-19 $X=5.815 $Y=1.765 $X2=0 $Y2=0
cc_235 N_B1_c_230_n N_A1_c_433_n 0.0161127f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_236 N_B1_c_235_n N_VPWR_M1012_s 0.0026705f $X=3.29 $Y=1.615 $X2=0 $Y2=0
cc_237 N_B1_c_228_n N_VPWR_M1012_s 4.74511e-19 $X=3.555 $Y=1.615 $X2=0 $Y2=0
cc_238 N_B1_c_230_n N_VPWR_M1016_s 0.00116552f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_239 N_B1_c_231_n N_VPWR_c_634_n 0.00494932f $X=2.465 $Y=1.765 $X2=0 $Y2=0
cc_240 N_B1_c_232_n N_VPWR_c_635_n 0.00336706f $X=2.915 $Y=1.765 $X2=0 $Y2=0
cc_241 N_B1_c_233_n N_VPWR_c_635_n 0.00285025f $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_242 N_B1_c_227_n N_VPWR_c_636_n 0.00487422f $X=5.815 $Y=1.765 $X2=0 $Y2=0
cc_243 N_B1_c_231_n N_VPWR_c_642_n 0.00445602f $X=2.465 $Y=1.765 $X2=0 $Y2=0
cc_244 N_B1_c_232_n N_VPWR_c_642_n 0.00445602f $X=2.915 $Y=1.765 $X2=0 $Y2=0
cc_245 N_B1_c_233_n N_VPWR_c_643_n 0.0044313f $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_246 N_B1_c_227_n N_VPWR_c_643_n 0.0044313f $X=5.815 $Y=1.765 $X2=0 $Y2=0
cc_247 N_B1_c_231_n N_VPWR_c_630_n 0.00857432f $X=2.465 $Y=1.765 $X2=0 $Y2=0
cc_248 N_B1_c_232_n N_VPWR_c_630_n 0.00437179f $X=2.915 $Y=1.765 $X2=0 $Y2=0
cc_249 N_B1_c_233_n N_VPWR_c_630_n 0.00437649f $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_250 N_B1_c_227_n N_VPWR_c_630_n 0.00854111f $X=5.815 $Y=1.765 $X2=0 $Y2=0
cc_251 N_B1_c_236_n N_Y_M1006_d 0.00197763f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_252 N_B1_c_236_n N_Y_M1026_d 0.00250873f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_253 N_B1_c_231_n N_Y_c_795_n 0.0196488f $X=2.465 $Y=1.765 $X2=0 $Y2=0
cc_254 N_B1_c_232_n N_Y_c_795_n 0.0112441f $X=2.915 $Y=1.765 $X2=0 $Y2=0
cc_255 N_B1_c_233_n N_Y_c_795_n 0.011193f $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_256 N_B1_c_235_n N_Y_c_795_n 0.0838702f $X=3.29 $Y=1.615 $X2=0 $Y2=0
cc_257 N_B1_c_229_n N_Y_c_795_n 0.00256297f $X=3.465 $Y=1.475 $X2=0 $Y2=0
cc_258 N_B1_c_236_n N_Y_c_815_n 0.0343548f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_259 N_B1_c_227_n N_Y_c_816_n 5.33746e-19 $X=5.815 $Y=1.765 $X2=0 $Y2=0
cc_260 N_B1_c_227_n N_Y_c_817_n 0.016066f $X=5.815 $Y=1.765 $X2=0 $Y2=0
cc_261 N_B1_c_236_n N_Y_c_817_n 0.00911646f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_262 N_B1_c_230_n N_Y_c_817_n 0.0341533f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_263 N_B1_c_229_n N_Y_c_764_n 0.00163472f $X=3.465 $Y=1.475 $X2=0 $Y2=0
cc_264 N_B1_c_236_n N_Y_c_821_n 0.0138391f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_265 N_B1_c_236_n N_Y_c_822_n 0.0203132f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_266 N_B1_c_235_n N_A_508_368#_M1001_d 0.00205254f $X=3.29 $Y=1.615 $X2=-0.19
+ $Y2=-0.245
cc_267 N_B1_c_236_n N_A_508_368#_M1014_d 0.00198204f $X=5.405 $Y=1.795 $X2=0
+ $Y2=0
cc_268 N_B1_c_236_n N_A_508_368#_M1010_s 0.00198204f $X=5.405 $Y=1.795 $X2=0
+ $Y2=0
cc_269 N_B1_c_230_n N_A_508_368#_M1036_s 0.00259823f $X=5.835 $Y=1.515 $X2=0
+ $Y2=0
cc_270 N_B1_c_232_n N_A_508_368#_c_914_n 0.00947174f $X=2.915 $Y=1.765 $X2=0
+ $Y2=0
cc_271 N_B1_c_233_n N_A_508_368#_c_914_n 0.00947174f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_272 N_B1_c_233_n N_A_508_368#_c_916_n 4.27119e-19 $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_273 N_B1_c_232_n N_A_508_368#_c_917_n 5.5844e-19 $X=2.915 $Y=1.765 $X2=0
+ $Y2=0
cc_274 N_B1_c_233_n N_A_508_368#_c_917_n 0.00497909f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_275 N_B1_c_233_n N_A_508_368#_c_906_n 0.00313312f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_276 N_B1_c_227_n N_A_508_368#_c_907_n 0.0033071f $X=5.815 $Y=1.765 $X2=0
+ $Y2=0
cc_277 N_B1_c_227_n N_A_508_368#_c_921_n 0.00512366f $X=5.815 $Y=1.765 $X2=0
+ $Y2=0
cc_278 N_B1_c_231_n N_A_508_368#_c_908_n 0.00618929f $X=2.465 $Y=1.765 $X2=0
+ $Y2=0
cc_279 N_B1_c_232_n N_A_508_368#_c_908_n 0.00650056f $X=2.915 $Y=1.765 $X2=0
+ $Y2=0
cc_280 N_B1_c_233_n N_A_508_368#_c_908_n 5.73918e-19 $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_281 N_B1_M1008_g N_A_27_84#_c_1030_n 0.00288917f $X=2.775 $Y=0.74 $X2=0 $Y2=0
cc_282 N_B1_M1008_g N_A_27_84#_c_1031_n 0.00289242f $X=2.775 $Y=0.74 $X2=0 $Y2=0
cc_283 N_B1_M1008_g N_A_27_84#_c_1032_n 0.0206145f $X=2.775 $Y=0.74 $X2=0 $Y2=0
cc_284 N_B1_c_235_n N_A_27_84#_c_1032_n 0.040357f $X=3.29 $Y=1.615 $X2=0 $Y2=0
cc_285 N_B1_c_229_n N_A_27_84#_c_1032_n 0.0137245f $X=3.465 $Y=1.475 $X2=0 $Y2=0
cc_286 N_B1_c_224_n N_A_27_84#_c_1034_n 0.00841735f $X=3.205 $Y=1.185 $X2=0
+ $Y2=0
cc_287 N_B1_c_225_n N_A_27_84#_c_1034_n 0.00950816f $X=3.635 $Y=1.185 $X2=0
+ $Y2=0
cc_288 N_B1_c_236_n N_A_27_84#_c_1034_n 0.00395856f $X=5.405 $Y=1.795 $X2=0
+ $Y2=0
cc_289 N_B1_c_229_n N_A_27_84#_c_1034_n 0.00317182f $X=3.465 $Y=1.475 $X2=0
+ $Y2=0
cc_290 N_B1_c_224_n N_A_27_84#_c_1036_n 0.00558702f $X=3.205 $Y=1.185 $X2=0
+ $Y2=0
cc_291 N_B1_c_225_n N_A_27_84#_c_1036_n 5.18778e-19 $X=3.635 $Y=1.185 $X2=0
+ $Y2=0
cc_292 N_B1_c_228_n N_A_27_84#_c_1036_n 0.040357f $X=3.555 $Y=1.615 $X2=0 $Y2=0
cc_293 N_B1_c_224_n N_A_27_84#_c_1037_n 6.02585e-19 $X=3.205 $Y=1.185 $X2=0
+ $Y2=0
cc_294 N_B1_c_225_n N_A_27_84#_c_1037_n 0.00612157f $X=3.635 $Y=1.185 $X2=0
+ $Y2=0
cc_295 N_B1_c_236_n N_A_27_84#_c_1037_n 0.0111311f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_296 N_B1_M1035_g N_A_27_84#_c_1061_n 0.00364331f $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_297 N_B1_c_230_n N_A_27_84#_c_1061_n 0.0149317f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_298 N_B1_M1008_g N_A_483_74#_c_1107_n 0.0102979f $X=2.775 $Y=0.74 $X2=0 $Y2=0
cc_299 N_B1_c_224_n N_A_483_74#_c_1107_n 0.0113119f $X=3.205 $Y=1.185 $X2=0
+ $Y2=0
cc_300 N_B1_c_225_n N_A_483_74#_c_1108_n 0.0112282f $X=3.635 $Y=1.185 $X2=0
+ $Y2=0
cc_301 N_B1_M1035_g N_A_483_74#_c_1108_n 0.0154814f $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_302 N_B1_M1035_g N_A_483_74#_c_1114_n 6.56207e-19 $X=5.785 $Y=0.74 $X2=0
+ $Y2=0
cc_303 N_B1_c_227_n N_A_483_74#_c_1114_n 6.57592e-19 $X=5.815 $Y=1.765 $X2=0
+ $Y2=0
cc_304 N_B1_c_230_n N_A_483_74#_c_1114_n 0.00538446f $X=5.835 $Y=1.515 $X2=0
+ $Y2=0
cc_305 N_B1_M1008_g N_VGND_c_1221_n 0.00291649f $X=2.775 $Y=0.74 $X2=0 $Y2=0
cc_306 N_B1_c_224_n N_VGND_c_1221_n 0.00291649f $X=3.205 $Y=1.185 $X2=0 $Y2=0
cc_307 N_B1_c_225_n N_VGND_c_1221_n 0.00291649f $X=3.635 $Y=1.185 $X2=0 $Y2=0
cc_308 N_B1_M1035_g N_VGND_c_1221_n 0.00291649f $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_309 N_B1_M1008_g N_VGND_c_1226_n 0.0036412f $X=2.775 $Y=0.74 $X2=0 $Y2=0
cc_310 N_B1_c_224_n N_VGND_c_1226_n 0.00359121f $X=3.205 $Y=1.185 $X2=0 $Y2=0
cc_311 N_B1_c_225_n N_VGND_c_1226_n 0.00359219f $X=3.635 $Y=1.185 $X2=0 $Y2=0
cc_312 N_B1_M1035_g N_VGND_c_1226_n 0.0035993f $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_313 N_B2_c_351_n N_VPWR_c_643_n 0.00278257f $X=3.915 $Y=1.765 $X2=0 $Y2=0
cc_314 N_B2_c_352_n N_VPWR_c_643_n 0.00278257f $X=4.365 $Y=1.765 $X2=0 $Y2=0
cc_315 N_B2_c_353_n N_VPWR_c_643_n 0.00278257f $X=4.815 $Y=1.765 $X2=0 $Y2=0
cc_316 N_B2_c_354_n N_VPWR_c_643_n 0.00278271f $X=5.315 $Y=1.765 $X2=0 $Y2=0
cc_317 N_B2_c_351_n N_VPWR_c_630_n 0.00353905f $X=3.915 $Y=1.765 $X2=0 $Y2=0
cc_318 N_B2_c_352_n N_VPWR_c_630_n 0.00353822f $X=4.365 $Y=1.765 $X2=0 $Y2=0
cc_319 N_B2_c_353_n N_VPWR_c_630_n 0.00354283f $X=4.815 $Y=1.765 $X2=0 $Y2=0
cc_320 N_B2_c_354_n N_VPWR_c_630_n 0.00354798f $X=5.315 $Y=1.765 $X2=0 $Y2=0
cc_321 N_B2_c_351_n N_Y_c_795_n 0.0126036f $X=3.915 $Y=1.765 $X2=0 $Y2=0
cc_322 N_B2_c_351_n N_Y_c_824_n 0.0045686f $X=3.915 $Y=1.765 $X2=0 $Y2=0
cc_323 N_B2_c_352_n N_Y_c_824_n 0.00457102f $X=4.365 $Y=1.765 $X2=0 $Y2=0
cc_324 N_B2_c_352_n N_Y_c_815_n 0.0126853f $X=4.365 $Y=1.765 $X2=0 $Y2=0
cc_325 N_B2_c_353_n N_Y_c_815_n 0.0151589f $X=4.815 $Y=1.765 $X2=0 $Y2=0
cc_326 N_B2_c_354_n N_Y_c_816_n 0.00716255f $X=5.315 $Y=1.765 $X2=0 $Y2=0
cc_327 N_B2_c_354_n N_Y_c_817_n 0.01222f $X=5.315 $Y=1.765 $X2=0 $Y2=0
cc_328 N_B2_c_350_n N_Y_c_821_n 9.15927e-19 $X=5.315 $Y=1.492 $X2=0 $Y2=0
cc_329 N_B2_c_354_n N_Y_c_822_n 4.12619e-19 $X=5.315 $Y=1.765 $X2=0 $Y2=0
cc_330 N_B2_c_351_n N_A_508_368#_c_916_n 0.00193591f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_331 N_B2_c_351_n N_A_508_368#_c_917_n 0.00472645f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_332 N_B2_c_352_n N_A_508_368#_c_917_n 4.88744e-19 $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_333 N_B2_c_351_n N_A_508_368#_c_905_n 0.0108414f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_334 N_B2_c_352_n N_A_508_368#_c_905_n 0.0108414f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_335 N_B2_c_351_n N_A_508_368#_c_906_n 0.00171731f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_336 N_B2_c_351_n N_A_508_368#_c_931_n 5.40723e-19 $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_337 N_B2_c_352_n N_A_508_368#_c_931_n 0.00665026f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_338 N_B2_c_353_n N_A_508_368#_c_931_n 0.00673784f $X=4.815 $Y=1.765 $X2=0
+ $Y2=0
cc_339 N_B2_c_354_n N_A_508_368#_c_931_n 4.54023e-19 $X=5.315 $Y=1.765 $X2=0
+ $Y2=0
cc_340 N_B2_c_353_n N_A_508_368#_c_907_n 0.0111147f $X=4.815 $Y=1.765 $X2=0
+ $Y2=0
cc_341 N_B2_c_354_n N_A_508_368#_c_907_n 0.0140663f $X=5.315 $Y=1.765 $X2=0
+ $Y2=0
cc_342 N_B2_c_352_n N_A_508_368#_c_909_n 0.00174703f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_343 N_B2_c_353_n N_A_508_368#_c_909_n 0.00174703f $X=4.815 $Y=1.765 $X2=0
+ $Y2=0
cc_344 N_B2_c_345_n N_A_27_84#_c_1037_n 0.00612289f $X=4.065 $Y=1.22 $X2=0 $Y2=0
cc_345 N_B2_c_346_n N_A_27_84#_c_1037_n 9.42328e-19 $X=4.495 $Y=1.22 $X2=0 $Y2=0
cc_346 N_B2_c_350_n N_A_27_84#_c_1037_n 0.00387271f $X=5.315 $Y=1.492 $X2=0
+ $Y2=0
cc_347 N_B2_c_348_n N_A_27_84#_c_1061_n 0.00202711f $X=5.355 $Y=1.22 $X2=0 $Y2=0
cc_348 N_B2_c_345_n N_A_27_84#_c_1067_n 0.0138321f $X=4.065 $Y=1.22 $X2=0 $Y2=0
cc_349 N_B2_c_346_n N_A_27_84#_c_1067_n 0.0103131f $X=4.495 $Y=1.22 $X2=0 $Y2=0
cc_350 N_B2_c_347_n N_A_27_84#_c_1067_n 0.0103131f $X=4.925 $Y=1.22 $X2=0 $Y2=0
cc_351 N_B2_c_348_n N_A_27_84#_c_1067_n 0.0130444f $X=5.355 $Y=1.22 $X2=0 $Y2=0
cc_352 B2 N_A_27_84#_c_1067_n 0.0699825f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_353 N_B2_c_350_n N_A_27_84#_c_1067_n 0.00192623f $X=5.315 $Y=1.492 $X2=0
+ $Y2=0
cc_354 N_B2_c_345_n N_A_483_74#_c_1108_n 0.0101343f $X=4.065 $Y=1.22 $X2=0 $Y2=0
cc_355 N_B2_c_346_n N_A_483_74#_c_1108_n 0.010218f $X=4.495 $Y=1.22 $X2=0 $Y2=0
cc_356 N_B2_c_347_n N_A_483_74#_c_1108_n 0.010218f $X=4.925 $Y=1.22 $X2=0 $Y2=0
cc_357 N_B2_c_348_n N_A_483_74#_c_1108_n 0.0101492f $X=5.355 $Y=1.22 $X2=0 $Y2=0
cc_358 N_B2_c_345_n N_VGND_c_1221_n 0.00291649f $X=4.065 $Y=1.22 $X2=0 $Y2=0
cc_359 N_B2_c_346_n N_VGND_c_1221_n 0.00291649f $X=4.495 $Y=1.22 $X2=0 $Y2=0
cc_360 N_B2_c_347_n N_VGND_c_1221_n 0.00291649f $X=4.925 $Y=1.22 $X2=0 $Y2=0
cc_361 N_B2_c_348_n N_VGND_c_1221_n 0.00291649f $X=5.355 $Y=1.22 $X2=0 $Y2=0
cc_362 N_B2_c_345_n N_VGND_c_1226_n 0.00358272f $X=4.065 $Y=1.22 $X2=0 $Y2=0
cc_363 N_B2_c_346_n N_VGND_c_1226_n 0.00359121f $X=4.495 $Y=1.22 $X2=0 $Y2=0
cc_364 N_B2_c_347_n N_VGND_c_1226_n 0.00359121f $X=4.925 $Y=1.22 $X2=0 $Y2=0
cc_365 N_B2_c_348_n N_VGND_c_1226_n 0.00359219f $X=5.355 $Y=1.22 $X2=0 $Y2=0
cc_366 N_A1_M1005_g N_A2_M1004_g 0.0240526f $X=6.285 $Y=0.74 $X2=0 $Y2=0
cc_367 N_A1_c_429_n N_A2_M1004_g 0.0179795f $X=6.365 $Y=1.765 $X2=0 $Y2=0
cc_368 N_A1_c_433_n N_A2_M1004_g 0.00517694f $X=6.575 $Y=1.175 $X2=0 $Y2=0
cc_369 N_A1_c_436_n N_A2_M1004_g 0.0128429f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_370 N_A1_c_429_n N_A2_c_549_n 0.0384825f $X=6.365 $Y=1.765 $X2=0 $Y2=0
cc_371 N_A1_c_436_n N_A2_M1011_g 0.0108858f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_372 N_A1_c_436_n N_A2_M1018_g 0.0108382f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_373 N_A1_c_437_n N_A2_M1018_g 4.14448e-19 $X=8.455 $Y=1.435 $X2=0 $Y2=0
cc_374 N_A1_M1029_g N_A2_M1022_g 0.0206073f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_375 N_A1_c_436_n N_A2_M1022_g 0.0104871f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_376 N_A1_c_437_n N_A2_M1022_g 0.00421415f $X=8.455 $Y=1.435 $X2=0 $Y2=0
cc_377 N_A1_c_439_n N_A2_c_552_n 0.0121151f $X=8.67 $Y=1.765 $X2=0 $Y2=0
cc_378 N_A1_c_437_n N_A2_c_552_n 8.12167e-19 $X=8.455 $Y=1.435 $X2=0 $Y2=0
cc_379 N_A1_c_429_n A2 0.0011864f $X=6.365 $Y=1.765 $X2=0 $Y2=0
cc_380 N_A1_c_433_n A2 0.00953035f $X=6.575 $Y=1.175 $X2=0 $Y2=0
cc_381 N_A1_c_436_n A2 0.0884035f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_382 N_A1_c_437_n A2 0.0220095f $X=8.455 $Y=1.435 $X2=0 $Y2=0
cc_383 N_A1_c_429_n N_A2_c_548_n 0.00742447f $X=6.365 $Y=1.765 $X2=0 $Y2=0
cc_384 N_A1_c_435_n N_A2_c_548_n 0.0317746f $X=9.57 $Y=1.512 $X2=0 $Y2=0
cc_385 N_A1_c_436_n N_A2_c_548_n 0.00936448f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_386 N_A1_c_437_n N_A2_c_548_n 0.0157984f $X=8.455 $Y=1.435 $X2=0 $Y2=0
cc_387 N_A1_c_429_n N_VPWR_c_636_n 0.00487422f $X=6.365 $Y=1.765 $X2=0 $Y2=0
cc_388 N_A1_c_439_n N_VPWR_c_637_n 0.00996098f $X=8.67 $Y=1.765 $X2=0 $Y2=0
cc_389 N_A1_c_440_n N_VPWR_c_637_n 0.00526215f $X=9.12 $Y=1.765 $X2=0 $Y2=0
cc_390 N_A1_c_441_n N_VPWR_c_639_n 0.00831454f $X=9.57 $Y=1.765 $X2=0 $Y2=0
cc_391 A1 N_VPWR_c_639_n 0.0219047f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_392 N_A1_c_429_n N_VPWR_c_644_n 0.0044313f $X=6.365 $Y=1.765 $X2=0 $Y2=0
cc_393 N_A1_c_439_n N_VPWR_c_644_n 0.00413917f $X=8.67 $Y=1.765 $X2=0 $Y2=0
cc_394 N_A1_c_440_n N_VPWR_c_645_n 0.00445602f $X=9.12 $Y=1.765 $X2=0 $Y2=0
cc_395 N_A1_c_441_n N_VPWR_c_645_n 0.00445602f $X=9.57 $Y=1.765 $X2=0 $Y2=0
cc_396 N_A1_c_429_n N_VPWR_c_630_n 0.00854152f $X=6.365 $Y=1.765 $X2=0 $Y2=0
cc_397 N_A1_c_439_n N_VPWR_c_630_n 0.0081781f $X=8.67 $Y=1.765 $X2=0 $Y2=0
cc_398 N_A1_c_440_n N_VPWR_c_630_n 0.00857589f $X=9.12 $Y=1.765 $X2=0 $Y2=0
cc_399 N_A1_c_441_n N_VPWR_c_630_n 0.008611f $X=9.57 $Y=1.765 $X2=0 $Y2=0
cc_400 N_A1_c_429_n N_Y_c_817_n 0.0177355f $X=6.365 $Y=1.765 $X2=0 $Y2=0
cc_401 N_A1_c_433_n N_Y_c_817_n 0.0104999f $X=6.575 $Y=1.175 $X2=0 $Y2=0
cc_402 N_A1_c_429_n Y 0.00224232f $X=6.365 $Y=1.765 $X2=0 $Y2=0
cc_403 N_A1_c_439_n N_A_1288_368#_c_973_n 0.00125031f $X=8.67 $Y=1.765 $X2=0
+ $Y2=0
cc_404 N_A1_c_437_n N_A_1288_368#_c_978_n 0.0153836f $X=8.455 $Y=1.435 $X2=0
+ $Y2=0
cc_405 N_A1_c_439_n N_A_1288_368#_c_979_n 0.0126853f $X=8.67 $Y=1.765 $X2=0
+ $Y2=0
cc_406 N_A1_c_440_n N_A_1288_368#_c_979_n 0.0119563f $X=9.12 $Y=1.765 $X2=0
+ $Y2=0
cc_407 A1 N_A_1288_368#_c_979_n 0.0443416f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_408 N_A1_c_435_n N_A_1288_368#_c_979_n 0.00108122f $X=9.57 $Y=1.512 $X2=0
+ $Y2=0
cc_409 N_A1_c_440_n N_A_1288_368#_c_983_n 4.27055e-19 $X=9.12 $Y=1.765 $X2=0
+ $Y2=0
cc_410 N_A1_c_441_n N_A_1288_368#_c_983_n 0.00203651f $X=9.57 $Y=1.765 $X2=0
+ $Y2=0
cc_411 A1 N_A_1288_368#_c_983_n 0.0241747f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_412 N_A1_c_435_n N_A_1288_368#_c_983_n 0.00118928f $X=9.57 $Y=1.512 $X2=0
+ $Y2=0
cc_413 N_A1_c_439_n N_A_1288_368#_c_974_n 6.69308e-19 $X=8.67 $Y=1.765 $X2=0
+ $Y2=0
cc_414 N_A1_c_440_n N_A_1288_368#_c_974_n 0.0105452f $X=9.12 $Y=1.765 $X2=0
+ $Y2=0
cc_415 N_A1_c_441_n N_A_1288_368#_c_974_n 0.00960826f $X=9.57 $Y=1.765 $X2=0
+ $Y2=0
cc_416 N_A1_c_429_n N_A_1288_368#_c_975_n 0.00612074f $X=6.365 $Y=1.765 $X2=0
+ $Y2=0
cc_417 N_A1_c_436_n N_A_483_74#_M1004_s 0.00176461f $X=8.285 $Y=1.435 $X2=0
+ $Y2=0
cc_418 N_A1_c_436_n N_A_483_74#_M1018_s 0.00176461f $X=8.285 $Y=1.435 $X2=0
+ $Y2=0
cc_419 N_A1_M1005_g N_A_483_74#_c_1129_n 0.0107566f $X=6.285 $Y=0.74 $X2=0 $Y2=0
cc_420 N_A1_c_429_n N_A_483_74#_c_1129_n 6.10063e-19 $X=6.365 $Y=1.765 $X2=0
+ $Y2=0
cc_421 N_A1_c_433_n N_A_483_74#_c_1129_n 0.0186469f $X=6.575 $Y=1.175 $X2=0
+ $Y2=0
cc_422 N_A1_c_436_n N_A_483_74#_c_1129_n 0.0195621f $X=8.285 $Y=1.435 $X2=0
+ $Y2=0
cc_423 N_A1_M1005_g N_A_483_74#_c_1109_n 5.78282e-19 $X=6.285 $Y=0.74 $X2=0
+ $Y2=0
cc_424 N_A1_c_436_n N_A_483_74#_c_1134_n 0.0357472f $X=8.285 $Y=1.435 $X2=0
+ $Y2=0
cc_425 N_A1_M1029_g N_A_483_74#_c_1135_n 0.0118367f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_426 A1 N_A_483_74#_c_1135_n 0.0123244f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_427 N_A1_c_436_n N_A_483_74#_c_1135_n 0.019324f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_428 N_A1_M1029_g N_A_483_74#_c_1111_n 0.00214936f $X=8.655 $Y=0.74 $X2=0
+ $Y2=0
cc_429 N_A1_M1031_g N_A_483_74#_c_1111_n 2.6509e-19 $X=9.155 $Y=0.74 $X2=0 $Y2=0
cc_430 N_A1_M1031_g N_A_483_74#_c_1112_n 0.0122595f $X=9.155 $Y=0.74 $X2=0 $Y2=0
cc_431 N_A1_M1034_g N_A_483_74#_c_1112_n 0.0122129f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_432 A1 N_A_483_74#_c_1112_n 0.0655704f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_433 N_A1_c_435_n N_A_483_74#_c_1112_n 0.00224206f $X=9.57 $Y=1.512 $X2=0
+ $Y2=0
cc_434 N_A1_M1034_g N_A_483_74#_c_1113_n 8.26992e-19 $X=9.585 $Y=0.74 $X2=0
+ $Y2=0
cc_435 N_A1_M1005_g N_A_483_74#_c_1114_n 0.0112264f $X=6.285 $Y=0.74 $X2=0 $Y2=0
cc_436 N_A1_c_433_n N_A_483_74#_c_1114_n 0.00188346f $X=6.575 $Y=1.175 $X2=0
+ $Y2=0
cc_437 N_A1_c_436_n N_A_483_74#_c_1147_n 0.0151907f $X=8.285 $Y=1.435 $X2=0
+ $Y2=0
cc_438 N_A1_c_436_n N_A_483_74#_c_1148_n 0.0151907f $X=8.285 $Y=1.435 $X2=0
+ $Y2=0
cc_439 A1 N_A_483_74#_c_1149_n 0.0206148f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_440 N_A1_c_435_n N_A_483_74#_c_1149_n 0.00396026f $X=9.57 $Y=1.512 $X2=0
+ $Y2=0
cc_441 N_A1_c_433_n N_VGND_M1005_s 0.0017364f $X=6.575 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_442 N_A1_c_436_n N_VGND_M1005_s 0.00158921f $X=8.285 $Y=1.435 $X2=-0.19
+ $Y2=-0.245
cc_443 N_A1_c_436_n N_VGND_M1011_d 0.00251484f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_444 N_A1_c_437_n N_VGND_M1022_d 0.00145497f $X=8.455 $Y=1.435 $X2=0 $Y2=0
cc_445 N_A1_M1005_g N_VGND_c_1217_n 0.00464693f $X=6.285 $Y=0.74 $X2=0 $Y2=0
cc_446 N_A1_M1029_g N_VGND_c_1219_n 0.00679571f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_447 N_A1_M1031_g N_VGND_c_1219_n 3.92591e-19 $X=9.155 $Y=0.74 $X2=0 $Y2=0
cc_448 N_A1_M1029_g N_VGND_c_1220_n 4.37937e-19 $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_449 N_A1_M1031_g N_VGND_c_1220_n 0.00869262f $X=9.155 $Y=0.74 $X2=0 $Y2=0
cc_450 N_A1_M1034_g N_VGND_c_1220_n 0.0114756f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_451 N_A1_M1005_g N_VGND_c_1221_n 0.00331438f $X=6.285 $Y=0.74 $X2=0 $Y2=0
cc_452 N_A1_M1029_g N_VGND_c_1224_n 0.00281141f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_453 N_A1_M1031_g N_VGND_c_1224_n 0.00383152f $X=9.155 $Y=0.74 $X2=0 $Y2=0
cc_454 N_A1_M1034_g N_VGND_c_1225_n 0.00383152f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_455 N_A1_M1005_g N_VGND_c_1226_n 0.0042805f $X=6.285 $Y=0.74 $X2=0 $Y2=0
cc_456 N_A1_M1029_g N_VGND_c_1226_n 0.00365724f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_457 N_A1_M1031_g N_VGND_c_1226_n 0.00758198f $X=9.155 $Y=0.74 $X2=0 $Y2=0
cc_458 N_A1_M1034_g N_VGND_c_1226_n 0.00761198f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_459 N_A2_c_549_n N_VPWR_c_644_n 0.00278271f $X=6.87 $Y=1.765 $X2=0 $Y2=0
cc_460 N_A2_c_550_n N_VPWR_c_644_n 0.00278271f $X=7.32 $Y=1.765 $X2=0 $Y2=0
cc_461 N_A2_c_551_n N_VPWR_c_644_n 0.00278271f $X=7.77 $Y=1.765 $X2=0 $Y2=0
cc_462 N_A2_c_552_n N_VPWR_c_644_n 0.00278271f $X=8.22 $Y=1.765 $X2=0 $Y2=0
cc_463 N_A2_c_549_n N_VPWR_c_630_n 0.00354378f $X=6.87 $Y=1.765 $X2=0 $Y2=0
cc_464 N_A2_c_550_n N_VPWR_c_630_n 0.00353823f $X=7.32 $Y=1.765 $X2=0 $Y2=0
cc_465 N_A2_c_551_n N_VPWR_c_630_n 0.00353823f $X=7.77 $Y=1.765 $X2=0 $Y2=0
cc_466 N_A2_c_552_n N_VPWR_c_630_n 0.00353907f $X=8.22 $Y=1.765 $X2=0 $Y2=0
cc_467 N_A2_c_549_n N_Y_c_817_n 0.00747335f $X=6.87 $Y=1.765 $X2=0 $Y2=0
cc_468 N_A2_c_550_n N_Y_c_836_n 0.0120074f $X=7.32 $Y=1.765 $X2=0 $Y2=0
cc_469 N_A2_c_551_n N_Y_c_836_n 0.0120074f $X=7.77 $Y=1.765 $X2=0 $Y2=0
cc_470 A2 N_Y_c_836_n 0.0386622f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_471 N_A2_c_548_n N_Y_c_836_n 0.00131353f $X=8.215 $Y=1.557 $X2=0 $Y2=0
cc_472 N_A2_c_550_n N_Y_c_840_n 5.70931e-19 $X=7.32 $Y=1.765 $X2=0 $Y2=0
cc_473 N_A2_c_551_n N_Y_c_840_n 0.0089154f $X=7.77 $Y=1.765 $X2=0 $Y2=0
cc_474 N_A2_c_552_n N_Y_c_840_n 0.00968337f $X=8.22 $Y=1.765 $X2=0 $Y2=0
cc_475 A2 N_Y_c_840_n 0.0151443f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_476 N_A2_c_548_n N_Y_c_840_n 0.00413059f $X=8.215 $Y=1.557 $X2=0 $Y2=0
cc_477 N_A2_c_549_n Y 0.0195004f $X=6.87 $Y=1.765 $X2=0 $Y2=0
cc_478 N_A2_c_550_n Y 0.00897905f $X=7.32 $Y=1.765 $X2=0 $Y2=0
cc_479 N_A2_c_551_n Y 5.70045e-19 $X=7.77 $Y=1.765 $X2=0 $Y2=0
cc_480 A2 Y 0.0300427f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_481 N_A2_c_548_n Y 0.00144162f $X=8.215 $Y=1.557 $X2=0 $Y2=0
cc_482 N_A2_c_549_n N_A_1288_368#_c_972_n 0.0118458f $X=6.87 $Y=1.765 $X2=0
+ $Y2=0
cc_483 N_A2_c_550_n N_A_1288_368#_c_972_n 0.0128043f $X=7.32 $Y=1.765 $X2=0
+ $Y2=0
cc_484 N_A2_c_551_n N_A_1288_368#_c_973_n 0.0127839f $X=7.77 $Y=1.765 $X2=0
+ $Y2=0
cc_485 N_A2_c_552_n N_A_1288_368#_c_973_n 0.012504f $X=8.22 $Y=1.765 $X2=0 $Y2=0
cc_486 N_A2_c_549_n N_A_1288_368#_c_975_n 6.69206e-19 $X=6.87 $Y=1.765 $X2=0
+ $Y2=0
cc_487 N_A2_M1004_g N_A_483_74#_c_1129_n 0.00941575f $X=6.855 $Y=0.74 $X2=0
+ $Y2=0
cc_488 N_A2_M1004_g N_A_483_74#_c_1109_n 0.00687331f $X=6.855 $Y=0.74 $X2=0
+ $Y2=0
cc_489 N_A2_M1011_g N_A_483_74#_c_1109_n 4.39567e-19 $X=7.285 $Y=0.74 $X2=0
+ $Y2=0
cc_490 N_A2_M1011_g N_A_483_74#_c_1134_n 0.0113092f $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_491 N_A2_M1018_g N_A_483_74#_c_1134_n 0.00916065f $X=7.785 $Y=0.74 $X2=0
+ $Y2=0
cc_492 N_A2_M1011_g N_A_483_74#_c_1110_n 6.09957e-19 $X=7.285 $Y=0.74 $X2=0
+ $Y2=0
cc_493 N_A2_M1018_g N_A_483_74#_c_1110_n 0.00657942f $X=7.785 $Y=0.74 $X2=0
+ $Y2=0
cc_494 N_A2_M1022_g N_A_483_74#_c_1110_n 4.39567e-19 $X=8.215 $Y=0.74 $X2=0
+ $Y2=0
cc_495 N_A2_M1022_g N_A_483_74#_c_1135_n 0.0109279f $X=8.215 $Y=0.74 $X2=0 $Y2=0
cc_496 N_A2_M1004_g N_A_483_74#_c_1114_n 0.00144055f $X=6.855 $Y=0.74 $X2=0
+ $Y2=0
cc_497 N_A2_M1004_g N_A_483_74#_c_1147_n 0.00181289f $X=6.855 $Y=0.74 $X2=0
+ $Y2=0
cc_498 N_A2_M1018_g N_A_483_74#_c_1148_n 0.00181289f $X=7.785 $Y=0.74 $X2=0
+ $Y2=0
cc_499 N_A2_M1004_g N_VGND_c_1217_n 0.00317556f $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_500 N_A2_M1004_g N_VGND_c_1218_n 4.44774e-19 $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_501 N_A2_M1011_g N_VGND_c_1218_n 0.00678063f $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_502 N_A2_M1018_g N_VGND_c_1218_n 0.0028836f $X=7.785 $Y=0.74 $X2=0 $Y2=0
cc_503 N_A2_M1018_g N_VGND_c_1219_n 4.44681e-19 $X=7.785 $Y=0.74 $X2=0 $Y2=0
cc_504 N_A2_M1022_g N_VGND_c_1219_n 0.00678207f $X=8.215 $Y=0.74 $X2=0 $Y2=0
cc_505 N_A2_M1004_g N_VGND_c_1222_n 0.00331438f $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_506 N_A2_M1011_g N_VGND_c_1222_n 0.00281141f $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_507 N_A2_M1018_g N_VGND_c_1223_n 0.00331438f $X=7.785 $Y=0.74 $X2=0 $Y2=0
cc_508 N_A2_M1022_g N_VGND_c_1223_n 0.00281141f $X=8.215 $Y=0.74 $X2=0 $Y2=0
cc_509 N_A2_M1004_g N_VGND_c_1226_n 0.00427339f $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_510 N_A2_M1011_g N_VGND_c_1226_n 0.00365066f $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_511 N_A2_M1018_g N_VGND_c_1226_n 0.00426745f $X=7.785 $Y=0.74 $X2=0 $Y2=0
cc_512 N_A2_M1022_g N_VGND_c_1226_n 0.00365066f $X=8.215 $Y=0.74 $X2=0 $Y2=0
cc_513 N_VPWR_c_632_n N_Y_c_772_n 0.0121024f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_514 N_VPWR_c_632_n N_Y_c_765_n 0.0576605f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_515 N_VPWR_c_633_n N_Y_c_765_n 0.0266809f $X=1.23 $Y=2.455 $X2=0 $Y2=0
cc_516 N_VPWR_c_640_n N_Y_c_765_n 0.014552f $X=1.065 $Y=3.33 $X2=0 $Y2=0
cc_517 N_VPWR_c_630_n N_Y_c_765_n 0.0119791f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_518 N_VPWR_M1023_s N_Y_c_787_n 0.00546838f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_519 N_VPWR_c_633_n N_Y_c_787_n 0.0220482f $X=1.23 $Y=2.455 $X2=0 $Y2=0
cc_520 N_VPWR_c_633_n N_Y_c_766_n 0.00148713f $X=1.23 $Y=2.455 $X2=0 $Y2=0
cc_521 N_VPWR_c_634_n N_Y_c_766_n 0.0395897f $X=2.19 $Y=2.475 $X2=0 $Y2=0
cc_522 N_VPWR_c_641_n N_Y_c_766_n 0.011066f $X=2.025 $Y=3.33 $X2=0 $Y2=0
cc_523 N_VPWR_c_630_n N_Y_c_766_n 0.00915947f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_524 N_VPWR_M1032_s N_Y_c_795_n 0.0115134f $X=2.04 $Y=1.84 $X2=0 $Y2=0
cc_525 N_VPWR_M1012_s N_Y_c_795_n 0.00600628f $X=2.99 $Y=1.84 $X2=0 $Y2=0
cc_526 N_VPWR_c_634_n N_Y_c_795_n 0.0202249f $X=2.19 $Y=2.475 $X2=0 $Y2=0
cc_527 N_VPWR_M1016_s N_Y_c_817_n 0.0122639f $X=5.89 $Y=1.84 $X2=0 $Y2=0
cc_528 N_VPWR_c_636_n N_Y_c_817_n 0.0232685f $X=6.09 $Y=2.475 $X2=0 $Y2=0
cc_529 N_VPWR_M1012_s N_A_508_368#_c_914_n 0.00639987f $X=2.99 $Y=1.84 $X2=0
+ $Y2=0
cc_530 N_VPWR_c_635_n N_A_508_368#_c_914_n 0.0226192f $X=3.19 $Y=2.815 $X2=0
+ $Y2=0
cc_531 N_VPWR_c_630_n N_A_508_368#_c_914_n 0.0117498f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_532 N_VPWR_c_643_n N_A_508_368#_c_905_n 0.03588f $X=5.925 $Y=3.33 $X2=0 $Y2=0
cc_533 N_VPWR_c_630_n N_A_508_368#_c_905_n 0.0201952f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_635_n N_A_508_368#_c_906_n 0.0119239f $X=3.19 $Y=2.815 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_643_n N_A_508_368#_c_906_n 0.0235643f $X=5.925 $Y=3.33 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_630_n N_A_508_368#_c_906_n 0.0126949f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_636_n N_A_508_368#_c_907_n 0.0119239f $X=6.09 $Y=2.475 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_643_n N_A_508_368#_c_907_n 0.0658922f $X=5.925 $Y=3.33 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_630_n N_A_508_368#_c_907_n 0.0366496f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_634_n N_A_508_368#_c_908_n 0.0165124f $X=2.19 $Y=2.475 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_635_n N_A_508_368#_c_908_n 0.0101711f $X=3.19 $Y=2.815 $X2=0
+ $Y2=0
cc_542 N_VPWR_c_642_n N_A_508_368#_c_908_n 0.0144033f $X=3.025 $Y=3.33 $X2=0
+ $Y2=0
cc_543 N_VPWR_c_630_n N_A_508_368#_c_908_n 0.0119211f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_643_n N_A_508_368#_c_909_n 0.0235642f $X=5.925 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_630_n N_A_508_368#_c_909_n 0.0126948f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_644_n N_A_1288_368#_c_972_n 0.0441612f $X=8.73 $Y=3.33 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_630_n N_A_1288_368#_c_972_n 0.0249452f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_637_n N_A_1288_368#_c_973_n 0.0123543f $X=8.895 $Y=2.455 $X2=0
+ $Y2=0
cc_549 N_VPWR_c_644_n N_A_1288_368#_c_973_n 0.0582805f $X=8.73 $Y=3.33 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_630_n N_A_1288_368#_c_973_n 0.0326824f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_637_n N_A_1288_368#_c_1001_n 0.039183f $X=8.895 $Y=2.455 $X2=0
+ $Y2=0
cc_552 N_VPWR_M1020_s N_A_1288_368#_c_979_n 0.00390065f $X=8.745 $Y=1.84 $X2=0
+ $Y2=0
cc_553 N_VPWR_c_637_n N_A_1288_368#_c_979_n 0.0154248f $X=8.895 $Y=2.455 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_639_n N_A_1288_368#_c_983_n 0.0121024f $X=9.795 $Y=2.115 $X2=0
+ $Y2=0
cc_555 N_VPWR_c_637_n N_A_1288_368#_c_974_n 0.0462948f $X=8.895 $Y=2.455 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_639_n N_A_1288_368#_c_974_n 0.0576605f $X=9.795 $Y=2.115 $X2=0
+ $Y2=0
cc_557 N_VPWR_c_645_n N_A_1288_368#_c_974_n 0.014552f $X=9.71 $Y=3.33 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_630_n N_A_1288_368#_c_974_n 0.0119791f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_636_n N_A_1288_368#_c_975_n 0.0214367f $X=6.09 $Y=2.475 $X2=0
+ $Y2=0
cc_560 N_VPWR_c_644_n N_A_1288_368#_c_975_n 0.0230495f $X=8.73 $Y=3.33 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_630_n N_A_1288_368#_c_975_n 0.0127846f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_562 N_VPWR_c_644_n N_A_1288_368#_c_976_n 0.0121867f $X=8.73 $Y=3.33 $X2=0
+ $Y2=0
cc_563 N_VPWR_c_630_n N_A_1288_368#_c_976_n 0.00660921f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_564 N_Y_c_795_n N_A_508_368#_M1001_d 0.00365946f $X=4.055 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_565 N_Y_c_795_n N_A_508_368#_M1014_d 0.00395925f $X=4.055 $Y=2.135 $X2=0
+ $Y2=0
cc_566 N_Y_c_815_n N_A_508_368#_M1010_s 0.00385254f $X=4.925 $Y=2.135 $X2=0
+ $Y2=0
cc_567 N_Y_c_817_n N_A_508_368#_M1036_s 0.00499657f $X=6.845 $Y=2.135 $X2=0
+ $Y2=0
cc_568 N_Y_c_795_n N_A_508_368#_c_914_n 0.039006f $X=4.055 $Y=2.135 $X2=0 $Y2=0
cc_569 N_Y_c_795_n N_A_508_368#_c_916_n 0.0173441f $X=4.055 $Y=2.135 $X2=0 $Y2=0
cc_570 N_Y_c_824_n N_A_508_368#_c_916_n 0.0117758f $X=4.14 $Y=2.57 $X2=0 $Y2=0
cc_571 N_Y_c_824_n N_A_508_368#_c_917_n 0.011366f $X=4.14 $Y=2.57 $X2=0 $Y2=0
cc_572 N_Y_M1006_d N_A_508_368#_c_905_n 0.00247267f $X=3.99 $Y=1.84 $X2=0 $Y2=0
cc_573 N_Y_c_824_n N_A_508_368#_c_905_n 0.0127942f $X=4.14 $Y=2.57 $X2=0 $Y2=0
cc_574 N_Y_c_824_n N_A_508_368#_c_931_n 0.0224722f $X=4.14 $Y=2.57 $X2=0 $Y2=0
cc_575 N_Y_c_815_n N_A_508_368#_c_931_n 0.0171916f $X=4.925 $Y=2.135 $X2=0 $Y2=0
cc_576 N_Y_M1026_d N_A_508_368#_c_907_n 0.00250873f $X=4.89 $Y=1.84 $X2=0 $Y2=0
cc_577 N_Y_c_816_n N_A_508_368#_c_907_n 0.0189337f $X=5.09 $Y=2.57 $X2=0 $Y2=0
cc_578 N_Y_c_817_n N_A_508_368#_c_921_n 0.0202371f $X=6.845 $Y=2.135 $X2=0 $Y2=0
cc_579 N_Y_c_795_n N_A_508_368#_c_908_n 0.0171364f $X=4.055 $Y=2.135 $X2=0 $Y2=0
cc_580 N_Y_c_817_n N_A_1288_368#_M1019_d 0.0115555f $X=6.845 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_581 N_Y_c_836_n N_A_1288_368#_M1013_s 0.00408911f $X=7.83 $Y=2.035 $X2=0
+ $Y2=0
cc_582 N_Y_M1007_d N_A_1288_368#_c_972_n 0.00197722f $X=6.945 $Y=1.84 $X2=0
+ $Y2=0
cc_583 Y N_A_1288_368#_c_972_n 0.0190187f $X=6.875 $Y=2.32 $X2=0 $Y2=0
cc_584 N_Y_c_836_n N_A_1288_368#_c_1018_n 0.0136682f $X=7.83 $Y=2.035 $X2=0
+ $Y2=0
cc_585 N_Y_c_840_n N_A_1288_368#_c_1018_n 0.0289859f $X=7.995 $Y=2.115 $X2=0
+ $Y2=0
cc_586 Y N_A_1288_368#_c_1018_n 0.0293817f $X=6.875 $Y=2.32 $X2=0 $Y2=0
cc_587 N_Y_M1027_d N_A_1288_368#_c_973_n 0.00197722f $X=7.845 $Y=1.84 $X2=0
+ $Y2=0
cc_588 N_Y_c_840_n N_A_1288_368#_c_973_n 0.0160777f $X=7.995 $Y=2.115 $X2=0
+ $Y2=0
cc_589 N_Y_c_840_n N_A_1288_368#_c_978_n 0.013092f $X=7.995 $Y=2.115 $X2=0 $Y2=0
cc_590 N_Y_c_840_n N_A_1288_368#_c_1001_n 0.039994f $X=7.995 $Y=2.115 $X2=0
+ $Y2=0
cc_591 N_Y_c_817_n N_A_1288_368#_c_975_n 0.00966092f $X=6.845 $Y=2.135 $X2=0
+ $Y2=0
cc_592 Y N_A_1288_368#_c_975_n 0.0044854f $X=6.875 $Y=2.32 $X2=0 $Y2=0
cc_593 N_Y_c_761_n N_A_27_84#_M1021_s 0.00176461f $X=1.405 $Y=1.095 $X2=0 $Y2=0
cc_594 N_Y_c_762_n N_A_27_84#_c_1027_n 0.00792678f $X=0.875 $Y=1.095 $X2=0 $Y2=0
cc_595 N_Y_M1000_d N_A_27_84#_c_1028_n 0.00176461f $X=0.57 $Y=0.42 $X2=0 $Y2=0
cc_596 N_Y_c_769_n N_A_27_84#_c_1028_n 0.0157965f $X=0.71 $Y=0.68 $X2=0 $Y2=0
cc_597 N_Y_c_761_n N_A_27_84#_c_1028_n 0.00304353f $X=1.405 $Y=1.095 $X2=0 $Y2=0
cc_598 N_Y_c_761_n N_A_27_84#_c_1078_n 0.0133411f $X=1.405 $Y=1.095 $X2=0 $Y2=0
cc_599 N_Y_M1038_d N_A_27_84#_c_1030_n 0.00176461f $X=1.43 $Y=0.42 $X2=0 $Y2=0
cc_600 N_Y_c_761_n N_A_27_84#_c_1030_n 0.00304353f $X=1.405 $Y=1.095 $X2=0 $Y2=0
cc_601 N_Y_c_791_n N_A_27_84#_c_1030_n 0.0165966f $X=1.57 $Y=0.68 $X2=0 $Y2=0
cc_602 N_Y_c_763_n N_A_27_84#_c_1033_n 0.00808484f $X=1.575 $Y=1.095 $X2=0 $Y2=0
cc_603 N_A_27_84#_c_1032_n N_A_483_74#_M1008_s 0.00441709f $X=2.95 $Y=0.975
+ $X2=-0.19 $Y2=-0.245
cc_604 N_A_27_84#_c_1034_n N_A_483_74#_M1009_s 0.00176461f $X=3.685 $Y=1.095
+ $X2=0 $Y2=0
cc_605 N_A_27_84#_c_1067_n N_A_483_74#_M1003_d 0.00332127f $X=5.405 $Y=0.91
+ $X2=0 $Y2=0
cc_606 N_A_27_84#_c_1067_n N_A_483_74#_M1017_d 0.00413357f $X=5.405 $Y=0.91
+ $X2=0 $Y2=0
cc_607 N_A_27_84#_M1008_d N_A_483_74#_c_1107_n 0.00179007f $X=2.85 $Y=0.37 $X2=0
+ $Y2=0
cc_608 N_A_27_84#_c_1030_n N_A_483_74#_c_1107_n 0.00560069f $X=1.915 $Y=0.34
+ $X2=0 $Y2=0
cc_609 N_A_27_84#_c_1031_n N_A_483_74#_c_1107_n 0.0121732f $X=2 $Y=0.565 $X2=0
+ $Y2=0
cc_610 N_A_27_84#_c_1032_n N_A_483_74#_c_1107_n 0.0445249f $X=2.95 $Y=0.975
+ $X2=0 $Y2=0
cc_611 N_A_27_84#_c_1034_n N_A_483_74#_c_1107_n 0.0174102f $X=3.685 $Y=1.095
+ $X2=0 $Y2=0
cc_612 N_A_27_84#_M1030_d N_A_483_74#_c_1108_n 0.00178571f $X=3.71 $Y=0.37 $X2=0
+ $Y2=0
cc_613 N_A_27_84#_M1015_s N_A_483_74#_c_1108_n 0.00170263f $X=4.57 $Y=0.37 $X2=0
+ $Y2=0
cc_614 N_A_27_84#_M1028_s N_A_483_74#_c_1108_n 0.00179007f $X=5.43 $Y=0.37 $X2=0
+ $Y2=0
cc_615 N_A_27_84#_c_1034_n N_A_483_74#_c_1108_n 0.00427478f $X=3.685 $Y=1.095
+ $X2=0 $Y2=0
cc_616 N_A_27_84#_c_1037_n N_A_483_74#_c_1108_n 0.0162997f $X=3.85 $Y=0.89 $X2=0
+ $Y2=0
cc_617 N_A_27_84#_c_1067_n N_A_483_74#_c_1108_n 0.0907973f $X=5.405 $Y=0.91
+ $X2=0 $Y2=0
cc_618 N_A_27_84#_c_1028_n N_VGND_c_1221_n 0.043102f $X=1.045 $Y=0.34 $X2=0
+ $Y2=0
cc_619 N_A_27_84#_c_1029_n N_VGND_c_1221_n 0.0186386f $X=0.375 $Y=0.34 $X2=0
+ $Y2=0
cc_620 N_A_27_84#_c_1030_n N_VGND_c_1221_n 0.0616678f $X=1.915 $Y=0.34 $X2=0
+ $Y2=0
cc_621 N_A_27_84#_c_1035_n N_VGND_c_1221_n 0.0134682f $X=1.14 $Y=0.34 $X2=0
+ $Y2=0
cc_622 N_A_27_84#_c_1028_n N_VGND_c_1226_n 0.0251825f $X=1.045 $Y=0.34 $X2=0
+ $Y2=0
cc_623 N_A_27_84#_c_1029_n N_VGND_c_1226_n 0.0101082f $X=0.375 $Y=0.34 $X2=0
+ $Y2=0
cc_624 N_A_27_84#_c_1030_n N_VGND_c_1226_n 0.0352779f $X=1.915 $Y=0.34 $X2=0
+ $Y2=0
cc_625 N_A_27_84#_c_1032_n N_VGND_c_1226_n 0.0105008f $X=2.95 $Y=0.975 $X2=0
+ $Y2=0
cc_626 N_A_27_84#_c_1035_n N_VGND_c_1226_n 0.00735812f $X=1.14 $Y=0.34 $X2=0
+ $Y2=0
cc_627 N_A_483_74#_c_1129_n N_VGND_M1005_s 0.00678566f $X=6.905 $Y=0.835
+ $X2=-0.19 $Y2=-0.245
cc_628 N_A_483_74#_c_1134_n N_VGND_M1011_d 0.00472947f $X=7.835 $Y=0.835 $X2=0
+ $Y2=0
cc_629 N_A_483_74#_c_1135_n N_VGND_M1022_d 0.00398331f $X=8.775 $Y=0.835 $X2=0
+ $Y2=0
cc_630 N_A_483_74#_c_1112_n N_VGND_M1031_s 0.00330483f $X=9.715 $Y=1.005 $X2=0
+ $Y2=0
cc_631 N_A_483_74#_c_1129_n N_VGND_c_1217_n 0.0240865f $X=6.905 $Y=0.835 $X2=0
+ $Y2=0
cc_632 N_A_483_74#_c_1109_n N_VGND_c_1217_n 0.00906117f $X=7.07 $Y=0.635 $X2=0
+ $Y2=0
cc_633 N_A_483_74#_c_1114_n N_VGND_c_1217_n 0.00942064f $X=6.07 $Y=0.475 $X2=0
+ $Y2=0
cc_634 N_A_483_74#_c_1109_n N_VGND_c_1218_n 0.00897147f $X=7.07 $Y=0.635 $X2=0
+ $Y2=0
cc_635 N_A_483_74#_c_1134_n N_VGND_c_1218_n 0.0203034f $X=7.835 $Y=0.835 $X2=0
+ $Y2=0
cc_636 N_A_483_74#_c_1110_n N_VGND_c_1218_n 0.00906117f $X=8 $Y=0.635 $X2=0
+ $Y2=0
cc_637 N_A_483_74#_c_1110_n N_VGND_c_1219_n 0.00900923f $X=8 $Y=0.635 $X2=0
+ $Y2=0
cc_638 N_A_483_74#_c_1135_n N_VGND_c_1219_n 0.0173074f $X=8.775 $Y=0.835 $X2=0
+ $Y2=0
cc_639 N_A_483_74#_c_1111_n N_VGND_c_1219_n 0.00942763f $X=8.94 $Y=0.515 $X2=0
+ $Y2=0
cc_640 N_A_483_74#_c_1111_n N_VGND_c_1220_n 0.0150645f $X=8.94 $Y=0.515 $X2=0
+ $Y2=0
cc_641 N_A_483_74#_c_1112_n N_VGND_c_1220_n 0.0171619f $X=9.715 $Y=1.005 $X2=0
+ $Y2=0
cc_642 N_A_483_74#_c_1113_n N_VGND_c_1220_n 0.0150645f $X=9.8 $Y=0.515 $X2=0
+ $Y2=0
cc_643 N_A_483_74#_c_1107_n N_VGND_c_1221_n 0.0454606f $X=3.335 $Y=0.475 $X2=0
+ $Y2=0
cc_644 N_A_483_74#_c_1108_n N_VGND_c_1221_n 0.0970299f $X=5.905 $Y=0.475 $X2=0
+ $Y2=0
cc_645 N_A_483_74#_c_1129_n N_VGND_c_1221_n 0.00190416f $X=6.905 $Y=0.835 $X2=0
+ $Y2=0
cc_646 N_A_483_74#_c_1114_n N_VGND_c_1221_n 0.0145639f $X=6.07 $Y=0.475 $X2=0
+ $Y2=0
cc_647 N_A_483_74#_c_1129_n N_VGND_c_1222_n 0.00189877f $X=6.905 $Y=0.835 $X2=0
+ $Y2=0
cc_648 N_A_483_74#_c_1109_n N_VGND_c_1222_n 0.0108551f $X=7.07 $Y=0.635 $X2=0
+ $Y2=0
cc_649 N_A_483_74#_c_1134_n N_VGND_c_1222_n 0.00197156f $X=7.835 $Y=0.835 $X2=0
+ $Y2=0
cc_650 N_A_483_74#_c_1134_n N_VGND_c_1223_n 0.00189877f $X=7.835 $Y=0.835 $X2=0
+ $Y2=0
cc_651 N_A_483_74#_c_1110_n N_VGND_c_1223_n 0.0108551f $X=8 $Y=0.635 $X2=0 $Y2=0
cc_652 N_A_483_74#_c_1135_n N_VGND_c_1223_n 0.00197156f $X=8.775 $Y=0.835 $X2=0
+ $Y2=0
cc_653 N_A_483_74#_c_1135_n N_VGND_c_1224_n 0.00190416f $X=8.775 $Y=0.835 $X2=0
+ $Y2=0
cc_654 N_A_483_74#_c_1111_n N_VGND_c_1224_n 0.011066f $X=8.94 $Y=0.515 $X2=0
+ $Y2=0
cc_655 N_A_483_74#_c_1113_n N_VGND_c_1225_n 0.011066f $X=9.8 $Y=0.515 $X2=0
+ $Y2=0
cc_656 N_A_483_74#_c_1107_n N_VGND_c_1226_n 0.0383078f $X=3.335 $Y=0.475 $X2=0
+ $Y2=0
cc_657 N_A_483_74#_c_1108_n N_VGND_c_1226_n 0.0814955f $X=5.905 $Y=0.475 $X2=0
+ $Y2=0
cc_658 N_A_483_74#_c_1129_n N_VGND_c_1226_n 0.00891641f $X=6.905 $Y=0.835 $X2=0
+ $Y2=0
cc_659 N_A_483_74#_c_1109_n N_VGND_c_1226_n 0.00898945f $X=7.07 $Y=0.635 $X2=0
+ $Y2=0
cc_660 N_A_483_74#_c_1134_n N_VGND_c_1226_n 0.00914714f $X=7.835 $Y=0.835 $X2=0
+ $Y2=0
cc_661 N_A_483_74#_c_1110_n N_VGND_c_1226_n 0.00898945f $X=8 $Y=0.635 $X2=0
+ $Y2=0
cc_662 N_A_483_74#_c_1135_n N_VGND_c_1226_n 0.00917295f $X=8.775 $Y=0.835 $X2=0
+ $Y2=0
cc_663 N_A_483_74#_c_1111_n N_VGND_c_1226_n 0.00915947f $X=8.94 $Y=0.515 $X2=0
+ $Y2=0
cc_664 N_A_483_74#_c_1113_n N_VGND_c_1226_n 0.00915947f $X=9.8 $Y=0.515 $X2=0
+ $Y2=0
cc_665 N_A_483_74#_c_1114_n N_VGND_c_1226_n 0.0119984f $X=6.07 $Y=0.475 $X2=0
+ $Y2=0
