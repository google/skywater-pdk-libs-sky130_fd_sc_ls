* File: sky130_fd_sc_ls__a32o_1.pxi.spice
* Created: Wed Sep  2 10:52:47 2020
* 
x_PM_SKY130_FD_SC_LS__A32O_1%A_84_48# N_A_84_48#_M1011_d N_A_84_48#_M1010_d
+ N_A_84_48#_M1009_g N_A_84_48#_c_55_n N_A_84_48#_M1003_g N_A_84_48#_c_56_n
+ N_A_84_48#_c_122_p N_A_84_48#_c_60_n N_A_84_48#_c_118_p N_A_84_48#_c_57_n
+ N_A_84_48#_c_58_n N_A_84_48#_c_67_p PM_SKY130_FD_SC_LS__A32O_1%A_84_48#
x_PM_SKY130_FD_SC_LS__A32O_1%A3 N_A3_c_137_n N_A3_M1001_g N_A3_c_138_n
+ N_A3_M1005_g A3 PM_SKY130_FD_SC_LS__A32O_1%A3
x_PM_SKY130_FD_SC_LS__A32O_1%A2 N_A2_c_168_n N_A2_M1002_g N_A2_c_169_n
+ N_A2_M1006_g A2 PM_SKY130_FD_SC_LS__A32O_1%A2
x_PM_SKY130_FD_SC_LS__A32O_1%A1 N_A1_c_195_n N_A1_M1011_g N_A1_c_196_n
+ N_A1_M1007_g A1 PM_SKY130_FD_SC_LS__A32O_1%A1
x_PM_SKY130_FD_SC_LS__A32O_1%B1 N_B1_c_224_n N_B1_M1010_g N_B1_c_225_n
+ N_B1_M1004_g B1 N_B1_c_226_n PM_SKY130_FD_SC_LS__A32O_1%B1
x_PM_SKY130_FD_SC_LS__A32O_1%B2 N_B2_c_252_n N_B2_M1008_g N_B2_c_253_n
+ N_B2_M1000_g B2 PM_SKY130_FD_SC_LS__A32O_1%B2
x_PM_SKY130_FD_SC_LS__A32O_1%X N_X_M1009_s N_X_M1003_s N_X_c_276_n N_X_c_277_n
+ N_X_c_273_n X X X PM_SKY130_FD_SC_LS__A32O_1%X
x_PM_SKY130_FD_SC_LS__A32O_1%VPWR N_VPWR_M1003_d N_VPWR_M1002_d N_VPWR_c_298_n
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n VPWR N_VPWR_c_302_n
+ N_VPWR_c_303_n N_VPWR_c_297_n N_VPWR_c_305_n PM_SKY130_FD_SC_LS__A32O_1%VPWR
x_PM_SKY130_FD_SC_LS__A32O_1%A_244_368# N_A_244_368#_M1001_d
+ N_A_244_368#_M1007_d N_A_244_368#_M1000_d N_A_244_368#_c_346_n
+ N_A_244_368#_c_347_n N_A_244_368#_c_356_n N_A_244_368#_c_340_n
+ N_A_244_368#_c_341_n N_A_244_368#_c_342_n N_A_244_368#_c_343_n
+ PM_SKY130_FD_SC_LS__A32O_1%A_244_368#
x_PM_SKY130_FD_SC_LS__A32O_1%VGND N_VGND_M1009_d N_VGND_M1008_d N_VGND_c_379_n
+ N_VGND_c_380_n N_VGND_c_381_n VGND N_VGND_c_382_n N_VGND_c_383_n
+ N_VGND_c_384_n PM_SKY130_FD_SC_LS__A32O_1%VGND
cc_1 VNB N_A_84_48#_M1009_g 0.029153f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_84_48#_c_55_n 0.0350036f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.765
cc_3 VNB N_A_84_48#_c_56_n 0.00309123f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.3
cc_4 VNB N_A_84_48#_c_57_n 0.00575673f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_5 VNB N_A_84_48#_c_58_n 0.00655964f $X=-0.19 $Y=-0.245 $X2=2.715 $Y2=0.595
cc_6 VNB N_A3_c_137_n 0.0367912f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.47
cc_7 VNB N_A3_c_138_n 0.0183757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB A3 0.0058955f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_9 VNB N_A2_c_168_n 0.0391488f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.47
cc_10 VNB N_A2_c_169_n 0.0173277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB A2 0.00343145f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_12 VNB N_A1_c_195_n 0.0199178f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.47
cc_13 VNB N_A1_c_196_n 0.044209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A1 0.00392553f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_15 VNB N_B1_c_224_n 0.0350175f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.47
cc_16 VNB N_B1_c_225_n 0.018627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_c_226_n 0.00901079f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.765
cc_18 VNB N_B2_c_252_n 0.020822f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.47
cc_19 VNB N_B2_c_253_n 0.0497475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB B2 0.0174691f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_21 VNB N_X_c_273_n 0.0247148f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.3
cc_22 VNB X 0.0265914f $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=0.935
cc_23 VNB X 0.0139041f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=0.935
cc_24 VNB N_VPWR_c_297_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_379_n 0.0134045f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.765
cc_26 VNB N_VGND_c_380_n 0.0130142f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_27 VNB N_VGND_c_381_n 0.0401609f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.3
cc_28 VNB N_VGND_c_382_n 0.0692324f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.805
cc_29 VNB N_VGND_c_383_n 0.0277248f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_30 VNB N_VGND_c_384_n 0.251223f $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=0.725
cc_31 VPB N_A_84_48#_c_55_n 0.0296995f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.765
cc_32 VPB N_A_84_48#_c_60_n 0.040771f $X=-0.19 $Y=1.66 $X2=2.895 $Y2=1.805
cc_33 VPB N_A_84_48#_c_57_n 0.0022822f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.465
cc_34 VPB N_A3_c_137_n 0.0225014f $X=-0.19 $Y=1.66 $X2=2.225 $Y2=0.47
cc_35 VPB N_A2_c_168_n 0.0233717f $X=-0.19 $Y=1.66 $X2=2.225 $Y2=0.47
cc_36 VPB N_A1_c_196_n 0.0227366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_B1_c_224_n 0.0209454f $X=-0.19 $Y=1.66 $X2=2.225 $Y2=0.47
cc_38 VPB N_B2_c_253_n 0.0291458f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_X_c_276_n 0.0420589f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.765
cc_40 VPB N_X_c_277_n 0.0143501f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.02
cc_41 VPB N_X_c_273_n 0.00757678f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.3
cc_42 VPB N_VPWR_c_298_n 0.0152241f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_43 VPB N_VPWR_c_299_n 0.0169573f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.3
cc_44 VPB N_VPWR_c_300_n 0.0228926f $X=-0.19 $Y=1.66 $X2=2.895 $Y2=1.805
cc_45 VPB N_VPWR_c_301_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=1.805
cc_46 VPB N_VPWR_c_302_n 0.0191572f $X=-0.19 $Y=1.66 $X2=3.06 $Y2=1.97
cc_47 VPB N_VPWR_c_303_n 0.044059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_297_n 0.0829063f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_305_n 0.00747566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_244_368#_c_340_n 0.0206603f $X=-0.19 $Y=1.66 $X2=2.2 $Y2=0.935
cc_51 VPB N_A_244_368#_c_341_n 0.00356803f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=0.935
cc_52 VPB N_A_244_368#_c_342_n 0.0445225f $X=-0.19 $Y=1.66 $X2=3.06 $Y2=1.89
cc_53 VPB N_A_244_368#_c_343_n 0.003137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 N_A_84_48#_M1009_g N_A3_c_137_n 0.00180795f $X=0.495 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_55 N_A_84_48#_c_55_n N_A3_c_137_n 0.0418995f $X=0.515 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_56 N_A_84_48#_c_56_n N_A3_c_137_n 6.05416e-19 $X=0.71 $Y=1.3 $X2=-0.19
+ $Y2=-0.245
cc_57 N_A_84_48#_c_60_n N_A3_c_137_n 0.0173499f $X=2.895 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_58 N_A_84_48#_c_57_n N_A3_c_137_n 0.0050083f $X=0.59 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_59 N_A_84_48#_c_67_p N_A3_c_137_n 0.00103446f $X=2.2 $Y=0.725 $X2=-0.19
+ $Y2=-0.245
cc_60 N_A_84_48#_M1009_g N_A3_c_138_n 0.0131011f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_61 N_A_84_48#_c_56_n N_A3_c_138_n 0.00325245f $X=0.71 $Y=1.3 $X2=0 $Y2=0
cc_62 N_A_84_48#_c_67_p N_A3_c_138_n 0.0126218f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_63 N_A_84_48#_c_55_n A3 2.8743e-19 $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_64 N_A_84_48#_c_56_n A3 0.00839161f $X=0.71 $Y=1.3 $X2=0 $Y2=0
cc_65 N_A_84_48#_c_60_n A3 0.0258645f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_66 N_A_84_48#_c_57_n A3 0.0201492f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_67 N_A_84_48#_c_67_p A3 0.0236883f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_68 N_A_84_48#_c_60_n N_A2_c_168_n 0.0137321f $X=2.895 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_69 N_A_84_48#_c_67_p N_A2_c_168_n 8.47471e-19 $X=2.2 $Y=0.725 $X2=-0.19
+ $Y2=-0.245
cc_70 N_A_84_48#_c_58_n N_A2_c_169_n 0.00192815f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_71 N_A_84_48#_c_67_p N_A2_c_169_n 0.0120996f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_72 N_A_84_48#_c_60_n A2 0.0242683f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_73 N_A_84_48#_c_67_p A2 0.0217461f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_74 N_A_84_48#_c_58_n N_A1_c_195_n 0.0107943f $X=2.715 $Y=0.595 $X2=-0.19
+ $Y2=-0.245
cc_75 N_A_84_48#_c_67_p N_A1_c_195_n 0.00902659f $X=2.2 $Y=0.725 $X2=-0.19
+ $Y2=-0.245
cc_76 N_A_84_48#_c_60_n N_A1_c_196_n 0.0155185f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_77 N_A_84_48#_c_58_n N_A1_c_196_n 0.00321057f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_78 N_A_84_48#_c_60_n A1 0.0244553f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_79 N_A_84_48#_c_67_p A1 0.0225348f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_80 N_A_84_48#_c_60_n N_B1_c_224_n 0.0198944f $X=2.895 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_81 N_A_84_48#_c_58_n N_B1_c_224_n 0.00112046f $X=2.715 $Y=0.595 $X2=-0.19
+ $Y2=-0.245
cc_82 N_A_84_48#_c_58_n N_B1_c_225_n 0.0111626f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_83 N_A_84_48#_c_60_n N_B1_c_226_n 0.0356446f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_84 N_A_84_48#_c_58_n N_B1_c_226_n 0.0260766f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_85 N_A_84_48#_c_58_n N_B2_c_252_n 0.0016581f $X=2.715 $Y=0.595 $X2=-0.19
+ $Y2=-0.245
cc_86 N_A_84_48#_c_60_n N_B2_c_253_n 0.00391145f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_87 N_A_84_48#_c_55_n N_X_c_276_n 0.0116317f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A_84_48#_c_55_n N_X_c_277_n 0.00438546f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A_84_48#_c_57_n N_X_c_277_n 0.00576634f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_90 N_A_84_48#_M1009_g N_X_c_273_n 0.0100159f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_91 N_A_84_48#_c_55_n N_X_c_273_n 0.0030582f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A_84_48#_c_56_n N_X_c_273_n 0.00523589f $X=0.71 $Y=1.3 $X2=0 $Y2=0
cc_93 N_A_84_48#_c_57_n N_X_c_273_n 0.0315479f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_94 N_A_84_48#_M1009_g X 0.0142066f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A_84_48#_M1009_g X 0.0028169f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_96 N_A_84_48#_c_56_n X 0.00468197f $X=0.71 $Y=1.3 $X2=0 $Y2=0
cc_97 N_A_84_48#_c_57_n X 0.00152458f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_98 N_A_84_48#_c_60_n N_VPWR_M1003_d 0.00252101f $X=2.895 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_99 N_A_84_48#_c_57_n N_VPWR_M1003_d 0.0020474f $X=0.59 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_100 N_A_84_48#_c_60_n N_VPWR_M1002_d 0.00561474f $X=2.895 $Y=1.805 $X2=0
+ $Y2=0
cc_101 N_A_84_48#_c_55_n N_VPWR_c_298_n 0.0118734f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_84_48#_c_60_n N_VPWR_c_298_n 0.0176997f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_103 N_A_84_48#_c_57_n N_VPWR_c_298_n 0.0133439f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_104 N_A_84_48#_c_55_n N_VPWR_c_302_n 0.00445602f $X=0.515 $Y=1.765 $X2=0
+ $Y2=0
cc_105 N_A_84_48#_c_55_n N_VPWR_c_297_n 0.00865246f $X=0.515 $Y=1.765 $X2=0
+ $Y2=0
cc_106 N_A_84_48#_c_60_n N_A_244_368#_M1001_d 0.00197722f $X=2.895 $Y=1.805
+ $X2=-0.19 $Y2=-0.245
cc_107 N_A_84_48#_c_60_n N_A_244_368#_M1007_d 0.00197722f $X=2.895 $Y=1.805
+ $X2=0 $Y2=0
cc_108 N_A_84_48#_c_60_n N_A_244_368#_c_346_n 0.0528064f $X=2.895 $Y=1.805 $X2=0
+ $Y2=0
cc_109 N_A_84_48#_c_60_n N_A_244_368#_c_347_n 0.0173337f $X=2.895 $Y=1.805 $X2=0
+ $Y2=0
cc_110 N_A_84_48#_c_118_p N_A_244_368#_c_340_n 0.0237369f $X=3.06 $Y=1.97 $X2=0
+ $Y2=0
cc_111 N_A_84_48#_c_60_n N_A_244_368#_c_342_n 0.0035248f $X=2.895 $Y=1.805 $X2=0
+ $Y2=0
cc_112 N_A_84_48#_c_60_n N_A_244_368#_c_343_n 0.0173337f $X=2.895 $Y=1.805 $X2=0
+ $Y2=0
cc_113 N_A_84_48#_c_56_n N_VGND_M1009_d 0.00198882f $X=0.71 $Y=1.3 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A_84_48#_c_122_p N_VGND_M1009_d 0.00372868f $X=0.795 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_115 N_A_84_48#_c_67_p N_VGND_M1009_d 0.0125332f $X=2.2 $Y=0.725 $X2=-0.19
+ $Y2=-0.245
cc_116 N_A_84_48#_M1009_g N_VGND_c_379_n 0.00811597f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_117 N_A_84_48#_c_55_n N_VGND_c_379_n 3.34594e-19 $X=0.515 $Y=1.765 $X2=0
+ $Y2=0
cc_118 N_A_84_48#_c_122_p N_VGND_c_379_n 0.0126823f $X=0.795 $Y=0.935 $X2=0
+ $Y2=0
cc_119 N_A_84_48#_c_67_p N_VGND_c_379_n 0.0201945f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_120 N_A_84_48#_c_58_n N_VGND_c_381_n 0.0197562f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_121 N_A_84_48#_c_58_n N_VGND_c_382_n 0.0224837f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_122 N_A_84_48#_M1009_g N_VGND_c_383_n 0.00434272f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_123 N_A_84_48#_M1009_g N_VGND_c_384_n 0.00829501f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_124 N_A_84_48#_c_122_p N_VGND_c_384_n 0.00149237f $X=0.795 $Y=0.935 $X2=0
+ $Y2=0
cc_125 N_A_84_48#_c_58_n N_VGND_c_384_n 0.0236713f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_126 N_A_84_48#_c_67_p N_VGND_c_384_n 0.0387864f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_127 N_A_84_48#_c_67_p A_259_94# 0.00736231f $X=2.2 $Y=0.725 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_84_48#_c_67_p A_337_94# 0.013672f $X=2.2 $Y=0.725 $X2=-0.19
+ $Y2=-0.245
cc_129 N_A3_c_137_n N_A2_c_168_n 0.0519528f $X=1.145 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_130 A3 N_A2_c_168_n 0.00188716f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_131 N_A3_c_138_n N_A2_c_169_n 0.049285f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_132 N_A3_c_137_n A2 3.99347e-19 $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_133 A3 A2 0.0264591f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_134 N_A3_c_137_n N_X_c_277_n 9.34777e-19 $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A3_c_137_n N_VPWR_c_298_n 0.00872653f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A3_c_137_n N_VPWR_c_300_n 0.00481995f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A3_c_137_n N_VPWR_c_297_n 0.00508379f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A3_c_137_n N_A_244_368#_c_343_n 0.0103165f $X=1.145 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A3_c_138_n N_VGND_c_379_n 0.010194f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_140 N_A3_c_138_n N_VGND_c_382_n 0.00507111f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_141 N_A3_c_138_n N_VGND_c_384_n 0.00514438f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_142 N_A2_c_169_n N_A1_c_195_n 0.0291659f $X=1.61 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_143 N_A2_c_168_n N_A1_c_196_n 0.0449869f $X=1.595 $Y=1.765 $X2=0 $Y2=0
cc_144 A2 N_A1_c_196_n 0.00118009f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_145 N_A2_c_168_n A1 0.00114936f $X=1.595 $Y=1.765 $X2=0 $Y2=0
cc_146 A2 A1 0.0230669f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_147 N_A2_c_168_n N_VPWR_c_299_n 0.00807742f $X=1.595 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A2_c_168_n N_VPWR_c_300_n 0.00481995f $X=1.595 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A2_c_168_n N_VPWR_c_297_n 0.00508379f $X=1.595 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A2_c_168_n N_A_244_368#_c_346_n 0.0130998f $X=1.595 $Y=1.765 $X2=0
+ $Y2=0
cc_151 N_A2_c_168_n N_A_244_368#_c_343_n 0.0153066f $X=1.595 $Y=1.765 $X2=0
+ $Y2=0
cc_152 N_A2_c_169_n N_VGND_c_382_n 0.00507111f $X=1.61 $Y=1.22 $X2=0 $Y2=0
cc_153 N_A2_c_169_n N_VGND_c_384_n 0.00514438f $X=1.61 $Y=1.22 $X2=0 $Y2=0
cc_154 N_A1_c_196_n N_B1_c_224_n 0.0475663f $X=2.335 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_155 A1 N_B1_c_224_n 3.04283e-19 $X=2.075 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_156 N_A1_c_195_n N_B1_c_225_n 0.00495039f $X=2.15 $Y=1.22 $X2=0 $Y2=0
cc_157 N_A1_c_196_n N_B1_c_226_n 0.002359f $X=2.335 $Y=1.765 $X2=0 $Y2=0
cc_158 A1 N_B1_c_226_n 0.0293561f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_159 N_A1_c_196_n N_VPWR_c_299_n 0.00621168f $X=2.335 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A1_c_196_n N_VPWR_c_303_n 0.00451897f $X=2.335 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A1_c_196_n N_VPWR_c_297_n 0.00457541f $X=2.335 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A1_c_196_n N_A_244_368#_c_346_n 0.0130998f $X=2.335 $Y=1.765 $X2=0
+ $Y2=0
cc_163 N_A1_c_196_n N_A_244_368#_c_347_n 4.27055e-19 $X=2.335 $Y=1.765 $X2=0
+ $Y2=0
cc_164 N_A1_c_196_n N_A_244_368#_c_356_n 0.0157962f $X=2.335 $Y=1.765 $X2=0
+ $Y2=0
cc_165 N_A1_c_196_n N_A_244_368#_c_341_n 0.00186581f $X=2.335 $Y=1.765 $X2=0
+ $Y2=0
cc_166 N_A1_c_195_n N_VGND_c_382_n 0.00484285f $X=2.15 $Y=1.22 $X2=0 $Y2=0
cc_167 N_A1_c_195_n N_VGND_c_384_n 0.00514438f $X=2.15 $Y=1.22 $X2=0 $Y2=0
cc_168 N_B1_c_225_n N_B2_c_252_n 0.031246f $X=2.93 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_169 N_B1_c_226_n N_B2_c_252_n 0.00143086f $X=2.84 $Y=1.385 $X2=-0.19
+ $Y2=-0.245
cc_170 N_B1_c_224_n N_B2_c_253_n 0.0659776f $X=2.785 $Y=1.765 $X2=0 $Y2=0
cc_171 N_B1_c_225_n B2 4.01112e-19 $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_172 N_B1_c_226_n B2 0.017611f $X=2.84 $Y=1.385 $X2=0 $Y2=0
cc_173 N_B1_c_224_n N_VPWR_c_303_n 7.44201e-19 $X=2.785 $Y=1.765 $X2=0 $Y2=0
cc_174 N_B1_c_224_n N_A_244_368#_c_347_n 0.00184286f $X=2.785 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_B1_c_224_n N_A_244_368#_c_356_n 0.010488f $X=2.785 $Y=1.765 $X2=0 $Y2=0
cc_176 N_B1_c_224_n N_A_244_368#_c_340_n 0.00990262f $X=2.785 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_B1_c_224_n N_A_244_368#_c_341_n 0.00114023f $X=2.785 $Y=1.765 $X2=0
+ $Y2=0
cc_178 N_B1_c_224_n N_A_244_368#_c_342_n 7.42913e-19 $X=2.785 $Y=1.765 $X2=0
+ $Y2=0
cc_179 N_B1_c_225_n N_VGND_c_381_n 0.0022187f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_180 N_B1_c_225_n N_VGND_c_382_n 0.00484285f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_181 N_B1_c_225_n N_VGND_c_384_n 0.00514438f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_182 N_B2_c_253_n N_VPWR_c_303_n 7.44201e-19 $X=3.335 $Y=1.765 $X2=0 $Y2=0
cc_183 N_B2_c_253_n N_A_244_368#_c_356_n 6.25647e-19 $X=3.335 $Y=1.765 $X2=0
+ $Y2=0
cc_184 N_B2_c_253_n N_A_244_368#_c_340_n 0.0115629f $X=3.335 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_B2_c_253_n N_A_244_368#_c_342_n 0.01879f $X=3.335 $Y=1.765 $X2=0 $Y2=0
cc_186 B2 N_A_244_368#_c_342_n 0.0194401f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_187 N_B2_c_252_n N_VGND_c_381_n 0.0151934f $X=3.32 $Y=1.22 $X2=0 $Y2=0
cc_188 N_B2_c_253_n N_VGND_c_381_n 0.0015621f $X=3.335 $Y=1.765 $X2=0 $Y2=0
cc_189 B2 N_VGND_c_381_n 0.0257644f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_190 N_B2_c_252_n N_VGND_c_382_n 0.00421418f $X=3.32 $Y=1.22 $X2=0 $Y2=0
cc_191 N_B2_c_252_n N_VGND_c_384_n 0.00432128f $X=3.32 $Y=1.22 $X2=0 $Y2=0
cc_192 N_X_c_276_n N_VPWR_c_298_n 0.0359411f $X=0.29 $Y=2.815 $X2=0 $Y2=0
cc_193 N_X_c_276_n N_VPWR_c_302_n 0.0163786f $X=0.29 $Y=2.815 $X2=0 $Y2=0
cc_194 N_X_c_276_n N_VPWR_c_297_n 0.0135239f $X=0.29 $Y=2.815 $X2=0 $Y2=0
cc_195 X N_VGND_c_379_n 0.0226903f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_196 X N_VGND_c_383_n 0.0159025f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_197 X N_VGND_c_384_n 0.0131064f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_198 N_VPWR_M1002_d N_A_244_368#_c_346_n 0.0160396f $X=1.67 $Y=1.84 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_299_n N_A_244_368#_c_346_n 0.0266856f $X=1.965 $Y=2.565 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_299_n N_A_244_368#_c_356_n 0.0279707f $X=1.965 $Y=2.565 $X2=0
+ $Y2=0
cc_201 N_VPWR_c_303_n N_A_244_368#_c_340_n 0.0667586f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_202 N_VPWR_c_297_n N_A_244_368#_c_340_n 0.0380121f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_203 N_VPWR_c_299_n N_A_244_368#_c_341_n 0.0107171f $X=1.965 $Y=2.565 $X2=0
+ $Y2=0
cc_204 N_VPWR_c_303_n N_A_244_368#_c_341_n 0.0236566f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_205 N_VPWR_c_297_n N_A_244_368#_c_341_n 0.0128296f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_206 N_VPWR_c_298_n N_A_244_368#_c_343_n 0.0223391f $X=0.85 $Y=2.225 $X2=0
+ $Y2=0
cc_207 N_VPWR_c_299_n N_A_244_368#_c_343_n 0.025439f $X=1.965 $Y=2.565 $X2=0
+ $Y2=0
cc_208 N_VPWR_c_300_n N_A_244_368#_c_343_n 0.00976219f $X=1.8 $Y=3.33 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_297_n N_A_244_368#_c_343_n 0.0111764f $X=3.6 $Y=3.33 $X2=0 $Y2=0
