# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ls__ha_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__ha_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.468000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.450000 0.255000 2.780000 0.670000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.468000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.765000 1.470000 2.095000 1.550000 ;
        RECT 1.765000 1.550000 3.300000 1.800000 ;
        RECT 2.970000 1.470000 3.300000 1.550000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.310000 0.475000 4.715000 1.180000 ;
        RECT 4.310000 1.850000 4.715000 2.980000 ;
        RECT 4.545000 1.180000 4.715000 1.850000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.350000 0.445000 1.130000 ;
        RECT 0.115000 1.130000 0.355000 1.820000 ;
        RECT 0.115000 1.820000 0.445000 2.980000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 4.800000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 1.745000 1.780000 ;
        RECT -0.190000 1.780000 4.990000 3.520000 ;
        RECT  3.110000 1.660000 4.990000 1.780000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.525000  1.300000 0.855000 1.630000 ;
      RECT 0.615000  2.650000 1.205000 3.245000 ;
      RECT 0.625000  0.085000 0.875000 0.795000 ;
      RECT 0.685000  1.130000 1.400000 1.300000 ;
      RECT 0.685000  1.630000 0.855000 2.310000 ;
      RECT 0.685000  2.310000 1.740000 2.480000 ;
      RECT 1.070000  0.910000 1.400000 1.130000 ;
      RECT 1.195000  1.470000 1.525000 1.970000 ;
      RECT 1.195000  1.970000 3.640000 2.140000 ;
      RECT 1.410000  2.480000 1.740000 2.800000 ;
      RECT 1.580000  0.630000 1.750000 1.130000 ;
      RECT 1.580000  1.130000 2.790000 1.300000 ;
      RECT 1.930000  0.085000 2.280000 0.960000 ;
      RECT 2.460000  0.840000 2.790000 1.130000 ;
      RECT 2.460000  1.300000 2.790000 1.355000 ;
      RECT 2.485000  2.310000 3.190000 3.245000 ;
      RECT 3.020000  0.575000 3.350000 1.085000 ;
      RECT 3.020000  1.085000 3.640000 1.255000 ;
      RECT 3.360000  2.140000 3.640000 2.980000 ;
      RECT 3.470000  1.255000 3.640000 1.350000 ;
      RECT 3.470000  1.350000 4.375000 1.680000 ;
      RECT 3.470000  1.680000 3.640000 1.970000 ;
      RECT 3.810000  0.085000 4.140000 1.180000 ;
      RECT 3.810000  2.100000 4.140000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_ls__ha_1
END LIBRARY
