* File: sky130_fd_sc_ls__dfxtp_2.pex.spice
* Created: Wed Sep  2 11:02:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DFXTP_2%CLK 3 5 7 8 12
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.34
+ $Y=1.465 $X2=0.34 $Y2=1.465
r33 8 12 6.06549 $w=3.78e-07 $l=2e-07 $layer=LI1_cond $X=0.315 $Y=1.665
+ $X2=0.315 $Y2=1.465
r34 5 11 57.3754 $w=3.5e-07 $l=3.54965e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.385 $Y2=1.465
r35 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r36 1 11 38.7839 $w=3.5e-07 $l=2.13014e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.385 $Y2=1.465
r37 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__DFXTP_2%A_27_74# 1 2 7 9 10 12 15 18 19 21 22 24 25
+ 30 34 36 38 40 41 42 45 48 49 51 52 53 55 56 57 59 61 63 64 67 69 72 73 86 90
+ 91 92 96
c262 96 0 6.76432e-20 $X=3.145 $Y=1.92
c263 90 0 6.36416e-20 $X=5.725 $Y=0.345
c264 88 0 2.82287e-20 $X=3.67 $Y=0.775
c265 61 0 1.41143e-20 $X=3.67 $Y=0.69
c266 15 0 5.64678e-20 $X=2.99 $Y=0.805
c267 7 0 8.02678e-20 $X=0.955 $Y=1.765
r268 91 100 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.725 $Y=0.345
+ $X2=5.725 $Y2=0.51
r269 90 92 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=0.382
+ $X2=5.56 $Y2=0.382
r270 90 91 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.725
+ $Y=0.345 $X2=5.725 $Y2=0.345
r271 84 86 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.455 $Y=1.37
+ $X2=3.67 $Y2=1.37
r272 80 96 27.1549 $w=2.84e-07 $l=1.6e-07 $layer=POLY_cond $X=3.305 $Y=1.92
+ $X2=3.145 $Y2=1.92
r273 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.305
+ $Y=1.92 $X2=3.305 $Y2=1.92
r274 75 77 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=1.385
+ $X2=0.905 $Y2=1.55
r275 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.385 $X2=0.97 $Y2=1.385
r276 72 75 8.84058 $w=4.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.905 $Y=1.045
+ $X2=0.905 $Y2=1.385
r277 72 73 7.19996 $w=4.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.905 $Y=1.045
+ $X2=0.905 $Y2=0.96
r278 69 92 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=4.575 $Y=0.34
+ $X2=5.56 $Y2=0.34
r279 66 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.49 $Y=0.425
+ $X2=4.575 $Y2=0.34
r280 66 67 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.49 $Y=0.425
+ $X2=4.49 $Y2=0.69
r281 65 88 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.755 $Y=0.775
+ $X2=3.67 $Y2=0.775
r282 64 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.405 $Y=0.775
+ $X2=4.49 $Y2=0.69
r283 64 65 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.405 $Y=0.775
+ $X2=3.755 $Y2=0.775
r284 63 86 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=1.285
+ $X2=3.67 $Y2=1.37
r285 62 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=0.86
+ $X2=3.67 $Y2=0.775
r286 62 63 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.67 $Y=0.86
+ $X2=3.67 $Y2=1.285
r287 61 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=0.69
+ $X2=3.67 $Y2=0.775
r288 60 61 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.67 $Y=0.425
+ $X2=3.67 $Y2=0.69
r289 59 79 6.77908 $w=2.53e-07 $l=1.5e-07 $layer=LI1_cond $X=3.455 $Y=1.957
+ $X2=3.305 $Y2=1.957
r290 58 84 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=1.455
+ $X2=3.455 $Y2=1.37
r291 58 59 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.455 $Y=1.455
+ $X2=3.455 $Y2=1.83
r292 56 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.585 $Y=0.34
+ $X2=3.67 $Y2=0.425
r293 56 57 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=3.585 $Y=0.34
+ $X2=2.52 $Y2=0.34
r294 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.435 $Y=0.425
+ $X2=2.52 $Y2=0.34
r295 54 55 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.435 $Y=0.425
+ $X2=2.435 $Y2=0.81
r296 52 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.35 $Y=0.895
+ $X2=2.435 $Y2=0.81
r297 52 53 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.35 $Y=0.895
+ $X2=1.815 $Y2=0.895
r298 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.73 $Y=0.81
+ $X2=1.815 $Y2=0.895
r299 50 51 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.73 $Y=0.425
+ $X2=1.73 $Y2=0.81
r300 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.645 $Y=0.34
+ $X2=1.73 $Y2=0.425
r301 48 49 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.645 $Y=0.34
+ $X2=1.135 $Y2=0.34
r302 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.05 $Y=0.425
+ $X2=1.135 $Y2=0.34
r303 46 73 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=1.05 $Y=0.425
+ $X2=1.05 $Y2=0.96
r304 45 77 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.76 $Y=1.95 $X2=0.76
+ $Y2=1.55
r305 43 71 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r306 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.76 $Y2=1.95
r307 42 43 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.445 $Y2=2.035
r308 40 72 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.675 $Y=1.045
+ $X2=0.905 $Y2=1.045
r309 40 41 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.675 $Y=1.045
+ $X2=0.365 $Y2=1.045
r310 36 71 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.12 $X2=0.28
+ $Y2=2.035
r311 36 38 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=2.815
r312 32 41 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.365 $Y2=1.045
r313 32 34 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.24 $Y2=0.515
r314 30 100 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.785 $Y=0.83
+ $X2=5.785 $Y2=0.51
r315 28 30 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.785 $Y=1.69
+ $X2=5.785 $Y2=0.83
r316 26 31 6.7465 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.11 $Y=1.765 $X2=5.02
+ $Y2=1.765
r317 25 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.71 $Y=1.765
+ $X2=5.785 $Y2=1.69
r318 25 26 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.71 $Y=1.765 $X2=5.11
+ $Y2=1.765
r319 22 31 77.5092 $w=1.77e-07 $l=2.8e-07 $layer=POLY_cond $X=5.02 $Y=2.045
+ $X2=5.02 $Y2=1.765
r320 22 24 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.02 $Y=2.045
+ $X2=5.02 $Y2=2.54
r321 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.145 $Y=2.445
+ $X2=3.145 $Y2=2.73
r322 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.145 $Y=2.355
+ $X2=3.145 $Y2=2.445
r323 17 96 13.4541 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=2.085
+ $X2=3.145 $Y2=1.92
r324 17 18 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=3.145 $Y=2.085
+ $X2=3.145 $Y2=2.355
r325 13 96 26.3063 $w=2.84e-07 $l=2.29783e-07 $layer=POLY_cond $X=2.99 $Y=1.755
+ $X2=3.145 $Y2=1.92
r326 13 15 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.99 $Y=1.755
+ $X2=2.99 $Y2=0.805
r327 10 76 38.666 $w=2.85e-07 $l=2.10286e-07 $layer=POLY_cond $X=1.085 $Y=1.22
+ $X2=0.982 $Y2=1.385
r328 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.085 $Y=1.22
+ $X2=1.085 $Y2=0.74
r329 7 76 75.0274 $w=2.85e-07 $l=3.93268e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.982 $Y2=1.385
r330 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r331 2 71 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r332 2 38 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r333 1 34 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFXTP_2%D 1 3 4 8 13 14 15 17 21
c63 21 0 1.22251e-19 $X=2.165 $Y=1.225
c64 17 0 5.64678e-20 $X=2.16 $Y=1.295
c65 13 0 2.01044e-19 $X=1.89 $Y=2.215
c66 4 0 1.77322e-19 $X=2.485 $Y=1.225
r67 21 24 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.165 $Y=1.225
+ $X2=2.165 $Y2=1.315
r68 17 27 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.16 $Y=1.315
+ $X2=1.97 $Y2=1.315
r69 17 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.165
+ $Y=1.315 $X2=2.165 $Y2=1.315
r70 14 20 25.1593 $w=3.64e-07 $l=1.9e-07 $layer=POLY_cond $X=1.89 $Y=2.257
+ $X2=2.08 $Y2=2.257
r71 13 15 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=2.215
+ $X2=1.89 $Y2=2.05
r72 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.89
+ $Y=2.215 $X2=1.89 $Y2=2.215
r73 10 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.97 $Y=1.48
+ $X2=1.97 $Y2=1.315
r74 10 15 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.97 $Y=1.48
+ $X2=1.97 $Y2=2.05
r75 6 8 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.56 $Y=1.15 $X2=2.56
+ $Y2=0.805
r76 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.33 $Y=1.225
+ $X2=2.165 $Y2=1.225
r77 4 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.485 $Y=1.225
+ $X2=2.56 $Y2=1.15
r78 4 5 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=2.485 $Y=1.225
+ $X2=2.33 $Y2=1.225
r79 1 20 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.08 $Y=2.465
+ $X2=2.08 $Y2=2.257
r80 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.08 $Y=2.465 $X2=2.08
+ $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_LS__DFXTP_2%A_206_368# 1 2 9 10 11 14 15 17 20 24 26 28
+ 30 32 35 37 39 41 43 44 45 49 53 56 59 63 70 71 75
c226 70 0 4.0193e-19 $X=5.25 $Y=1.315
c227 53 0 1.22251e-19 $X=1.39 $Y=1.65
c228 26 0 1.43814e-19 $X=5.55 $Y=2.465
c229 15 0 1.20776e-19 $X=2.615 $Y=2.07
r230 71 72 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.905 $Y=2.71
+ $X2=4.905 $Y2=2.99
r231 70 78 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.25 $Y=1.315
+ $X2=5.125 $Y2=1.315
r232 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.25
+ $Y=1.315 $X2=5.25 $Y2=1.315
r233 63 65 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.455 $Y=2.71
+ $X2=3.455 $Y2=2.84
r234 59 61 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.19 $Y=2.71
+ $X2=2.19 $Y2=2.84
r235 56 76 40.0724 $w=3.6e-07 $l=2.5e-07 $layer=POLY_cond $X=1.58 $Y=1.515
+ $X2=1.58 $Y2=1.765
r236 56 75 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.58 $Y=1.515
+ $X2=1.58 $Y2=1.35
r237 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=1.515 $X2=1.565 $Y2=1.515
r238 53 55 5.81744 $w=3.67e-07 $l=1.75e-07 $layer=LI1_cond $X=1.39 $Y=1.65
+ $X2=1.565 $Y2=1.65
r239 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.71
+ $Y=2.215 $X2=5.71 $Y2=2.215
r240 47 49 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=5.71 $Y=2.905
+ $X2=5.71 $Y2=2.215
r241 46 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=2.99
+ $X2=4.905 $Y2=2.99
r242 45 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.545 $Y=2.99
+ $X2=5.71 $Y2=2.905
r243 45 46 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.545 $Y=2.99
+ $X2=4.99 $Y2=2.99
r244 44 71 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=2.625
+ $X2=4.905 $Y2=2.71
r245 43 69 14.4144 $w=2.92e-07 $l=4.31625e-07 $layer=LI1_cond $X=4.905 $Y=1.54
+ $X2=5.25 $Y2=1.345
r246 43 44 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=4.905 $Y=1.54
+ $X2=4.905 $Y2=2.625
r247 42 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=2.71
+ $X2=3.455 $Y2=2.71
r248 41 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.82 $Y=2.71
+ $X2=4.905 $Y2=2.71
r249 41 42 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=4.82 $Y=2.71
+ $X2=3.54 $Y2=2.71
r250 40 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=2.84
+ $X2=2.19 $Y2=2.84
r251 39 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.37 $Y=2.84
+ $X2=3.455 $Y2=2.84
r252 39 40 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=3.37 $Y=2.84
+ $X2=2.275 $Y2=2.84
r253 38 58 5.73712 $w=1.7e-07 $l=2.7214e-07 $layer=LI1_cond $X=1.475 $Y=2.71
+ $X2=1.245 $Y2=2.802
r254 37 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=2.71
+ $X2=2.19 $Y2=2.71
r255 37 38 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.105 $Y=2.71
+ $X2=1.475 $Y2=2.71
r256 33 53 5.25812 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=1.39 $Y=1.35 $X2=1.39
+ $Y2=1.65
r257 33 35 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.39 $Y=1.35
+ $X2=1.39 $Y2=0.86
r258 30 58 3.15363 $w=4.6e-07 $l=1.77e-07 $layer=LI1_cond $X=1.245 $Y=2.625
+ $X2=1.245 $Y2=2.802
r259 30 32 16.6411 $w=4.58e-07 $l=6.4e-07 $layer=LI1_cond $X=1.245 $Y=2.625
+ $X2=1.245 $Y2=1.985
r260 29 53 4.82016 $w=3.67e-07 $l=3.65377e-07 $layer=LI1_cond $X=1.245 $Y=1.95
+ $X2=1.39 $Y2=1.65
r261 29 32 0.91006 $w=4.58e-07 $l=3.5e-08 $layer=LI1_cond $X=1.245 $Y=1.95
+ $X2=1.245 $Y2=1.985
r262 26 50 50.1894 $w=3.66e-07 $l=3.02903e-07 $layer=POLY_cond $X=5.55 $Y=2.465
+ $X2=5.667 $Y2=2.215
r263 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.55 $Y=2.465
+ $X2=5.55 $Y2=2.75
r264 22 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.125 $Y=1.15
+ $X2=5.125 $Y2=1.315
r265 22 24 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=5.125 $Y=1.15
+ $X2=5.125 $Y2=0.65
r266 18 20 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.465 $Y=0.255
+ $X2=3.465 $Y2=0.715
r267 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.615 $Y=2.07
+ $X2=2.615 $Y2=2.355
r268 14 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.615 $Y=1.98
+ $X2=2.615 $Y2=2.07
r269 13 14 54.4194 $w=1.8e-07 $l=1.4e-07 $layer=POLY_cond $X=2.615 $Y=1.84
+ $X2=2.615 $Y2=1.98
r270 12 76 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.76 $Y=1.765
+ $X2=1.58 $Y2=1.765
r271 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.525 $Y=1.765
+ $X2=2.615 $Y2=1.84
r272 11 12 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.525 $Y=1.765
+ $X2=1.76 $Y2=1.765
r273 9 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.39 $Y=0.18
+ $X2=3.465 $Y2=0.255
r274 9 10 835.809 $w=1.5e-07 $l=1.63e-06 $layer=POLY_cond $X=3.39 $Y=0.18
+ $X2=1.76 $Y2=0.18
r275 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.685 $Y=0.255
+ $X2=1.76 $Y2=0.18
r276 7 75 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=1.685 $Y=0.255
+ $X2=1.685 $Y2=1.35
r277 2 58 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.815
r278 2 32 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=1.985
r279 1 35 182 $w=1.7e-07 $l=5.9397e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.37 $X2=1.39 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__DFXTP_2%A_695_459# 1 2 7 9 11 14 18 20 25 26 30 36
c86 26 0 1.31176e-19 $X=4.565 $Y=2.125
c87 14 0 1.80864e-19 $X=3.855 $Y=0.715
c88 11 0 5.9515e-20 $X=3.755 $Y=2.295
r89 28 30 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.475 $Y=2.29
+ $X2=4.565 $Y2=2.29
r90 26 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.565 $Y=2.125
+ $X2=4.565 $Y2=2.29
r91 25 26 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.565 $Y=1.415
+ $X2=4.565 $Y2=2.125
r92 23 36 38.0101 $w=2.98e-07 $l=2.35e-07 $layer=POLY_cond $X=4.09 $Y=1.25
+ $X2=3.855 $Y2=1.25
r93 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.09
+ $Y=1.25 $X2=4.09 $Y2=1.25
r94 20 25 10.1681 $w=2.93e-07 $l=2.31633e-07 $layer=LI1_cond $X=4.48 $Y=1.222
+ $X2=4.565 $Y2=1.415
r95 20 33 18.8205 $w=2.93e-07 $l=5.81849e-07 $layer=LI1_cond $X=4.48 $Y=1.222
+ $X2=4.777 $Y2=0.77
r96 20 22 11.6741 $w=3.83e-07 $l=3.9e-07 $layer=LI1_cond $X=4.48 $Y=1.222
+ $X2=4.09 $Y2=1.222
r97 16 18 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.565 $Y=2.37
+ $X2=3.755 $Y2=2.37
r98 12 36 18.8112 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.085
+ $X2=3.855 $Y2=1.25
r99 12 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.855 $Y=1.085
+ $X2=3.855 $Y2=0.715
r100 11 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.755 $Y=2.295
+ $X2=3.755 $Y2=2.37
r101 10 36 16.1745 $w=2.98e-07 $l=2.09105e-07 $layer=POLY_cond $X=3.755 $Y=1.415
+ $X2=3.855 $Y2=1.25
r102 10 11 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.755 $Y=1.415
+ $X2=3.755 $Y2=2.295
r103 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.565 $Y=2.445
+ $X2=3.565 $Y2=2.37
r104 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.565 $Y=2.445
+ $X2=3.565 $Y2=2.73
r105 2 28 600 $w=1.7e-07 $l=2.35053e-07 $layer=licon1_PDIFF $count=1 $X=4.32
+ $Y=2.12 $X2=4.475 $Y2=2.29
r106 1 33 182 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_NDIFF $count=1 $X=4.77
+ $Y=0.375 $X2=4.91 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LS__DFXTP_2%A_538_429# 1 2 7 9 11 12 14 17 21 24 26 27
+ 28 34 39 44 48
c105 39 0 1.80864e-19 $X=3.225 $Y=0.78
c106 24 0 2.36837e-19 $X=3.115 $Y=1.49
r107 48 49 44.0028 $w=3.56e-07 $l=3.25e-07 $layer=POLY_cond $X=4.245 $Y=1.835
+ $X2=4.57 $Y2=1.835
r108 45 48 5.41573 $w=3.56e-07 $l=4e-08 $layer=POLY_cond $X=4.205 $Y=1.835
+ $X2=4.245 $Y2=1.835
r109 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.205
+ $Y=1.79 $X2=4.205 $Y2=1.79
r110 41 44 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=4.05 $Y=1.79
+ $X2=4.205 $Y2=1.79
r111 36 39 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.115 $Y=0.78
+ $X2=3.225 $Y2=0.78
r112 32 34 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.87 $Y=1.575
+ $X2=3.115 $Y2=1.575
r113 27 30 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=2.855 $Y=2.34
+ $X2=2.855 $Y2=2.355
r114 27 28 12.2041 $w=1.98e-07 $l=2.15e-07 $layer=LI1_cond $X=2.855 $Y=2.34
+ $X2=2.855 $Y2=2.125
r115 25 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=1.955
+ $X2=4.05 $Y2=1.79
r116 25 26 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.05 $Y=1.955
+ $X2=4.05 $Y2=2.255
r117 24 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=1.49
+ $X2=3.115 $Y2=1.575
r118 23 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=0.945
+ $X2=3.115 $Y2=0.78
r119 23 24 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.115 $Y=0.945
+ $X2=3.115 $Y2=1.49
r120 22 27 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.955 $Y=2.34
+ $X2=2.855 $Y2=2.34
r121 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.965 $Y=2.34
+ $X2=4.05 $Y2=2.255
r122 21 22 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.965 $Y=2.34
+ $X2=2.955 $Y2=2.34
r123 19 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=1.66
+ $X2=2.87 $Y2=1.575
r124 19 28 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.87 $Y=1.66
+ $X2=2.87 $Y2=2.125
r125 15 17 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=4.57 $Y=1.075
+ $X2=4.695 $Y2=1.075
r126 12 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.695 $Y=1
+ $X2=4.695 $Y2=1.075
r127 12 14 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.695 $Y=1
+ $X2=4.695 $Y2=0.65
r128 11 49 23.0368 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.57 $Y=1.625
+ $X2=4.57 $Y2=1.835
r129 10 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.57 $Y=1.15
+ $X2=4.57 $Y2=1.075
r130 10 11 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=4.57 $Y=1.15
+ $X2=4.57 $Y2=1.625
r131 7 48 23.0368 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.245 $Y=2.045
+ $X2=4.245 $Y2=1.835
r132 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.245 $Y=2.045
+ $X2=4.245 $Y2=2.54
r133 2 30 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=2.69
+ $Y=2.145 $X2=2.84 $Y2=2.355
r134 1 39 182 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.595 $X2=3.225 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LS__DFXTP_2%A_1217_314# 1 2 9 11 13 14 16 19 21 23 26 30
+ 33 37 41 45 47 48 52 53 54 56 58 65
c136 65 0 1.78913e-19 $X=8.135 $Y=1.557
c137 53 0 2.92783e-19 $X=6.25 $Y=1.735
c138 9 0 6.36416e-20 $X=6.175 $Y=0.83
r139 65 66 1.3027 $w=3.7e-07 $l=1e-08 $layer=POLY_cond $X=8.135 $Y=1.557
+ $X2=8.145 $Y2=1.557
r140 64 65 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=7.715 $Y=1.557
+ $X2=8.135 $Y2=1.557
r141 63 64 3.90811 $w=3.7e-07 $l=3e-08 $layer=POLY_cond $X=7.685 $Y=1.557
+ $X2=7.715 $Y2=1.557
r142 57 63 5.21081 $w=3.7e-07 $l=4e-08 $layer=POLY_cond $X=7.645 $Y=1.557
+ $X2=7.685 $Y2=1.557
r143 56 59 8.8128 $w=3.38e-07 $l=2.6e-07 $layer=LI1_cond $X=7.595 $Y=1.515
+ $X2=7.595 $Y2=1.775
r144 56 58 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=7.595 $Y=1.515
+ $X2=7.595 $Y2=1.35
r145 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.645
+ $Y=1.515 $X2=7.645 $Y2=1.515
r146 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.25
+ $Y=1.735 $X2=6.25 $Y2=1.735
r147 49 58 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.51 $Y=1.02
+ $X2=7.51 $Y2=1.35
r148 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.425 $Y=0.935
+ $X2=7.51 $Y2=1.02
r149 47 48 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.425 $Y=0.935
+ $X2=7.115 $Y2=0.935
r150 46 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.04 $Y=1.775
+ $X2=6.915 $Y2=1.775
r151 45 59 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=7.425 $Y=1.775
+ $X2=7.595 $Y2=1.775
r152 45 46 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.425 $Y=1.775
+ $X2=7.04 $Y2=1.775
r153 41 43 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=6.915 $Y=1.985
+ $X2=6.915 $Y2=2.695
r154 39 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.915 $Y=1.86
+ $X2=6.915 $Y2=1.775
r155 39 41 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.915 $Y=1.86
+ $X2=6.915 $Y2=1.985
r156 35 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.95 $Y=0.85
+ $X2=7.115 $Y2=0.935
r157 35 37 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=6.95 $Y=0.85
+ $X2=6.95 $Y2=0.645
r158 34 52 4.72267 $w=1.7e-07 $l=1.92678e-07 $layer=LI1_cond $X=6.415 $Y=1.775
+ $X2=6.25 $Y2=1.715
r159 33 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.79 $Y=1.775
+ $X2=6.915 $Y2=1.775
r160 33 34 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.79 $Y=1.775
+ $X2=6.415 $Y2=1.775
r161 30 53 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.25 $Y=2.075
+ $X2=6.25 $Y2=1.735
r162 29 53 43.7316 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.25 $Y=1.57
+ $X2=6.25 $Y2=1.735
r163 24 66 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.145 $Y=1.35
+ $X2=8.145 $Y2=1.557
r164 24 26 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.145 $Y=1.35
+ $X2=8.145 $Y2=0.74
r165 21 65 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.135 $Y=1.765
+ $X2=8.135 $Y2=1.557
r166 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.135 $Y=1.765
+ $X2=8.135 $Y2=2.4
r167 17 64 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.715 $Y=1.35
+ $X2=7.715 $Y2=1.557
r168 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.715 $Y=1.35
+ $X2=7.715 $Y2=0.74
r169 14 63 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.685 $Y=1.765
+ $X2=7.685 $Y2=1.557
r170 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.685 $Y=1.765
+ $X2=7.685 $Y2=2.4
r171 11 30 77.358 $w=2.43e-07 $l=4.25852e-07 $layer=POLY_cond $X=6.175 $Y=2.465
+ $X2=6.25 $Y2=2.075
r172 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.175 $Y=2.465
+ $X2=6.175 $Y2=2.75
r173 9 29 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.175 $Y=0.83
+ $X2=6.175 $Y2=1.57
r174 2 43 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=1.84 $X2=6.955 $Y2=2.695
r175 2 41 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=1.84 $X2=6.955 $Y2=1.985
r176 1 37 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=6.805
+ $Y=0.37 $X2=6.95 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__DFXTP_2%A_1019_424# 1 2 9 12 13 15 18 20 24 25 27 29
+ 32 34 35 36
c106 36 0 1.43814e-19 $X=6.91 $Y=1.355
c107 34 0 1.78913e-19 $X=7.075 $Y=1.355
c108 29 0 1.52685e-19 $X=5.67 $Y=1.71
c109 25 0 1.79753e-19 $X=5.33 $Y=1.795
c110 24 0 2.31098e-19 $X=5.585 $Y=1.795
c111 9 0 2.55617e-20 $X=7.165 $Y=0.645
r112 35 40 40.8642 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.09 $Y=1.355
+ $X2=7.09 $Y2=1.52
r113 35 39 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.09 $Y=1.355
+ $X2=7.09 $Y2=1.19
r114 34 36 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.075 $Y=1.355
+ $X2=6.91 $Y2=1.355
r115 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.075
+ $Y=1.355 $X2=7.075 $Y2=1.355
r116 31 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.755 $Y=1.315
+ $X2=5.67 $Y2=1.315
r117 31 36 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=5.755 $Y=1.315
+ $X2=6.91 $Y2=1.315
r118 28 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.67 $Y=1.4 $X2=5.67
+ $Y2=1.315
r119 28 29 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.67 $Y=1.4
+ $X2=5.67 $Y2=1.71
r120 27 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.67 $Y=1.23
+ $X2=5.67 $Y2=1.315
r121 26 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.67 $Y=0.945
+ $X2=5.67 $Y2=1.23
r122 24 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.585 $Y=1.795
+ $X2=5.67 $Y2=1.71
r123 24 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.585 $Y=1.795
+ $X2=5.33 $Y2=1.795
r124 20 26 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.585 $Y=0.82
+ $X2=5.67 $Y2=0.945
r125 20 22 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=5.585 $Y=0.82
+ $X2=5.49 $Y2=0.82
r126 16 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.245 $Y=1.88
+ $X2=5.33 $Y2=1.795
r127 16 18 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.245 $Y=1.88
+ $X2=5.245 $Y2=2.495
r128 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.18 $Y=1.765
+ $X2=7.18 $Y2=2.34
r129 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.18 $Y=1.675
+ $X2=7.18 $Y2=1.765
r130 12 40 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=7.18 $Y=1.675
+ $X2=7.18 $Y2=1.52
r131 9 39 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.165 $Y=0.645
+ $X2=7.165 $Y2=1.19
r132 2 18 600 $w=1.7e-07 $l=4.43706e-07 $layer=licon1_PDIFF $count=1 $X=5.095
+ $Y=2.12 $X2=5.245 $Y2=2.495
r133 1 22 182 $w=1.7e-07 $l=5.30542e-07 $layer=licon1_NDIFF $count=1 $X=5.2
+ $Y=0.375 $X2=5.49 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LS__DFXTP_2%VPWR 1 2 3 4 5 6 23 27 31 33 35 39 41 46 54
+ 59 64 70 73 80 87 90 94
r105 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r106 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r107 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r108 83 84 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r109 80 83 8.27395 $w=3.88e-07 $l=2.8e-07 $layer=LI1_cond $X=3.905 $Y=3.05
+ $X2=3.905 $Y2=3.33
r110 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r111 73 76 8.96345 $w=3.58e-07 $l=2.8e-07 $layer=LI1_cond $X=1.755 $Y=3.05
+ $X2=1.755 $Y2=3.33
r112 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 68 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r114 68 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r115 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r116 65 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.57 $Y=3.33
+ $X2=7.405 $Y2=3.33
r117 65 67 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.57 $Y=3.33
+ $X2=7.92 $Y2=3.33
r118 64 93 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.275 $Y=3.33
+ $X2=8.457 $Y2=3.33
r119 64 67 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.275 $Y=3.33
+ $X2=7.92 $Y2=3.33
r120 63 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r121 63 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r122 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r123 60 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.565 $Y=3.33
+ $X2=6.4 $Y2=3.33
r124 60 62 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.565 $Y=3.33
+ $X2=6.96 $Y2=3.33
r125 59 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.24 $Y=3.33
+ $X2=7.405 $Y2=3.33
r126 59 62 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.24 $Y=3.33
+ $X2=6.96 $Y2=3.33
r127 58 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r128 57 58 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r129 55 83 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.1 $Y=3.33
+ $X2=3.905 $Y2=3.33
r130 55 57 123.957 $w=1.68e-07 $l=1.9e-06 $layer=LI1_cond $X=4.1 $Y=3.33 $X2=6
+ $Y2=3.33
r131 54 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.235 $Y=3.33
+ $X2=6.4 $Y2=3.33
r132 54 57 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.235 $Y=3.33
+ $X2=6 $Y2=3.33
r133 53 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r134 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r135 50 53 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r136 50 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r137 49 52 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r138 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r139 47 76 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=1.755 $Y2=3.33
r140 47 49 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=2.16 $Y2=3.33
r141 46 83 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.71 $Y=3.33
+ $X2=3.905 $Y2=3.33
r142 46 52 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.71 $Y=3.33
+ $X2=3.6 $Y2=3.33
r143 45 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r144 45 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r145 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r146 42 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.73 $Y2=3.33
r147 42 44 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r148 41 76 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.755 $Y2=3.33
r149 41 44 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r150 39 58 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=6 $Y2=3.33
r151 39 84 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r152 35 38 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.4 $Y=1.985
+ $X2=8.4 $Y2=2.815
r153 33 93 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.4 $Y=3.245
+ $X2=8.457 $Y2=3.33
r154 33 38 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.4 $Y=3.245 $X2=8.4
+ $Y2=2.815
r155 29 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.405 $Y=3.245
+ $X2=7.405 $Y2=3.33
r156 29 31 36.6686 $w=3.28e-07 $l=1.05e-06 $layer=LI1_cond $X=7.405 $Y=3.245
+ $X2=7.405 $Y2=2.195
r157 25 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=3.245 $X2=6.4
+ $Y2=3.33
r158 25 27 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=6.4 $Y=3.245
+ $X2=6.4 $Y2=2.75
r159 21 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r160 21 23 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.455
r161 6 38 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.84 $X2=8.36 $Y2=2.815
r162 6 35 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.84 $X2=8.36 $Y2=1.985
r163 5 31 300 $w=1.7e-07 $l=4.23409e-07 $layer=licon1_PDIFF $count=2 $X=7.255
+ $Y=1.84 $X2=7.405 $Y2=2.195
r164 4 27 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=6.25
+ $Y=2.54 $X2=6.4 $Y2=2.75
r165 3 80 600 $w=1.7e-07 $l=6.49115e-07 $layer=licon1_PDIFF $count=1 $X=3.64
+ $Y=2.52 $X2=3.905 $Y2=3.05
r166 2 73 600 $w=1.7e-07 $l=5.84551e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=2.54 $X2=1.755 $Y2=3.05
r167 1 23 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__DFXTP_2%A_431_508# 1 2 9 15 17 18 21
c45 9 0 6.76432e-20 $X=2.39 $Y=2.29
r46 19 21 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.53 $Y=1.235
+ $X2=2.775 $Y2=1.235
r47 17 18 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.42 $Y=1.65
+ $X2=2.42 $Y2=1.82
r48 13 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=1.15
+ $X2=2.775 $Y2=1.235
r49 13 15 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.775 $Y=1.15
+ $X2=2.775 $Y2=0.815
r50 11 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=1.32
+ $X2=2.53 $Y2=1.235
r51 11 17 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.53 $Y=1.32
+ $X2=2.53 $Y2=1.65
r52 9 18 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=2.39 $Y=2.29 $X2=2.39
+ $Y2=1.82
r53 2 9 600 $w=1.7e-07 $l=3.4821e-07 $layer=licon1_PDIFF $count=1 $X=2.155
+ $Y=2.54 $X2=2.39 $Y2=2.29
r54 1 15 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.635
+ $Y=0.595 $X2=2.775 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LS__DFXTP_2%Q 1 2 9 15 16 17 18 19
c35 17 0 2.55617e-20 $X=7.935 $Y=1.13
r36 18 19 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=7.925 $Y=2.405
+ $X2=7.925 $Y2=2.775
r37 16 17 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=8.02 $Y=2.03 $X2=8.02
+ $Y2=1.13
r38 15 16 6.59029 $w=3.58e-07 $l=1.05e-07 $layer=LI1_cond $X=7.925 $Y=2.135
+ $X2=7.925 $Y2=2.03
r39 13 18 6.2424 $w=3.58e-07 $l=1.95e-07 $layer=LI1_cond $X=7.925 $Y=2.21
+ $X2=7.925 $Y2=2.405
r40 13 15 2.40092 $w=3.58e-07 $l=7.5e-08 $layer=LI1_cond $X=7.925 $Y=2.21
+ $X2=7.925 $Y2=2.135
r41 7 17 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=7.935 $Y=0.96
+ $X2=7.935 $Y2=1.13
r42 7 9 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=7.935 $Y=0.96
+ $X2=7.935 $Y2=0.515
r43 2 19 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=1.84 $X2=7.91 $Y2=2.815
r44 2 15 400 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=1.84 $X2=7.91 $Y2=2.135
r45 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.79
+ $Y=0.37 $X2=7.93 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DFXTP_2%VGND 1 2 3 4 5 6 21 25 29 33 37 39 41 44 45
+ 46 48 53 58 70 74 80 83 86 89 93
r116 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r117 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r118 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r119 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r120 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r121 78 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r122 78 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r123 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r124 75 89 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.447 $Y2=0
r125 75 77 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.92 $Y2=0
r126 74 92 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.275 $Y=0
+ $X2=8.457 $Y2=0
r127 74 77 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.275 $Y=0
+ $X2=7.92 $Y2=0
r128 73 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r129 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r130 70 89 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=7.3 $Y=0 $X2=7.447
+ $Y2=0
r131 70 72 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.3 $Y=0 $X2=6.96
+ $Y2=0
r132 69 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r133 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r134 66 69 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r135 65 68 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r136 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r137 63 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.235 $Y=0 $X2=4.11
+ $Y2=0
r138 63 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.235 $Y=0
+ $X2=4.56 $Y2=0
r139 62 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r140 62 84 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.16
+ $Y2=0
r141 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r142 59 83 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.082
+ $Y2=0
r143 59 61 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=2.18 $Y=0 $X2=3.6
+ $Y2=0
r144 58 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.985 $Y=0 $X2=4.11
+ $Y2=0
r145 58 61 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.985 $Y=0 $X2=3.6
+ $Y2=0
r146 57 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r147 57 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r148 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r149 54 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.67
+ $Y2=0
r150 54 56 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.68
+ $Y2=0
r151 53 83 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=1.985 $Y=0 $X2=2.082
+ $Y2=0
r152 53 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=0
+ $X2=1.68 $Y2=0
r153 51 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r154 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r155 48 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.67
+ $Y2=0
r156 48 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r157 46 66 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r158 46 87 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r159 44 68 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.225 $Y=0 $X2=6
+ $Y2=0
r160 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.225 $Y=0 $X2=6.39
+ $Y2=0
r161 43 72 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.555 $Y=0
+ $X2=6.96 $Y2=0
r162 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.555 $Y=0 $X2=6.39
+ $Y2=0
r163 39 92 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.4 $Y=0.085
+ $X2=8.457 $Y2=0
r164 39 41 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.4 $Y=0.085 $X2=8.4
+ $Y2=0.515
r165 35 89 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=7.447 $Y=0.085
+ $X2=7.447 $Y2=0
r166 35 37 16.7983 $w=2.93e-07 $l=4.3e-07 $layer=LI1_cond $X=7.447 $Y=0.085
+ $X2=7.447 $Y2=0.515
r167 31 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=0.085
+ $X2=6.39 $Y2=0
r168 31 33 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=6.39 $Y=0.085
+ $X2=6.39 $Y2=0.83
r169 27 86 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=0.085
+ $X2=4.11 $Y2=0
r170 27 29 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=4.11 $Y=0.085
+ $X2=4.11 $Y2=0.355
r171 23 83 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.082 $Y=0.085
+ $X2=2.082 $Y2=0
r172 23 25 22.1818 $w=1.93e-07 $l=3.9e-07 $layer=LI1_cond $X=2.082 $Y=0.085
+ $X2=2.082 $Y2=0.475
r173 19 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r174 19 21 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.57
r175 6 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.22
+ $Y=0.37 $X2=8.36 $Y2=0.515
r176 5 37 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=7.24
+ $Y=0.37 $X2=7.405 $Y2=0.515
r177 4 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.25
+ $Y=0.62 $X2=6.39 $Y2=0.83
r178 3 29 182 $w=1.7e-07 $l=2.85307e-07 $layer=licon1_NDIFF $count=1 $X=3.93
+ $Y=0.505 $X2=4.15 $Y2=0.355
r179 2 25 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.33 $X2=2.08 $Y2=0.475
r180 1 21 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.57
.ends

