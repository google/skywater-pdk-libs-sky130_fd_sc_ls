* File: sky130_fd_sc_ls__a311o_1.spice
* Created: Fri Aug 28 12:57:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a311o_1.pex.spice"
.subckt sky130_fd_sc_ls__a311o_1  VNB VPB A3 A2 A1 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_89_270#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.74
+ AD=0.137758 AS=0.1961 PD=1.17971 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1001 A_264_120# N_A3_M1001_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.64
+ AD=0.105312 AS=0.119142 PD=0.98 PS=1.02029 NRD=20.532 NRS=14.988 M=1 R=4.26667
+ SA=75000.7 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1008 A_359_123# N_A2_M1008_g A_264_120# VNB NSHORT L=0.15 W=0.64 AD=0.1024
+ AS=0.105312 PD=0.96 PS=0.98 NRD=19.68 NRS=20.532 M=1 R=4.26667 SA=75001.2
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1004 N_A_89_270#_M1004_d N_A1_M1004_g A_359_123# VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1024 PD=0.92 PS=0.96 NRD=0 NRS=19.68 M=1 R=4.26667 SA=75001.6
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_B1_M1011_g N_A_89_270#_M1004_d VNB NSHORT L=0.15 W=0.64
+ AD=0.136 AS=0.0896 PD=1.065 PS=0.92 NRD=14.988 NRS=0 M=1 R=4.26667 SA=75002.1
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1000 N_A_89_270#_M1000_d N_C1_M1000_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1696 AS=0.136 PD=1.81 PS=1.065 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75002.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1010 N_VPWR_M1010_d N_A_89_270#_M1010_g N_X_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2968 AS=0.308 PD=1.7434 PS=2.79 NRD=21.9852 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1009 N_A_258_392#_M1009_d N_A3_M1009_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.265 PD=1.3 PS=1.5566 NRD=1.9503 NRS=24.6053 M=1 R=6.66667
+ SA=75000.9 SB=75002 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_258_392#_M1009_d VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.15 PD=1.39 PS=1.3 NRD=5.8903 NRS=1.9503 M=1 R=6.66667 SA=75001.3
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1005 N_A_258_392#_M1005_d N_A1_M1005_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.195 PD=1.3 PS=1.39 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75001.9 SB=75001 A=0.15 P=2.3 MULT=1
MM1006 A_546_392# N_B1_M1006_g N_A_258_392#_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.12 AS=0.15 PD=1.24 PS=1.3 NRD=12.7853 NRS=1.9503 M=1 R=6.66667 SA=75002.3
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1007 N_A_89_270#_M1007_d N_C1_M1007_g A_546_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.275 AS=0.12 PD=2.55 PS=1.24 NRD=1.9503 NRS=12.7853 M=1 R=6.66667
+ SA=75002.7 SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ls__a311o_1.pxi.spice"
*
.ends
*
*
