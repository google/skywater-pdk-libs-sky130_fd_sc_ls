* File: sky130_fd_sc_ls__clkdlyinv5sd3_1.pxi.spice
* Created: Fri Aug 28 13:10:20 2020
* 
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%A N_A_M1007_g N_A_c_74_n N_A_c_78_n
+ N_A_M1009_g A A N_A_c_76_n PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%A
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%A_28_74# N_A_28_74#_M1007_s
+ N_A_28_74#_M1009_s N_A_28_74#_c_110_n N_A_28_74#_M1002_g N_A_28_74#_c_111_n
+ N_A_28_74#_M1005_g N_A_28_74#_c_113_n N_A_28_74#_c_117_n N_A_28_74#_c_118_n
+ N_A_28_74#_c_129_n N_A_28_74#_c_114_n N_A_28_74#_c_115_n N_A_28_74#_c_137_n
+ PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%A_28_74#
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%A_288_74# N_A_288_74#_M1002_d
+ N_A_288_74#_M1005_d N_A_288_74#_c_168_n N_A_288_74#_c_169_n
+ N_A_288_74#_c_170_n N_A_288_74#_c_174_n N_A_288_74#_c_171_n
+ N_A_288_74#_M1006_g N_A_288_74#_M1001_g
+ PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%A_288_74#
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%A_549_74# N_A_549_74#_M1006_d
+ N_A_549_74#_M1001_d N_A_549_74#_c_206_n N_A_549_74#_M1004_g
+ N_A_549_74#_M1008_g N_A_549_74#_c_209_n N_A_549_74#_c_210_n
+ N_A_549_74#_c_211_n N_A_549_74#_c_212_n
+ PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%A_549_74#
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%A_682_74# N_A_682_74#_M1008_s
+ N_A_682_74#_M1004_s N_A_682_74#_M1003_g N_A_682_74#_c_254_n
+ N_A_682_74#_M1000_g N_A_682_74#_c_255_n N_A_682_74#_c_262_n
+ N_A_682_74#_c_256_n N_A_682_74#_c_257_n N_A_682_74#_c_258_n
+ N_A_682_74#_c_259_n N_A_682_74#_c_260_n
+ PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%A_682_74#
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%VPWR N_VPWR_M1009_d N_VPWR_M1001_s
+ N_VPWR_M1004_d N_VPWR_c_309_n N_VPWR_c_310_n N_VPWR_c_311_n VPWR
+ N_VPWR_c_312_n N_VPWR_c_313_n N_VPWR_c_314_n N_VPWR_c_315_n N_VPWR_c_308_n
+ N_VPWR_c_317_n N_VPWR_c_318_n N_VPWR_c_319_n VPWR
+ PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%VPWR
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%Y N_Y_M1003_d N_Y_M1000_d Y Y Y Y Y Y Y Y
+ PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%Y
x_PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%VGND N_VGND_M1007_d N_VGND_M1006_s
+ N_VGND_M1008_d N_VGND_c_372_n N_VGND_c_373_n N_VGND_c_374_n VGND
+ N_VGND_c_375_n N_VGND_c_376_n N_VGND_c_377_n N_VGND_c_378_n N_VGND_c_379_n
+ N_VGND_c_380_n N_VGND_c_381_n N_VGND_c_382_n VGND
+ PM_SKY130_FD_SC_LS__CLKDLYINV5SD3_1%VGND
cc_1 VNB N_A_M1007_g 0.0436663f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.58
cc_2 VNB N_A_c_74_n 0.00890285f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.675
cc_3 VNB A 0.0265853f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A_c_76_n 0.035867f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_5 VNB N_A_28_74#_c_110_n 0.0390458f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_6 VNB N_A_28_74#_c_111_n 0.048705f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_A_28_74#_M1005_g 0.0269704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_28_74#_c_113_n 0.0226356f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_9 VNB N_A_28_74#_c_114_n 0.0123049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_28_74#_c_115_n 0.0121635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_288_74#_c_168_n 0.0172077f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_12 VNB N_A_288_74#_c_169_n 0.00548306f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_13 VNB N_A_288_74#_c_170_n 0.0255344f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.19
cc_14 VNB N_A_288_74#_c_171_n 0.00614775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_288_74#_M1006_g 0.128182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_549_74#_c_206_n 0.0609527f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_17 VNB N_A_549_74#_M1004_g 0.0116394f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_18 VNB N_A_549_74#_M1008_g 0.0602032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_549_74#_c_209_n 0.0155677f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.19
cc_20 VNB N_A_549_74#_c_210_n 0.0111173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_549_74#_c_211_n 0.0373197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_549_74#_c_212_n 0.00227058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_682_74#_M1003_g 0.0444659f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_24 VNB N_A_682_74#_c_254_n 0.0391593f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_25 VNB N_A_682_74#_c_255_n 0.00645043f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_26 VNB N_A_682_74#_c_256_n 0.00438081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_682_74#_c_257_n 0.00366902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_682_74#_c_258_n 0.0134028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_682_74#_c_259_n 0.00543637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_682_74#_c_260_n 0.00272046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_308_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB Y 0.0204118f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_33 VNB Y 0.0466962f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_34 VNB N_VGND_c_372_n 0.00963665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_373_n 0.0113129f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_36 VNB N_VGND_c_374_n 0.00662038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_375_n 0.0180717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_376_n 0.0296852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_377_n 0.0620127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_378_n 0.0189455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_379_n 0.315628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_380_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_381_n 0.00654723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_382_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_A_c_74_n 8.9669e-19 $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.675
cc_46 VPB N_A_c_78_n 0.0271587f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_47 VPB A 0.0105602f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_48 VPB N_A_28_74#_M1005_g 0.0608692f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_28_74#_c_117_n 0.0079884f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.52
cc_50 VPB N_A_28_74#_c_118_n 0.0205617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_288_74#_c_169_n 0.0145364f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.355
cc_52 VPB N_A_288_74#_c_174_n 0.00255514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_288_74#_M1006_g 0.0663125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_549_74#_M1004_g 0.0643005f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_55 VPB N_A_549_74#_c_210_n 0.0106835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_682_74#_c_254_n 0.0254953f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_57 VPB N_A_682_74#_c_262_n 0.00826349f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_682_74#_c_256_n 0.00876445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_682_74#_c_257_n 9.90711e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_309_n 0.00996699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_310_n 0.0220323f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.355
cc_62 VPB N_VPWR_c_311_n 0.00777218f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.355
cc_63 VPB N_VPWR_c_312_n 0.018958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_313_n 0.0298867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_314_n 0.0623064f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_315_n 0.0184442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_308_n 0.0946668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_317_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_318_n 0.00652134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_319_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB Y 0.0121098f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_72 VPB Y 0.0526708f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_73 A N_A_28_74#_M1009_s 0.00256075f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A_M1007_g N_A_28_74#_c_110_n 0.0151729f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_75 N_A_M1007_g N_A_28_74#_c_111_n 0.0021171f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_76 A N_A_28_74#_c_111_n 0.00125289f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A_c_76_n N_A_28_74#_c_111_n 0.0208561f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_78 N_A_c_74_n N_A_28_74#_M1005_g 0.00769658f $X=0.495 $Y=1.675 $X2=0 $Y2=0
cc_79 N_A_c_78_n N_A_28_74#_M1005_g 0.0299649f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_80 A N_A_28_74#_M1005_g 0.00301665f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A_M1007_g N_A_28_74#_c_113_n 0.00871827f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_82 A N_A_28_74#_c_117_n 0.0237727f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A_c_78_n N_A_28_74#_c_129_n 0.0136074f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_84 A N_A_28_74#_c_129_n 0.0197054f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A_c_76_n N_A_28_74#_c_129_n 6.00585e-19 $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_86 N_A_M1007_g N_A_28_74#_c_114_n 0.010935f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_87 A N_A_28_74#_c_114_n 0.0251751f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_88 N_A_c_76_n N_A_28_74#_c_114_n 0.00146806f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_89 N_A_M1007_g N_A_28_74#_c_115_n 0.00415005f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_90 A N_A_28_74#_c_115_n 0.0289843f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A_M1007_g N_A_28_74#_c_137_n 9.21332e-19 $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_92 N_A_c_74_n N_A_28_74#_c_137_n 2.44702e-19 $X=0.495 $Y=1.675 $X2=0 $Y2=0
cc_93 N_A_c_78_n N_A_28_74#_c_137_n 0.00102987f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_94 A N_A_28_74#_c_137_n 0.0410047f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_95 N_A_c_76_n N_A_28_74#_c_137_n 0.00110237f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_96 A N_VPWR_M1009_d 0.00133607f $X=0.155 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_97 N_A_c_78_n N_VPWR_c_309_n 0.00387645f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A_c_78_n N_VPWR_c_312_n 0.00461464f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_c_78_n N_VPWR_c_308_n 0.00911783f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A_M1007_g N_VGND_c_372_n 0.00248511f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_101 N_A_M1007_g N_VGND_c_375_n 0.00456766f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_102 N_A_M1007_g N_VGND_c_379_n 0.00454566f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_103 N_A_28_74#_c_110_n N_A_288_74#_c_168_n 0.0133513f $X=1.19 $Y=0.88 $X2=0
+ $Y2=0
cc_104 N_A_28_74#_c_111_n N_A_288_74#_c_168_n 2.87835e-19 $X=1.195 $Y=1.38 $X2=0
+ $Y2=0
cc_105 N_A_28_74#_c_114_n N_A_288_74#_c_168_n 0.01637f $X=0.975 $Y=0.92 $X2=0
+ $Y2=0
cc_106 N_A_28_74#_c_137_n N_A_288_74#_c_168_n 0.0091978f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_107 N_A_28_74#_M1005_g N_A_288_74#_c_169_n 0.0142889f $X=1.195 $Y=2.46 $X2=0
+ $Y2=0
cc_108 N_A_28_74#_c_137_n N_A_288_74#_c_169_n 0.0406706f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_109 N_A_28_74#_M1005_g N_A_288_74#_c_174_n 0.0079719f $X=1.195 $Y=2.46 $X2=0
+ $Y2=0
cc_110 N_A_28_74#_c_111_n N_A_288_74#_c_171_n 0.00987877f $X=1.195 $Y=1.38 $X2=0
+ $Y2=0
cc_111 N_A_28_74#_c_137_n N_A_288_74#_c_171_n 0.0277877f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_112 N_A_28_74#_c_129_n N_VPWR_M1009_d 0.00987397f $X=0.975 $Y=2.117 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A_28_74#_M1005_g N_VPWR_c_309_n 0.00818817f $X=1.195 $Y=2.46 $X2=0
+ $Y2=0
cc_114 N_A_28_74#_c_129_n N_VPWR_c_309_n 0.0208193f $X=0.975 $Y=2.117 $X2=0
+ $Y2=0
cc_115 N_A_28_74#_M1005_g N_VPWR_c_310_n 0.00488034f $X=1.195 $Y=2.46 $X2=0
+ $Y2=0
cc_116 N_A_28_74#_c_118_n N_VPWR_c_312_n 0.00593336f $X=0.265 $Y=2.56 $X2=0
+ $Y2=0
cc_117 N_A_28_74#_M1005_g N_VPWR_c_313_n 0.0150739f $X=1.195 $Y=2.46 $X2=0 $Y2=0
cc_118 N_A_28_74#_M1005_g N_VPWR_c_308_n 0.0291737f $X=1.195 $Y=2.46 $X2=0 $Y2=0
cc_119 N_A_28_74#_c_118_n N_VPWR_c_308_n 0.00940928f $X=0.265 $Y=2.56 $X2=0
+ $Y2=0
cc_120 N_A_28_74#_c_110_n N_VGND_c_372_n 0.0031236f $X=1.19 $Y=0.88 $X2=0 $Y2=0
cc_121 N_A_28_74#_c_113_n N_VGND_c_372_n 0.0151665f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_122 N_A_28_74#_c_114_n N_VGND_c_372_n 0.0242038f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_123 N_A_28_74#_c_110_n N_VGND_c_373_n 0.00268449f $X=1.19 $Y=0.88 $X2=0 $Y2=0
cc_124 N_A_28_74#_c_113_n N_VGND_c_375_n 0.0170785f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_125 N_A_28_74#_c_110_n N_VGND_c_376_n 0.0153821f $X=1.19 $Y=0.88 $X2=0 $Y2=0
cc_126 N_A_28_74#_c_110_n N_VGND_c_379_n 0.0192653f $X=1.19 $Y=0.88 $X2=0 $Y2=0
cc_127 N_A_28_74#_c_113_n N_VGND_c_379_n 0.0118627f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_128 N_A_28_74#_c_114_n N_VGND_c_379_n 0.0189117f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_129 N_A_288_74#_c_170_n N_A_549_74#_c_209_n 0.00419423f $X=2.425 $Y=1.305
+ $X2=0 $Y2=0
cc_130 N_A_288_74#_M1006_g N_A_549_74#_c_209_n 0.0184465f $X=2.495 $Y=0.58 $X2=0
+ $Y2=0
cc_131 N_A_288_74#_c_170_n N_A_549_74#_c_210_n 0.00419423f $X=2.425 $Y=1.305
+ $X2=0 $Y2=0
cc_132 N_A_288_74#_M1006_g N_A_549_74#_c_210_n 0.0247631f $X=2.495 $Y=0.58 $X2=0
+ $Y2=0
cc_133 N_A_288_74#_c_170_n N_A_549_74#_c_212_n 0.0101411f $X=2.425 $Y=1.305
+ $X2=0 $Y2=0
cc_134 N_A_288_74#_M1006_g N_A_549_74#_c_212_n 0.00534783f $X=2.495 $Y=0.58
+ $X2=0 $Y2=0
cc_135 N_A_288_74#_c_169_n N_VPWR_c_310_n 0.0793701f $X=1.58 $Y=2.105 $X2=0
+ $Y2=0
cc_136 N_A_288_74#_c_170_n N_VPWR_c_310_n 0.0150336f $X=2.425 $Y=1.305 $X2=0
+ $Y2=0
cc_137 N_A_288_74#_M1006_g N_VPWR_c_310_n 0.0348189f $X=2.495 $Y=0.58 $X2=0
+ $Y2=0
cc_138 N_A_288_74#_c_174_n N_VPWR_c_313_n 0.00976575f $X=1.58 $Y=2.815 $X2=0
+ $Y2=0
cc_139 N_A_288_74#_M1006_g N_VPWR_c_314_n 0.0147528f $X=2.495 $Y=0.58 $X2=0
+ $Y2=0
cc_140 N_A_288_74#_c_174_n N_VPWR_c_308_n 0.0112865f $X=1.58 $Y=2.815 $X2=0
+ $Y2=0
cc_141 N_A_288_74#_M1006_g N_VPWR_c_308_n 0.0290091f $X=2.495 $Y=0.58 $X2=0
+ $Y2=0
cc_142 N_A_288_74#_c_168_n N_VGND_c_372_n 0.00224734f $X=1.58 $Y=0.58 $X2=0
+ $Y2=0
cc_143 N_A_288_74#_c_168_n N_VGND_c_373_n 0.0326859f $X=1.58 $Y=0.58 $X2=0 $Y2=0
cc_144 N_A_288_74#_c_170_n N_VGND_c_373_n 0.0150716f $X=2.425 $Y=1.305 $X2=0
+ $Y2=0
cc_145 N_A_288_74#_M1006_g N_VGND_c_373_n 0.0200848f $X=2.495 $Y=0.58 $X2=0
+ $Y2=0
cc_146 N_A_288_74#_c_168_n N_VGND_c_376_n 0.0132196f $X=1.58 $Y=0.58 $X2=0 $Y2=0
cc_147 N_A_288_74#_M1006_g N_VGND_c_377_n 0.0147528f $X=2.495 $Y=0.58 $X2=0
+ $Y2=0
cc_148 N_A_288_74#_c_168_n N_VGND_c_379_n 0.00920999f $X=1.58 $Y=0.58 $X2=0
+ $Y2=0
cc_149 N_A_288_74#_M1006_g N_VGND_c_379_n 0.0290091f $X=2.495 $Y=0.58 $X2=0
+ $Y2=0
cc_150 N_A_549_74#_M1008_g N_A_682_74#_M1003_g 0.0206725f $X=3.925 $Y=0.58 $X2=0
+ $Y2=0
cc_151 N_A_549_74#_c_206_n N_A_682_74#_c_254_n 0.0131837f $X=3.92 $Y=1.545 $X2=0
+ $Y2=0
cc_152 N_A_549_74#_M1004_g N_A_682_74#_c_254_n 0.0207651f $X=3.92 $Y=2.46 $X2=0
+ $Y2=0
cc_153 N_A_549_74#_c_211_n N_A_682_74#_c_254_n 2.99954e-19 $X=3.84 $Y=1.305
+ $X2=0 $Y2=0
cc_154 N_A_549_74#_M1008_g N_A_682_74#_c_255_n 0.0198301f $X=3.925 $Y=0.58 $X2=0
+ $Y2=0
cc_155 N_A_549_74#_c_209_n N_A_682_74#_c_255_n 0.0198272f $X=2.885 $Y=0.58 $X2=0
+ $Y2=0
cc_156 N_A_549_74#_M1004_g N_A_682_74#_c_262_n 0.0111545f $X=3.92 $Y=2.46 $X2=0
+ $Y2=0
cc_157 N_A_549_74#_c_210_n N_A_682_74#_c_262_n 0.046582f $X=2.885 $Y=2.105 $X2=0
+ $Y2=0
cc_158 N_A_549_74#_M1004_g N_A_682_74#_c_256_n 0.0445213f $X=3.92 $Y=2.46 $X2=0
+ $Y2=0
cc_159 N_A_549_74#_c_211_n N_A_682_74#_c_256_n 0.0237983f $X=3.84 $Y=1.305 $X2=0
+ $Y2=0
cc_160 N_A_549_74#_c_210_n N_A_682_74#_c_257_n 0.0073655f $X=2.885 $Y=2.105
+ $X2=0 $Y2=0
cc_161 N_A_549_74#_c_211_n N_A_682_74#_c_257_n 0.0202705f $X=3.84 $Y=1.305 $X2=0
+ $Y2=0
cc_162 N_A_549_74#_c_206_n N_A_682_74#_c_258_n 0.00843713f $X=3.92 $Y=1.545
+ $X2=0 $Y2=0
cc_163 N_A_549_74#_M1008_g N_A_682_74#_c_258_n 0.0303022f $X=3.925 $Y=0.58 $X2=0
+ $Y2=0
cc_164 N_A_549_74#_c_211_n N_A_682_74#_c_258_n 0.0206391f $X=3.84 $Y=1.305 $X2=0
+ $Y2=0
cc_165 N_A_549_74#_c_206_n N_A_682_74#_c_259_n 4.80213e-19 $X=3.92 $Y=1.545
+ $X2=0 $Y2=0
cc_166 N_A_549_74#_M1008_g N_A_682_74#_c_259_n 0.00369944f $X=3.925 $Y=0.58
+ $X2=0 $Y2=0
cc_167 N_A_549_74#_c_209_n N_A_682_74#_c_259_n 0.0079307f $X=2.885 $Y=0.58 $X2=0
+ $Y2=0
cc_168 N_A_549_74#_c_211_n N_A_682_74#_c_259_n 0.0275619f $X=3.84 $Y=1.305 $X2=0
+ $Y2=0
cc_169 N_A_549_74#_c_206_n N_A_682_74#_c_260_n 0.00564593f $X=3.92 $Y=1.545
+ $X2=0 $Y2=0
cc_170 N_A_549_74#_c_211_n N_A_682_74#_c_260_n 0.00545692f $X=3.84 $Y=1.305
+ $X2=0 $Y2=0
cc_171 N_A_549_74#_c_210_n N_VPWR_c_310_n 0.0160312f $X=2.885 $Y=2.105 $X2=0
+ $Y2=0
cc_172 N_A_549_74#_M1004_g N_VPWR_c_311_n 0.0197872f $X=3.92 $Y=2.46 $X2=0 $Y2=0
cc_173 N_A_549_74#_M1004_g N_VPWR_c_314_n 0.0153821f $X=3.92 $Y=2.46 $X2=0 $Y2=0
cc_174 N_A_549_74#_c_210_n N_VPWR_c_314_n 0.00749631f $X=2.885 $Y=2.105 $X2=0
+ $Y2=0
cc_175 N_A_549_74#_M1004_g N_VPWR_c_308_n 0.030237f $X=3.92 $Y=2.46 $X2=0 $Y2=0
cc_176 N_A_549_74#_c_210_n N_VPWR_c_308_n 0.0062048f $X=2.885 $Y=2.105 $X2=0
+ $Y2=0
cc_177 N_A_549_74#_M1008_g N_VGND_c_374_n 0.00843039f $X=3.925 $Y=0.58 $X2=0
+ $Y2=0
cc_178 N_A_549_74#_M1008_g N_VGND_c_377_n 0.0151209f $X=3.925 $Y=0.58 $X2=0
+ $Y2=0
cc_179 N_A_549_74#_c_209_n N_VGND_c_377_n 0.00573605f $X=2.885 $Y=0.58 $X2=0
+ $Y2=0
cc_180 N_A_549_74#_M1008_g N_VGND_c_379_n 0.0293656f $X=3.925 $Y=0.58 $X2=0
+ $Y2=0
cc_181 N_A_549_74#_c_209_n N_VGND_c_379_n 0.00594877f $X=2.885 $Y=0.58 $X2=0
+ $Y2=0
cc_182 N_A_682_74#_c_254_n N_VPWR_c_311_n 0.0163879f $X=4.72 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A_682_74#_c_262_n N_VPWR_c_311_n 0.0164467f $X=3.535 $Y=2.105 $X2=0
+ $Y2=0
cc_184 N_A_682_74#_c_256_n N_VPWR_c_311_n 0.0255637f $X=4.53 $Y=1.645 $X2=0
+ $Y2=0
cc_185 N_A_682_74#_c_262_n N_VPWR_c_314_n 0.0106198f $X=3.535 $Y=2.105 $X2=0
+ $Y2=0
cc_186 N_A_682_74#_c_254_n N_VPWR_c_315_n 0.00413917f $X=4.72 $Y=1.765 $X2=0
+ $Y2=0
cc_187 N_A_682_74#_c_254_n N_VPWR_c_308_n 0.00821389f $X=4.72 $Y=1.765 $X2=0
+ $Y2=0
cc_188 N_A_682_74#_c_262_n N_VPWR_c_308_n 0.00879013f $X=3.535 $Y=2.105 $X2=0
+ $Y2=0
cc_189 N_A_682_74#_M1003_g Y 8.21909e-19 $X=4.71 $Y=0.58 $X2=0 $Y2=0
cc_190 N_A_682_74#_M1003_g Y 0.0124475f $X=4.71 $Y=0.58 $X2=0 $Y2=0
cc_191 N_A_682_74#_c_254_n Y 0.0163621f $X=4.72 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A_682_74#_c_256_n Y 0.0140324f $X=4.53 $Y=1.645 $X2=0 $Y2=0
cc_193 N_A_682_74#_c_258_n Y 0.0133247f $X=4.53 $Y=0.965 $X2=0 $Y2=0
cc_194 N_A_682_74#_c_260_n Y 0.0384675f $X=4.67 $Y=1.46 $X2=0 $Y2=0
cc_195 N_A_682_74#_c_254_n Y 0.00229934f $X=4.72 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A_682_74#_M1003_g N_VGND_c_374_n 0.0112059f $X=4.71 $Y=0.58 $X2=0 $Y2=0
cc_197 N_A_682_74#_c_254_n N_VGND_c_374_n 3.24916e-19 $X=4.72 $Y=1.765 $X2=0
+ $Y2=0
cc_198 N_A_682_74#_c_255_n N_VGND_c_374_n 0.00743402f $X=3.535 $Y=0.565 $X2=0
+ $Y2=0
cc_199 N_A_682_74#_c_258_n N_VGND_c_374_n 0.0218411f $X=4.53 $Y=0.965 $X2=0
+ $Y2=0
cc_200 N_A_682_74#_c_255_n N_VGND_c_377_n 0.0108145f $X=3.535 $Y=0.565 $X2=0
+ $Y2=0
cc_201 N_A_682_74#_M1003_g N_VGND_c_378_n 0.00383152f $X=4.71 $Y=0.58 $X2=0
+ $Y2=0
cc_202 N_A_682_74#_M1003_g N_VGND_c_379_n 0.00761428f $X=4.71 $Y=0.58 $X2=0
+ $Y2=0
cc_203 N_A_682_74#_c_255_n N_VGND_c_379_n 0.0115915f $X=3.535 $Y=0.565 $X2=0
+ $Y2=0
cc_204 N_VPWR_c_311_n Y 0.0476994f $X=4.495 $Y=1.985 $X2=0 $Y2=0
cc_205 N_VPWR_c_315_n Y 0.0234396f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_206 N_VPWR_c_308_n Y 0.0138183f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_207 Y N_VGND_c_374_n 0.0124097f $X=4.95 $Y=0.47 $X2=0 $Y2=0
cc_208 Y N_VGND_c_378_n 0.0155069f $X=4.95 $Y=0.47 $X2=0 $Y2=0
cc_209 Y N_VGND_c_379_n 0.013122f $X=4.95 $Y=0.47 $X2=0 $Y2=0
