* File: sky130_fd_sc_ls__o22a_2.pex.spice
* Created: Fri Aug 28 13:48:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O22A_2%A_82_48# 1 2 9 11 13 16 18 20 24 26 27 28 29
+ 31 34 36 39 40 47
c92 39 0 8.46476e-20 $X=2.115 $Y=0.965
r93 46 47 15.5484 $w=3.41e-07 $l=1.1e-07 $layer=POLY_cond $X=0.915 $Y=1.532
+ $X2=1.025 $Y2=1.532
r94 45 46 48.0587 $w=3.41e-07 $l=3.4e-07 $layer=POLY_cond $X=0.575 $Y=1.532
+ $X2=0.915 $Y2=1.532
r95 39 40 4.54614 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=2.115 $Y=0.965
+ $X2=2.005 $Y2=0.965
r96 35 47 16.2551 $w=3.41e-07 $l=1.15e-07 $layer=POLY_cond $X=1.14 $Y=1.532
+ $X2=1.025 $Y2=1.532
r97 34 37 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.14 $Y=1.465
+ $X2=1.14 $Y2=1.63
r98 34 36 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.14 $Y=1.465
+ $X2=1.14 $Y2=1.3
r99 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.465 $X2=1.14 $Y2=1.465
r100 29 43 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=2.12
+ $X2=2.515 $Y2=2.035
r101 29 31 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=2.515 $Y=2.12
+ $X2=2.515 $Y2=2.775
r102 27 43 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=2.035
+ $X2=2.515 $Y2=2.035
r103 27 28 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=2.35 $Y=2.035
+ $X2=1.305 $Y2=2.035
r104 26 40 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=1.305 $Y=1.005
+ $X2=2.005 $Y2=1.005
r105 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.22 $Y=1.95
+ $X2=1.305 $Y2=2.035
r106 24 37 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.22 $Y=1.95
+ $X2=1.22 $Y2=1.63
r107 21 26 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.22 $Y=1.13
+ $X2=1.305 $Y2=1.005
r108 21 36 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.22 $Y=1.13
+ $X2=1.22 $Y2=1.3
r109 18 47 22.0049 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.025 $Y=1.765
+ $X2=1.025 $Y2=1.532
r110 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.025 $Y=1.765
+ $X2=1.025 $Y2=2.4
r111 14 46 22.0049 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.915 $Y=1.3
+ $X2=0.915 $Y2=1.532
r112 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.915 $Y=1.3
+ $X2=0.915 $Y2=0.74
r113 11 45 22.0049 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.575 $Y=1.765
+ $X2=0.575 $Y2=1.532
r114 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.575 $Y=1.765
+ $X2=0.575 $Y2=2.4
r115 7 45 12.7214 $w=3.41e-07 $l=9e-08 $layer=POLY_cond $X=0.485 $Y=1.532
+ $X2=0.575 $Y2=1.532
r116 7 9 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=0.485 $Y=1.39
+ $X2=0.485 $Y2=0.74
r117 2 43 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=2.365
+ $Y=1.92 $X2=2.515 $Y2=2.095
r118 2 31 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.365
+ $Y=1.92 $X2=2.515 $Y2=2.775
r119 1 39 182 $w=1.7e-07 $l=6.68019e-07 $layer=licon1_NDIFF $count=1 $X=1.96
+ $Y=0.37 $X2=2.115 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_2%B1 1 3 6 8
r33 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.595 $X2=1.71 $Y2=1.595
r34 4 11 38.9954 $w=3.66e-07 $l=2.21743e-07 $layer=POLY_cond $X=1.885 $Y=1.43
+ $X2=1.752 $Y2=1.595
r35 4 6 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.885 $Y=1.43
+ $X2=1.885 $Y2=0.74
r36 1 11 50.1894 $w=3.66e-07 $l=2.90689e-07 $layer=POLY_cond $X=1.84 $Y=1.845
+ $X2=1.752 $Y2=1.595
r37 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.84 $Y=1.845
+ $X2=1.84 $Y2=2.42
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_2%B2 1 3 6 8 12
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.335
+ $Y=1.595 $X2=2.335 $Y2=1.595
r34 8 12 5.76222 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=2.16 $Y=1.605
+ $X2=2.335 $Y2=1.605
r35 4 11 38.5562 $w=2.99e-07 $l=1.69926e-07 $layer=POLY_cond $X=2.345 $Y=1.43
+ $X2=2.335 $Y2=1.595
r36 4 6 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.345 $Y=1.43
+ $X2=2.345 $Y2=0.74
r37 1 11 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.29 $Y=1.845
+ $X2=2.335 $Y2=1.595
r38 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.29 $Y=1.845
+ $X2=2.29 $Y2=2.42
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_2%A2 1 3 6 8
c32 6 0 8.46476e-20 $X=2.845 $Y=0.74
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.875
+ $Y=1.595 $X2=2.875 $Y2=1.595
r34 8 12 8.0671 $w=3.48e-07 $l=2.45e-07 $layer=LI1_cond $X=3.12 $Y=1.605
+ $X2=2.875 $Y2=1.605
r35 4 11 38.5562 $w=2.99e-07 $l=1.79374e-07 $layer=POLY_cond $X=2.845 $Y=1.43
+ $X2=2.875 $Y2=1.595
r36 4 6 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.845 $Y=1.43
+ $X2=2.845 $Y2=0.74
r37 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.8 $Y=1.845
+ $X2=2.875 $Y2=1.595
r38 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.8 $Y=1.845 $X2=2.8
+ $Y2=2.42
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_2%A1 1 3 6 8 12
c24 6 0 7.64167e-20 $X=3.345 $Y=0.74
r25 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.465 $X2=3.57 $Y2=1.465
r26 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.57 $Y=1.665 $X2=3.57
+ $Y2=1.465
r27 4 11 38.9663 $w=3.64e-07 $l=2.26892e-07 $layer=POLY_cond $X=3.345 $Y=1.3
+ $X2=3.492 $Y2=1.465
r28 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.345 $Y=1.3 $X2=3.345
+ $Y2=0.74
r29 1 11 67.4361 $w=3.64e-07 $l=4.49622e-07 $layer=POLY_cond $X=3.34 $Y=1.845
+ $X2=3.492 $Y2=1.465
r30 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.34 $Y=1.845
+ $X2=3.34 $Y2=2.42
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_2%VPWR 1 2 3 10 12 16 20 22 24 28 30 42 48
r43 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r44 43 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 42 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 40 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 37 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r50 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 33 36 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r53 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 31 42 13.1831 $w=1.7e-07 $l=3.28e-07 $layer=LI1_cond $X=1.79 $Y=3.33
+ $X2=1.462 $Y2=3.33
r55 31 33 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.79 $Y=3.33 $X2=2.16
+ $Y2=3.33
r56 30 47 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=3.4 $Y=3.33 $X2=3.62
+ $Y2=3.33
r57 30 36 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.4 $Y=3.33 $X2=3.12
+ $Y2=3.33
r58 28 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 28 43 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 24 27 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.565 $Y=2.095
+ $X2=3.565 $Y2=2.775
r61 22 47 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=3.565 $Y=3.245
+ $X2=3.62 $Y2=3.33
r62 22 27 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=3.565 $Y=3.245
+ $X2=3.565 $Y2=2.775
r63 18 42 2.719 $w=6.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.462 $Y=3.245
+ $X2=1.462 $Y2=3.33
r64 18 20 15.2477 $w=6.53e-07 $l=8.35e-07 $layer=LI1_cond $X=1.462 $Y=3.245
+ $X2=1.462 $Y2=2.41
r65 17 39 4.68787 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.232 $Y2=3.33
r66 16 42 13.1831 $w=1.7e-07 $l=3.27e-07 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=1.462 $Y2=3.33
r67 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=0.465 $Y2=3.33
r68 12 15 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.3 $Y=1.985 $X2=0.3
+ $Y2=2.815
r69 10 39 3.0783 $w=3.3e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.3 $Y=3.245
+ $X2=0.232 $Y2=3.33
r70 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.3 $Y=3.245 $X2=0.3
+ $Y2=2.815
r71 3 27 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.415
+ $Y=1.92 $X2=3.565 $Y2=2.775
r72 3 24 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=3.415
+ $Y=1.92 $X2=3.565 $Y2=2.095
r73 2 20 150 $w=1.7e-07 $l=7.86416e-07 $layer=licon1_PDIFF $count=4 $X=1.1
+ $Y=1.84 $X2=1.615 $Y2=2.41
r74 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.84 $X2=0.3 $Y2=2.815
r75 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.84 $X2=0.3 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_2%X 1 2 9 15 17 19 20
r34 20 26 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.7 $Y=0.925
+ $X2=0.7 $Y2=1.13
r35 20 23 4.29215 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=0.7 $Y=0.925
+ $X2=0.7 $Y2=0.82
r36 19 26 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.72 $Y=1.82 $X2=0.72
+ $Y2=1.13
r37 15 19 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.8 $Y=1.985
+ $X2=0.8 $Y2=1.82
r38 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.8 $Y=1.985 $X2=0.8
+ $Y2=2.815
r39 9 23 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=0.662 $Y=0.515
+ $X2=0.662 $Y2=0.82
r40 2 17 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.84 $X2=0.8 $Y2=2.815
r41 2 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.84 $X2=0.8 $Y2=1.985
r42 1 20 182 $w=1.7e-07 $l=6.26099e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.37 $X2=0.7 $Y2=0.93
r43 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.37 $X2=0.7 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_2%VGND 1 2 3 10 12 16 20 22 24 29 39 40 46 49
r50 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r51 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r52 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r53 40 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r54 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=0 $X2=3.13
+ $Y2=0
r56 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.295 $Y=0 $X2=3.6
+ $Y2=0
r57 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r58 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r59 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r60 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r61 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r62 30 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.295 $Y=0 $X2=1.13
+ $Y2=0
r63 30 32 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.295 $Y=0 $X2=1.68
+ $Y2=0
r64 29 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=3.13
+ $Y2=0
r65 29 35 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=2.64
+ $Y2=0
r66 28 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r67 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r68 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r69 25 43 4.11164 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r70 25 27 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r71 24 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=1.13
+ $Y2=0
r72 24 27 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=0.72
+ $Y2=0
r73 22 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r74 22 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r75 18 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=0.085
+ $X2=3.13 $Y2=0
r76 18 20 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=3.13 $Y=0.085
+ $X2=3.13 $Y2=0.625
r77 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=0.085
+ $X2=1.13 $Y2=0
r78 14 16 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.13 $Y=0.085
+ $X2=1.13 $Y2=0.535
r79 10 43 3.10058 $w=2.6e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.235 $Y=0.085
+ $X2=0.182 $Y2=0
r80 10 12 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=0.235 $Y=0.085
+ $X2=0.235 $Y2=0.535
r81 3 20 182 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_NDIFF $count=1 $X=2.92
+ $Y=0.37 $X2=3.13 $Y2=0.625
r82 2 16 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.99
+ $Y=0.37 $X2=1.13 $Y2=0.535
r83 1 12 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.27 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_2%A_307_74# 1 2 3 10 12 13 14 15 18 20
c46 12 0 7.64167e-20 $X=2.63 $Y=0.52
r47 20 23 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.67 $Y=0.435
+ $X2=1.67 $Y2=0.57
r48 16 18 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=3.6 $Y=0.96 $X2=3.6
+ $Y2=0.515
r49 14 16 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.475 $Y=1.045
+ $X2=3.6 $Y2=0.96
r50 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.475 $Y=1.045
+ $X2=2.795 $Y2=1.045
r51 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.63 $Y=0.96
+ $X2=2.795 $Y2=1.045
r52 12 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=0.52 $X2=2.63
+ $Y2=0.435
r53 12 13 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.63 $Y=0.52
+ $X2=2.63 $Y2=0.96
r54 11 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=0.435
+ $X2=1.67 $Y2=0.435
r55 10 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0.435
+ $X2=2.63 $Y2=0.435
r56 10 11 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.465 $Y=0.435
+ $X2=1.835 $Y2=0.435
r57 3 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.42
+ $Y=0.37 $X2=3.56 $Y2=0.515
r58 2 26 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.42
+ $Y=0.37 $X2=2.63 $Y2=0.515
r59 1 23 182 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.37 $X2=1.67 $Y2=0.57
.ends

