* File: sky130_fd_sc_ls__o32ai_4.pex.spice
* Created: Wed Sep  2 11:23:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O32AI_4%B2 3 5 7 10 12 14 15 17 20 22 24 27 29 30 31
+ 32 52
c86 32 0 1.05621e-20 $X=1.68 $Y=1.665
c87 22 0 1.19081e-19 $X=1.855 $Y=1.765
r88 52 53 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=1.855 $Y=1.557
+ $X2=1.87 $Y2=1.557
r89 50 52 33.2189 $w=3.7e-07 $l=2.55e-07 $layer=POLY_cond $X=1.6 $Y=1.557
+ $X2=1.855 $Y2=1.557
r90 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.515 $X2=1.6 $Y2=1.515
r91 48 50 22.7973 $w=3.7e-07 $l=1.75e-07 $layer=POLY_cond $X=1.425 $Y=1.557
+ $X2=1.6 $Y2=1.557
r92 47 48 2.60541 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=1.405 $Y=1.557
+ $X2=1.425 $Y2=1.557
r93 46 51 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.26 $Y=1.605
+ $X2=1.6 $Y2=1.605
r94 45 47 18.8892 $w=3.7e-07 $l=1.45e-07 $layer=POLY_cond $X=1.26 $Y=1.557
+ $X2=1.405 $Y2=1.557
r95 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.26
+ $Y=1.515 $X2=1.26 $Y2=1.515
r96 43 45 39.7324 $w=3.7e-07 $l=3.05e-07 $layer=POLY_cond $X=0.955 $Y=1.557
+ $X2=1.26 $Y2=1.557
r97 42 43 3.90811 $w=3.7e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.557
+ $X2=0.955 $Y2=1.557
r98 40 42 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=0.92 $Y=1.557
+ $X2=0.925 $Y2=1.557
r99 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.92
+ $Y=1.515 $X2=0.92 $Y2=1.515
r100 38 40 54.0622 $w=3.7e-07 $l=4.15e-07 $layer=POLY_cond $X=0.505 $Y=1.557
+ $X2=0.92 $Y2=1.557
r101 37 38 1.3027 $w=3.7e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.505 $Y2=1.557
r102 32 51 2.63416 $w=3.48e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=1.605 $X2=1.6
+ $Y2=1.605
r103 31 46 1.97562 $w=3.48e-07 $l=6e-08 $layer=LI1_cond $X=1.2 $Y=1.605 $X2=1.26
+ $Y2=1.605
r104 31 41 9.21954 $w=3.48e-07 $l=2.8e-07 $layer=LI1_cond $X=1.2 $Y=1.605
+ $X2=0.92 $Y2=1.605
r105 30 41 6.58539 $w=3.48e-07 $l=2e-07 $layer=LI1_cond $X=0.72 $Y=1.605
+ $X2=0.92 $Y2=1.605
r106 29 30 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.605
+ $X2=0.72 $Y2=1.605
r107 25 53 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.87 $Y=1.35
+ $X2=1.87 $Y2=1.557
r108 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.87 $Y=1.35
+ $X2=1.87 $Y2=0.74
r109 22 52 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.557
r110 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r111 18 48 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=1.557
r112 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=0.74
r113 15 47 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.557
r114 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r115 12 43 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.557
r116 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r117 8 42 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=1.557
r118 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=0.74
r119 5 38 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.557
r120 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r121 1 37 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r122 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 33 56
c96 33 0 1.94211e-19 $X=4.08 $Y=1.665
c97 1 0 1.05621e-20 $X=2.305 $Y=1.765
r98 56 58 15.1863 $w=3.65e-07 $l=1.15e-07 $layer=POLY_cond $X=3.74 $Y=1.557
+ $X2=3.855 $Y2=1.557
r99 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.74
+ $Y=1.515 $X2=3.74 $Y2=1.515
r100 54 56 9.90411 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=3.665 $Y=1.557
+ $X2=3.74 $Y2=1.557
r101 52 54 34.9945 $w=3.65e-07 $l=2.65e-07 $layer=POLY_cond $X=3.4 $Y=1.557
+ $X2=3.665 $Y2=1.557
r102 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.4
+ $Y=1.515 $X2=3.4 $Y2=1.515
r103 50 52 5.94247 $w=3.65e-07 $l=4.5e-08 $layer=POLY_cond $X=3.355 $Y=1.557
+ $X2=3.4 $Y2=1.557
r104 49 50 19.8082 $w=3.65e-07 $l=1.5e-07 $layer=POLY_cond $X=3.205 $Y=1.557
+ $X2=3.355 $Y2=1.557
r105 47 49 19.1479 $w=3.65e-07 $l=1.45e-07 $layer=POLY_cond $X=3.06 $Y=1.557
+ $X2=3.205 $Y2=1.557
r106 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.06
+ $Y=1.515 $X2=3.06 $Y2=1.515
r107 45 47 27.0712 $w=3.65e-07 $l=2.05e-07 $layer=POLY_cond $X=2.855 $Y=1.557
+ $X2=3.06 $Y2=1.557
r108 44 45 13.2055 $w=3.65e-07 $l=1e-07 $layer=POLY_cond $X=2.755 $Y=1.557
+ $X2=2.855 $Y2=1.557
r109 43 48 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.72 $Y=1.605
+ $X2=3.06 $Y2=1.605
r110 42 44 4.62192 $w=3.65e-07 $l=3.5e-08 $layer=POLY_cond $X=2.72 $Y=1.557
+ $X2=2.755 $Y2=1.557
r111 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.72
+ $Y=1.515 $X2=2.72 $Y2=1.515
r112 40 42 48.2 $w=3.65e-07 $l=3.65e-07 $layer=POLY_cond $X=2.355 $Y=1.557
+ $X2=2.72 $Y2=1.557
r113 39 40 6.60274 $w=3.65e-07 $l=5e-08 $layer=POLY_cond $X=2.305 $Y=1.557
+ $X2=2.355 $Y2=1.557
r114 33 57 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=4.08 $Y=1.605
+ $X2=3.74 $Y2=1.605
r115 32 57 4.60977 $w=3.48e-07 $l=1.4e-07 $layer=LI1_cond $X=3.6 $Y=1.605
+ $X2=3.74 $Y2=1.605
r116 32 53 6.58539 $w=3.48e-07 $l=2e-07 $layer=LI1_cond $X=3.6 $Y=1.605 $X2=3.4
+ $Y2=1.605
r117 31 53 9.21954 $w=3.48e-07 $l=2.8e-07 $layer=LI1_cond $X=3.12 $Y=1.605
+ $X2=3.4 $Y2=1.605
r118 31 48 1.97562 $w=3.48e-07 $l=6e-08 $layer=LI1_cond $X=3.12 $Y=1.605
+ $X2=3.06 $Y2=1.605
r119 30 43 2.63416 $w=3.48e-07 $l=8e-08 $layer=LI1_cond $X=2.64 $Y=1.605
+ $X2=2.72 $Y2=1.605
r120 29 30 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.605
+ $X2=2.64 $Y2=1.605
r121 25 58 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.855 $Y=1.35
+ $X2=3.855 $Y2=1.557
r122 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.855 $Y=1.35
+ $X2=3.855 $Y2=0.74
r123 22 54 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.665 $Y=1.765
+ $X2=3.665 $Y2=1.557
r124 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.665 $Y=1.765
+ $X2=3.665 $Y2=2.4
r125 18 50 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.355 $Y=1.35
+ $X2=3.355 $Y2=1.557
r126 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.355 $Y=1.35
+ $X2=3.355 $Y2=0.74
r127 15 49 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.205 $Y=1.765
+ $X2=3.205 $Y2=1.557
r128 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.205 $Y=1.765
+ $X2=3.205 $Y2=2.4
r129 11 45 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.855 $Y=1.35
+ $X2=2.855 $Y2=1.557
r130 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.855 $Y=1.35
+ $X2=2.855 $Y2=0.74
r131 8 44 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=1.557
r132 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=2.4
r133 4 40 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.355 $Y=1.35
+ $X2=2.355 $Y2=1.557
r134 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.355 $Y=1.35
+ $X2=2.355 $Y2=0.74
r135 1 39 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.305 $Y2=1.557
r136 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.305 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_4%A3 3 5 6 7 9 12 14 16 19 21 23 26 28 30 31
+ 32 33 48
c95 28 0 1.24804e-19 $X=6.025 $Y=1.765
c96 7 0 2.43974e-19 $X=4.675 $Y=1.765
r97 48 49 20.6571 $w=3.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.875 $Y=1.557
+ $X2=6.025 $Y2=1.557
r98 47 48 41.3143 $w=3.5e-07 $l=3e-07 $layer=POLY_cond $X=5.575 $Y=1.557
+ $X2=5.875 $Y2=1.557
r99 46 47 18.5914 $w=3.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.44 $Y=1.557
+ $X2=5.575 $Y2=1.557
r100 44 46 1.37714 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=5.43 $Y=1.557
+ $X2=5.44 $Y2=1.557
r101 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.43
+ $Y=1.515 $X2=5.43 $Y2=1.515
r102 42 44 42.0029 $w=3.5e-07 $l=3.05e-07 $layer=POLY_cond $X=5.125 $Y=1.557
+ $X2=5.43 $Y2=1.557
r103 41 45 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=5.09 $Y=1.605
+ $X2=5.43 $Y2=1.605
r104 40 42 4.82 $w=3.5e-07 $l=3.5e-08 $layer=POLY_cond $X=5.09 $Y=1.557
+ $X2=5.125 $Y2=1.557
r105 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.09
+ $Y=1.515 $X2=5.09 $Y2=1.515
r106 38 40 19.9686 $w=3.5e-07 $l=1.45e-07 $layer=POLY_cond $X=4.945 $Y=1.557
+ $X2=5.09 $Y2=1.557
r107 37 38 37.1829 $w=3.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.675 $Y=1.557
+ $X2=4.945 $Y2=1.557
r108 33 45 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=5.52 $Y=1.605
+ $X2=5.43 $Y2=1.605
r109 32 41 1.64635 $w=3.48e-07 $l=5e-08 $layer=LI1_cond $X=5.04 $Y=1.605
+ $X2=5.09 $Y2=1.605
r110 31 32 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.605
+ $X2=5.04 $Y2=1.605
r111 28 49 22.6286 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.025 $Y=1.765
+ $X2=6.025 $Y2=1.557
r112 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.025 $Y=1.765
+ $X2=6.025 $Y2=2.4
r113 24 48 22.6286 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.875 $Y=1.35
+ $X2=5.875 $Y2=1.557
r114 24 26 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.875 $Y=1.35
+ $X2=5.875 $Y2=0.74
r115 21 47 22.6286 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.575 $Y=1.765
+ $X2=5.575 $Y2=1.557
r116 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.575 $Y=1.765
+ $X2=5.575 $Y2=2.4
r117 17 46 22.6286 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.44 $Y=1.35
+ $X2=5.44 $Y2=1.557
r118 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.44 $Y=1.35
+ $X2=5.44 $Y2=0.74
r119 14 42 22.6286 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.125 $Y=1.765
+ $X2=5.125 $Y2=1.557
r120 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.125 $Y=1.765
+ $X2=5.125 $Y2=2.4
r121 10 38 22.6286 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.945 $Y=1.35
+ $X2=4.945 $Y2=1.557
r122 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.945 $Y=1.35
+ $X2=4.945 $Y2=0.74
r123 7 37 22.6286 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.675 $Y=1.765
+ $X2=4.675 $Y2=1.557
r124 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.675 $Y=1.765
+ $X2=4.675 $Y2=2.4
r125 5 37 28.4554 $w=3.5e-07 $l=1.71184e-07 $layer=POLY_cond $X=4.585 $Y=1.425
+ $X2=4.675 $Y2=1.557
r126 5 6 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=4.585 $Y=1.425
+ $X2=4.43 $Y2=1.425
r127 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.355 $Y=1.35
+ $X2=4.43 $Y2=1.425
r128 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.355 $Y=1.35
+ $X2=4.355 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 33 50
c95 33 0 1.88749e-19 $X=8.4 $Y=1.665
c96 22 0 4.83678e-20 $X=8.025 $Y=1.765
r97 50 52 33.5655 $w=3.59e-07 $l=2.5e-07 $layer=POLY_cond $X=8.04 $Y=1.557
+ $X2=8.29 $Y2=1.557
r98 50 51 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=8.04
+ $Y=1.515 $X2=8.04 $Y2=1.515
r99 48 50 2.01393 $w=3.59e-07 $l=1.5e-08 $layer=POLY_cond $X=8.025 $Y=1.557
+ $X2=8.04 $Y2=1.557
r100 47 48 40.9499 $w=3.59e-07 $l=3.05e-07 $layer=POLY_cond $X=7.72 $Y=1.557
+ $X2=8.025 $Y2=1.557
r101 46 47 26.1811 $w=3.59e-07 $l=1.95e-07 $layer=POLY_cond $X=7.525 $Y=1.557
+ $X2=7.72 $Y2=1.557
r102 45 46 31.5515 $w=3.59e-07 $l=2.35e-07 $layer=POLY_cond $X=7.29 $Y=1.557
+ $X2=7.525 $Y2=1.557
r103 44 45 35.5794 $w=3.59e-07 $l=2.65e-07 $layer=POLY_cond $X=7.025 $Y=1.557
+ $X2=7.29 $Y2=1.557
r104 43 44 40.9499 $w=3.59e-07 $l=3.05e-07 $layer=POLY_cond $X=6.72 $Y=1.557
+ $X2=7.025 $Y2=1.557
r105 41 43 5.37047 $w=3.59e-07 $l=4e-08 $layer=POLY_cond $X=6.68 $Y=1.557
+ $X2=6.72 $Y2=1.557
r106 41 42 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.68
+ $Y=1.515 $X2=6.68 $Y2=1.515
r107 39 41 14.0975 $w=3.59e-07 $l=1.05e-07 $layer=POLY_cond $X=6.575 $Y=1.557
+ $X2=6.68 $Y2=1.557
r108 33 51 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.04 $Y2=1.565
r109 32 51 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=8.04 $Y2=1.565
r110 31 32 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.92 $Y2=1.565
r111 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r112 30 42 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.68 $Y2=1.565
r113 29 42 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=6.48 $Y=1.565 $X2=6.68
+ $Y2=1.565
r114 25 52 23.2387 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.29 $Y=1.35
+ $X2=8.29 $Y2=1.557
r115 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.29 $Y=1.35
+ $X2=8.29 $Y2=0.74
r116 22 48 23.2387 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.025 $Y=1.765
+ $X2=8.025 $Y2=1.557
r117 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.025 $Y=1.765
+ $X2=8.025 $Y2=2.4
r118 18 47 23.2387 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.72 $Y=1.35
+ $X2=7.72 $Y2=1.557
r119 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.72 $Y=1.35
+ $X2=7.72 $Y2=0.74
r120 15 46 23.2387 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.525 $Y=1.765
+ $X2=7.525 $Y2=1.557
r121 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.525 $Y=1.765
+ $X2=7.525 $Y2=2.4
r122 11 45 23.2387 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.29 $Y=1.35
+ $X2=7.29 $Y2=1.557
r123 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.29 $Y=1.35
+ $X2=7.29 $Y2=0.74
r124 8 44 23.2387 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.025 $Y=1.765
+ $X2=7.025 $Y2=1.557
r125 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.025 $Y=1.765
+ $X2=7.025 $Y2=2.4
r126 4 43 23.2387 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.72 $Y=1.35
+ $X2=6.72 $Y2=1.557
r127 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.72 $Y=1.35 $X2=6.72
+ $Y2=0.74
r128 1 39 23.2387 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.575 $Y=1.765
+ $X2=6.575 $Y2=1.557
r129 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.575 $Y=1.765
+ $X2=6.575 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_4%A1 3 5 7 10 12 14 17 19 21 24 26 28 29 30 31
+ 32 33 51
c81 33 0 4.83678e-20 $X=10.8 $Y=1.665
c82 5 0 6.39445e-20 $X=9.085 $Y=1.765
r83 51 52 46.0091 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=10.22 $Y=1.557
+ $X2=10.535 $Y2=1.557
r84 50 51 19.7182 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=10.085 $Y=1.557
+ $X2=10.22 $Y2=1.557
r85 48 50 19.7182 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=9.95 $Y=1.557
+ $X2=10.085 $Y2=1.557
r86 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.95
+ $Y=1.515 $X2=9.95 $Y2=1.515
r87 46 48 33.5939 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=9.72 $Y=1.557
+ $X2=9.95 $Y2=1.557
r88 45 46 27.0212 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=9.535 $Y=1.557
+ $X2=9.72 $Y2=1.557
r89 44 45 35.7848 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=9.29 $Y=1.557
+ $X2=9.535 $Y2=1.557
r90 42 44 2.92121 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=9.27 $Y=1.557 $X2=9.29
+ $Y2=1.557
r91 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.27
+ $Y=1.515 $X2=9.27 $Y2=1.515
r92 40 42 27.0212 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=9.085 $Y=1.557
+ $X2=9.27 $Y2=1.557
r93 39 40 43.0879 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=8.79 $Y=1.557
+ $X2=9.085 $Y2=1.557
r94 32 33 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=10.32 $Y=1.565
+ $X2=10.8 $Y2=1.565
r95 32 49 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.32 $Y=1.565
+ $X2=9.95 $Y2=1.565
r96 31 49 2.94811 $w=4.28e-07 $l=1.1e-07 $layer=LI1_cond $X=9.84 $Y=1.565
+ $X2=9.95 $Y2=1.565
r97 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.84 $Y2=1.565
r98 30 43 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=9.36 $Y=1.565 $X2=9.27
+ $Y2=1.565
r99 29 43 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.27 $Y2=1.565
r100 26 52 21.2229 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=10.535 $Y=1.765
+ $X2=10.535 $Y2=1.557
r101 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.535 $Y=1.765
+ $X2=10.535 $Y2=2.4
r102 22 51 21.2229 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.22 $Y=1.35
+ $X2=10.22 $Y2=1.557
r103 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.22 $Y=1.35
+ $X2=10.22 $Y2=0.74
r104 19 50 21.2229 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=10.085 $Y=1.765
+ $X2=10.085 $Y2=1.557
r105 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.085 $Y=1.765
+ $X2=10.085 $Y2=2.4
r106 15 46 21.2229 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.72 $Y=1.35
+ $X2=9.72 $Y2=1.557
r107 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.72 $Y=1.35
+ $X2=9.72 $Y2=0.74
r108 12 45 21.2229 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.535 $Y=1.765
+ $X2=9.535 $Y2=1.557
r109 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.535 $Y=1.765
+ $X2=9.535 $Y2=2.4
r110 8 44 21.2229 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.29 $Y=1.35
+ $X2=9.29 $Y2=1.557
r111 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.29 $Y=1.35
+ $X2=9.29 $Y2=0.74
r112 5 40 21.2229 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.085 $Y=1.765
+ $X2=9.085 $Y2=1.557
r113 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.085 $Y=1.765
+ $X2=9.085 $Y2=2.4
r114 1 39 21.2229 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.79 $Y=1.35
+ $X2=8.79 $Y2=1.557
r115 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.79 $Y=1.35 $X2=8.79
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_4%A_27_368# 1 2 3 4 5 18 22 23 26 28 30 31 32
+ 36 40 44 46
c74 46 0 1.68844e-19 $X=3.89 $Y=2.455
r75 37 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=2.375
+ $X2=2.98 $Y2=2.375
r76 36 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.725 $Y=2.375
+ $X2=3.89 $Y2=2.375
r77 36 37 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.725 $Y=2.375
+ $X2=3.145 $Y2=2.375
r78 33 42 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.245 $Y=2.375
+ $X2=2.12 $Y2=2.375
r79 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=2.375
+ $X2=2.98 $Y2=2.375
r80 32 33 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.815 $Y=2.375
+ $X2=2.245 $Y2=2.375
r81 30 42 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=2.46 $X2=2.12
+ $Y2=2.375
r82 30 31 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.12 $Y=2.46
+ $X2=2.12 $Y2=2.905
r83 29 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.265 $Y=2.99
+ $X2=1.14 $Y2=2.99
r84 28 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.995 $Y=2.99
+ $X2=2.12 $Y2=2.905
r85 28 29 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.995 $Y=2.99
+ $X2=1.265 $Y2=2.99
r86 24 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.905
+ $X2=1.14 $Y2=2.99
r87 24 26 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=1.14 $Y=2.905
+ $X2=1.14 $Y2=2.455
r88 22 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.015 $Y=2.99
+ $X2=1.14 $Y2=2.99
r89 22 23 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.015 $Y=2.99
+ $X2=0.445 $Y2=2.99
r90 18 21 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115 $X2=0.28
+ $Y2=2.815
r91 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r92 16 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905 $X2=0.28
+ $Y2=2.815
r93 5 46 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=3.74
+ $Y=1.84 $X2=3.89 $Y2=2.455
r94 4 44 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=2.83
+ $Y=1.84 $X2=2.98 $Y2=2.455
r95 3 42 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.455
r96 2 26 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.455
r97 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r98 1 18 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_4%Y 1 2 3 4 5 6 7 8 27 31 33 34 37 39 41 45 47
+ 51 53 57 62 64 67 68 69 70 72 74 75
r168 65 75 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.63 $Y=2.12
+ $X2=1.63 $Y2=2.405
r169 65 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=2.12
+ $X2=1.63 $Y2=2.035
r170 62 74 3.70735 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.89 $Y=1.95
+ $X2=5.805 $Y2=2.035
r171 61 62 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.89 $Y=1.26
+ $X2=5.89 $Y2=1.95
r172 58 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.065 $Y=2.035
+ $X2=4.9 $Y2=2.035
r173 57 74 2.76166 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.635 $Y=2.035
+ $X2=5.805 $Y2=2.035
r174 57 58 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.635 $Y=2.035
+ $X2=5.065 $Y2=2.035
r175 54 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.805 $Y=1.175
+ $X2=3.64 $Y2=1.175
r176 53 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.805 $Y=1.175
+ $X2=5.89 $Y2=1.26
r177 53 54 130.481 $w=1.68e-07 $l=2e-06 $layer=LI1_cond $X=5.805 $Y=1.175
+ $X2=3.805 $Y2=1.175
r178 49 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=1.09
+ $X2=3.64 $Y2=1.175
r179 49 51 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.64 $Y=1.09
+ $X2=3.64 $Y2=0.86
r180 48 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=1.175
+ $X2=2.64 $Y2=1.175
r181 47 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.475 $Y=1.175
+ $X2=3.64 $Y2=1.175
r182 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.475 $Y=1.175
+ $X2=2.805 $Y2=1.175
r183 43 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=1.09
+ $X2=2.64 $Y2=1.175
r184 43 45 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.64 $Y=1.09
+ $X2=2.64 $Y2=0.86
r185 42 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=1.175
+ $X2=1.68 $Y2=1.175
r186 41 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=1.175
+ $X2=2.64 $Y2=1.175
r187 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=1.175
+ $X2=1.805 $Y2=1.175
r188 40 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=2.035
+ $X2=1.63 $Y2=2.035
r189 39 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.735 $Y=2.035
+ $X2=4.9 $Y2=2.035
r190 39 40 191.807 $w=1.68e-07 $l=2.94e-06 $layer=LI1_cond $X=4.735 $Y=2.035
+ $X2=1.795 $Y2=2.035
r191 35 68 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=1.09
+ $X2=1.68 $Y2=1.175
r192 35 37 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=1.68 $Y=1.09
+ $X2=1.68 $Y2=0.86
r193 33 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.555 $Y=1.175
+ $X2=1.68 $Y2=1.175
r194 33 34 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.555 $Y=1.175
+ $X2=0.875 $Y2=1.175
r195 32 64 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=2.035
+ $X2=0.73 $Y2=2.035
r196 31 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=1.63 $Y2=2.035
r197 31 32 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=0.815 $Y2=2.035
r198 25 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.71 $Y=1.09
+ $X2=0.875 $Y2=1.175
r199 25 27 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.71 $Y=1.09
+ $X2=0.71 $Y2=0.86
r200 8 74 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=5.65
+ $Y=1.84 $X2=5.8 $Y2=2.115
r201 7 72 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=4.75
+ $Y=1.84 $X2=4.9 $Y2=2.115
r202 6 67 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.115
r203 5 64 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.115
r204 4 51 182 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=1 $X=3.43
+ $Y=0.37 $X2=3.64 $Y2=0.86
r205 3 45 182 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.37 $X2=2.64 $Y2=0.86
r206 2 37 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.86
r207 1 27 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_4%VPWR 1 2 3 4 5 18 22 26 30 32 34 39 40 42 43
+ 45 46 47 65 69 75 79
r121 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r122 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r123 73 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r124 73 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r125 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r126 70 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.975 $Y=3.33
+ $X2=9.81 $Y2=3.33
r127 70 72 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.975 $Y=3.33
+ $X2=10.32 $Y2=3.33
r128 69 78 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.675 $Y=3.33
+ $X2=10.857 $Y2=3.33
r129 69 72 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.675 $Y=3.33
+ $X2=10.32 $Y2=3.33
r130 68 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r131 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r132 65 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.645 $Y=3.33
+ $X2=9.81 $Y2=3.33
r133 65 67 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.645 $Y=3.33
+ $X2=9.36 $Y2=3.33
r134 64 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r135 63 64 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r136 60 63 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=8.4
+ $Y2=3.33
r137 60 61 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r138 58 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r139 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r140 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r141 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r142 51 55 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r143 50 54 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r144 50 51 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r145 47 64 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=8.4 $Y2=3.33
r146 47 61 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=3.6 $Y2=3.33
r147 45 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.695 $Y=3.33
+ $X2=8.4 $Y2=3.33
r148 45 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.695 $Y=3.33
+ $X2=8.82 $Y2=3.33
r149 44 67 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.945 $Y=3.33
+ $X2=9.36 $Y2=3.33
r150 44 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.945 $Y=3.33
+ $X2=8.82 $Y2=3.33
r151 42 57 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.345 $Y=3.33
+ $X2=3.12 $Y2=3.33
r152 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.345 $Y=3.33
+ $X2=3.43 $Y2=3.33
r153 41 60 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=3.33
+ $X2=3.6 $Y2=3.33
r154 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=3.33
+ $X2=3.43 $Y2=3.33
r155 39 54 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.16 $Y2=3.33
r156 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.53 $Y2=3.33
r157 38 57 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=3.12 $Y2=3.33
r158 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=2.53 $Y2=3.33
r159 34 37 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=10.8 $Y=2.115
+ $X2=10.8 $Y2=2.815
r160 32 78 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.8 $Y=3.245
+ $X2=10.857 $Y2=3.33
r161 32 37 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.8 $Y=3.245
+ $X2=10.8 $Y2=2.815
r162 28 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.81 $Y=3.245
+ $X2=9.81 $Y2=3.33
r163 28 30 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=9.81 $Y=3.245
+ $X2=9.81 $Y2=2.455
r164 24 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.82 $Y=3.245
+ $X2=8.82 $Y2=3.33
r165 24 26 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=8.82 $Y=3.245
+ $X2=8.82 $Y2=2.455
r166 20 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=3.33
r167 20 22 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=2.805
r168 16 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=3.245
+ $X2=2.53 $Y2=3.33
r169 16 18 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.53 $Y=3.245
+ $X2=2.53 $Y2=2.805
r170 5 37 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.61
+ $Y=1.84 $X2=10.76 $Y2=2.815
r171 5 34 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=10.61
+ $Y=1.84 $X2=10.76 $Y2=2.115
r172 4 30 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=9.61
+ $Y=1.84 $X2=9.81 $Y2=2.455
r173 3 26 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=8.715
+ $Y=1.84 $X2=8.86 $Y2=2.455
r174 2 22 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.84 $X2=3.43 $Y2=2.805
r175 1 18 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=1.84 $X2=2.53 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_4%A_861_368# 1 2 3 4 5 18 20 21 24 26 30 34 38
+ 40 44 46 47 48
r62 42 44 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.3 $Y=2.905 $X2=8.3
+ $Y2=2.455
r63 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.465 $Y=2.99
+ $X2=7.3 $Y2=2.99
r64 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.135 $Y=2.99
+ $X2=8.3 $Y2=2.905
r65 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.135 $Y=2.99
+ $X2=7.465 $Y2=2.99
r66 36 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.3 $Y=2.905 $X2=7.3
+ $Y2=2.99
r67 36 38 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.3 $Y=2.905 $X2=7.3
+ $Y2=2.455
r68 35 47 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.465 $Y=2.99
+ $X2=6.305 $Y2=2.99
r69 34 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.135 $Y=2.99
+ $X2=7.3 $Y2=2.99
r70 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.135 $Y=2.99
+ $X2=6.465 $Y2=2.99
r71 30 33 25.2097 $w=3.18e-07 $l=7e-07 $layer=LI1_cond $X=6.305 $Y=2.115
+ $X2=6.305 $Y2=2.815
r72 28 47 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.305 $Y=2.905
+ $X2=6.305 $Y2=2.99
r73 28 33 3.24125 $w=3.18e-07 $l=9e-08 $layer=LI1_cond $X=6.305 $Y=2.905
+ $X2=6.305 $Y2=2.815
r74 27 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.435 $Y=2.99
+ $X2=5.35 $Y2=2.99
r75 26 47 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.145 $Y=2.99
+ $X2=6.305 $Y2=2.99
r76 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=6.145 $Y=2.99
+ $X2=5.435 $Y2=2.99
r77 22 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.35 $Y=2.905
+ $X2=5.35 $Y2=2.99
r78 22 24 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.35 $Y=2.905
+ $X2=5.35 $Y2=2.455
r79 20 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.265 $Y=2.99
+ $X2=5.35 $Y2=2.99
r80 20 21 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.265 $Y=2.99
+ $X2=4.535 $Y2=2.99
r81 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.41 $Y=2.905
+ $X2=4.535 $Y2=2.99
r82 16 18 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=4.41 $Y=2.905
+ $X2=4.41 $Y2=2.455
r83 5 44 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=8.1
+ $Y=1.84 $X2=8.3 $Y2=2.455
r84 4 38 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=7.1
+ $Y=1.84 $X2=7.3 $Y2=2.455
r85 3 33 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=6.1
+ $Y=1.84 $X2=6.3 $Y2=2.815
r86 3 30 400 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=6.1
+ $Y=1.84 $X2=6.3 $Y2=2.115
r87 2 24 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=5.2
+ $Y=1.84 $X2=5.35 $Y2=2.455
r88 1 18 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=4.305
+ $Y=1.84 $X2=4.45 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_4%A_1330_368# 1 2 3 4 15 19 23 25 27 29 32 34
+ 36
r60 27 38 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.31 $Y=2.12
+ $X2=10.31 $Y2=2.035
r61 27 29 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=10.31 $Y=2.12
+ $X2=10.31 $Y2=2.815
r62 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.475 $Y=2.035
+ $X2=9.31 $Y2=2.035
r63 25 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.145 $Y=2.035
+ $X2=10.31 $Y2=2.035
r64 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.145 $Y=2.035
+ $X2=9.475 $Y2=2.035
r65 21 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.31 $Y=2.12 $X2=9.31
+ $Y2=2.035
r66 21 23 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=9.31 $Y=2.12
+ $X2=9.31 $Y2=2.815
r67 20 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.965 $Y=2.035
+ $X2=7.8 $Y2=2.035
r68 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.145 $Y=2.035
+ $X2=9.31 $Y2=2.035
r69 19 20 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=9.145 $Y=2.035
+ $X2=7.965 $Y2=2.035
r70 16 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.965 $Y=2.035
+ $X2=6.8 $Y2=2.035
r71 15 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.635 $Y=2.035
+ $X2=7.8 $Y2=2.035
r72 15 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.635 $Y=2.035
+ $X2=6.965 $Y2=2.035
r73 4 38 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=10.16
+ $Y=1.84 $X2=10.31 $Y2=2.115
r74 4 29 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.16
+ $Y=1.84 $X2=10.31 $Y2=2.815
r75 3 36 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=9.16
+ $Y=1.84 $X2=9.31 $Y2=2.115
r76 3 23 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.16
+ $Y=1.84 $X2=9.31 $Y2=2.815
r77 2 34 300 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=2 $X=7.6
+ $Y=1.84 $X2=7.8 $Y2=2.115
r78 1 32 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=6.65
+ $Y=1.84 $X2=6.8 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_4%A_27_74# 1 2 3 4 5 6 7 8 9 10 11 36 38 39 42
+ 44 48 50 54 56 61 62 63 66 68 70 74 76 80 82 86 88 92 94 95 96 98 102 104 105
+ 106
r184 102 103 4.15909 $w=5.72e-07 $l=1.95e-07 $layer=LI1_cond $X=6.332 $Y=0.9
+ $X2=6.332 $Y2=1.095
r185 100 102 1.38636 $w=5.72e-07 $l=6.5e-08 $layer=LI1_cond $X=6.332 $Y=0.835
+ $X2=6.332 $Y2=0.9
r186 90 92 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.505 $Y=1.01
+ $X2=10.505 $Y2=0.515
r187 89 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.67 $Y=1.095
+ $X2=9.505 $Y2=1.095
r188 88 90 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.34 $Y=1.095
+ $X2=10.505 $Y2=1.01
r189 88 89 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.34 $Y=1.095
+ $X2=9.67 $Y2=1.095
r190 84 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.505 $Y=1.01
+ $X2=9.505 $Y2=1.095
r191 84 86 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=9.505 $Y=1.01
+ $X2=9.505 $Y2=0.515
r192 83 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.67 $Y=1.095
+ $X2=8.505 $Y2=1.095
r193 82 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.34 $Y=1.095
+ $X2=9.505 $Y2=1.095
r194 82 83 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.34 $Y=1.095
+ $X2=8.67 $Y2=1.095
r195 78 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.505 $Y=1.01
+ $X2=8.505 $Y2=1.095
r196 78 80 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=8.505 $Y=1.01
+ $X2=8.505 $Y2=0.515
r197 77 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.67 $Y=1.095
+ $X2=7.505 $Y2=1.095
r198 76 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.34 $Y=1.095
+ $X2=8.505 $Y2=1.095
r199 76 77 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.34 $Y=1.095
+ $X2=7.67 $Y2=1.095
r200 72 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.505 $Y=1.01
+ $X2=7.505 $Y2=1.095
r201 72 74 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=7.505 $Y=1.01
+ $X2=7.505 $Y2=0.515
r202 71 103 8.0097 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=6.67 $Y=1.095
+ $X2=6.332 $Y2=1.095
r203 70 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.34 $Y=1.095
+ $X2=7.505 $Y2=1.095
r204 70 71 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.34 $Y=1.095
+ $X2=6.67 $Y2=1.095
r205 69 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.325 $Y=0.835
+ $X2=5.16 $Y2=0.835
r206 68 100 8.0097 $w=1.7e-07 $l=3.37e-07 $layer=LI1_cond $X=5.995 $Y=0.835
+ $X2=6.332 $Y2=0.835
r207 68 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.995 $Y=0.835
+ $X2=5.325 $Y2=0.835
r208 64 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.16 $Y=0.75
+ $X2=5.16 $Y2=0.835
r209 64 66 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.16 $Y=0.75
+ $X2=5.16 $Y2=0.495
r210 62 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.995 $Y=0.835
+ $X2=5.16 $Y2=0.835
r211 62 63 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.995 $Y=0.835
+ $X2=4.305 $Y2=0.835
r212 59 63 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.14 $Y=0.75
+ $X2=4.305 $Y2=0.835
r213 59 61 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.14 $Y=0.75
+ $X2=4.14 $Y2=0.635
r214 58 61 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=4.14 $Y=0.425
+ $X2=4.14 $Y2=0.635
r215 57 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=0.34
+ $X2=3.14 $Y2=0.34
r216 56 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.975 $Y=0.34
+ $X2=4.14 $Y2=0.425
r217 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.975 $Y=0.34
+ $X2=3.305 $Y2=0.34
r218 52 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=0.425
+ $X2=3.14 $Y2=0.34
r219 52 54 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.14 $Y=0.425
+ $X2=3.14 $Y2=0.635
r220 51 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0.34
+ $X2=2.14 $Y2=0.34
r221 50 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=0.34
+ $X2=3.14 $Y2=0.34
r222 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.975 $Y=0.34
+ $X2=2.305 $Y2=0.34
r223 46 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.425
+ $X2=2.14 $Y2=0.34
r224 46 48 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.14 $Y=0.425
+ $X2=2.14 $Y2=0.635
r225 45 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.34
+ $X2=1.21 $Y2=0.34
r226 44 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0.34
+ $X2=2.14 $Y2=0.34
r227 44 45 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.975 $Y=0.34
+ $X2=1.375 $Y2=0.34
r228 40 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.425
+ $X2=1.21 $Y2=0.34
r229 40 42 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.21 $Y=0.425
+ $X2=1.21 $Y2=0.635
r230 38 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=1.21 $Y2=0.34
r231 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=0.365 $Y2=0.34
r232 34 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.425
+ $X2=0.365 $Y2=0.34
r233 34 36 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.24 $Y=0.425
+ $X2=0.24 $Y2=0.515
r234 11 92 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=10.295
+ $Y=0.37 $X2=10.505 $Y2=0.515
r235 10 86 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.365
+ $Y=0.37 $X2=9.505 $Y2=0.515
r236 9 80 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.365
+ $Y=0.37 $X2=8.505 $Y2=0.515
r237 8 74 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.365
+ $Y=0.37 $X2=7.505 $Y2=0.515
r238 7 102 121.333 $w=1.7e-07 $l=7.75999e-07 $layer=licon1_NDIFF $count=1
+ $X=5.95 $Y=0.37 $X2=6.505 $Y2=0.9
r239 7 100 121.333 $w=1.7e-07 $l=5.60245e-07 $layer=licon1_NDIFF $count=1
+ $X=5.95 $Y=0.37 $X2=6.16 $Y2=0.835
r240 6 98 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=5.02
+ $Y=0.37 $X2=5.16 $Y2=0.835
r241 6 66 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.02
+ $Y=0.37 $X2=5.16 $Y2=0.495
r242 5 61 182 $w=1.7e-07 $l=3.54789e-07 $layer=licon1_NDIFF $count=1 $X=3.93
+ $Y=0.37 $X2=4.14 $Y2=0.635
r243 4 54 182 $w=1.7e-07 $l=3.54789e-07 $layer=licon1_NDIFF $count=1 $X=2.93
+ $Y=0.37 $X2=3.14 $Y2=0.635
r244 3 48 182 $w=1.7e-07 $l=3.49142e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.37 $X2=2.14 $Y2=0.635
r245 2 42 182 $w=1.7e-07 $l=3.54789e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.37 $X2=1.21 $Y2=0.635
r246 1 36 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O32AI_4%VGND 1 2 3 4 5 6 21 23 27 31 33 37 39 43 45
+ 49 51 53 58 65 66 69 72 75 78 81 84
r134 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r135 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r136 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r137 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r138 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r139 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r140 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r141 69 70 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r142 66 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0 $X2=9.84
+ $Y2=0
r143 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r144 63 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.17 $Y=0
+ $X2=10.005 $Y2=0
r145 63 65 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=10.17 $Y=0 $X2=10.8
+ $Y2=0
r146 62 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r147 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r148 59 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.825 $Y=0 $X2=5.66
+ $Y2=0
r149 59 61 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.825 $Y=0
+ $X2=6.48 $Y2=0
r150 58 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.84 $Y=0 $X2=7.005
+ $Y2=0
r151 58 61 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.84 $Y=0 $X2=6.48
+ $Y2=0
r152 56 70 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=4.56
+ $Y2=0
r153 55 56 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r154 53 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.485 $Y=0 $X2=4.65
+ $Y2=0
r155 53 55 276.947 $w=1.68e-07 $l=4.245e-06 $layer=LI1_cond $X=4.485 $Y=0
+ $X2=0.24 $Y2=0
r156 51 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r157 51 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r158 51 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r159 47 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.005 $Y=0.085
+ $X2=10.005 $Y2=0
r160 47 49 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=10.005 $Y=0.085
+ $X2=10.005 $Y2=0.595
r161 46 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.17 $Y=0 $X2=9.005
+ $Y2=0
r162 45 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.84 $Y=0
+ $X2=10.005 $Y2=0
r163 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.84 $Y=0 $X2=9.17
+ $Y2=0
r164 41 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.005 $Y=0.085
+ $X2=9.005 $Y2=0
r165 41 43 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=9.005 $Y=0.085
+ $X2=9.005 $Y2=0.595
r166 40 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.17 $Y=0 $X2=8.005
+ $Y2=0
r167 39 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.84 $Y=0 $X2=9.005
+ $Y2=0
r168 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.84 $Y=0 $X2=8.17
+ $Y2=0
r169 35 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.005 $Y=0.085
+ $X2=8.005 $Y2=0
r170 35 37 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=8.005 $Y=0.085
+ $X2=8.005 $Y2=0.595
r171 34 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.17 $Y=0 $X2=7.005
+ $Y2=0
r172 33 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.84 $Y=0 $X2=8.005
+ $Y2=0
r173 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.84 $Y=0 $X2=7.17
+ $Y2=0
r174 29 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.005 $Y=0.085
+ $X2=7.005 $Y2=0
r175 29 31 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=7.005 $Y=0.085
+ $X2=7.005 $Y2=0.595
r176 25 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.66 $Y=0.085
+ $X2=5.66 $Y2=0
r177 25 27 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.66 $Y=0.085
+ $X2=5.66 $Y2=0.495
r178 24 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=0 $X2=4.65
+ $Y2=0
r179 23 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.495 $Y=0 $X2=5.66
+ $Y2=0
r180 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.495 $Y=0
+ $X2=4.815 $Y2=0
r181 19 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=0.085
+ $X2=4.65 $Y2=0
r182 19 21 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=4.65 $Y=0.085
+ $X2=4.65 $Y2=0.415
r183 6 49 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=9.795
+ $Y=0.37 $X2=10.005 $Y2=0.595
r184 5 43 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=8.865
+ $Y=0.37 $X2=9.005 $Y2=0.595
r185 4 37 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=7.795
+ $Y=0.37 $X2=8.005 $Y2=0.595
r186 3 31 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=6.795
+ $Y=0.37 $X2=7.005 $Y2=0.595
r187 2 27 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.515
+ $Y=0.37 $X2=5.66 $Y2=0.495
r188 1 21 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.37 $X2=4.65 $Y2=0.415
.ends

