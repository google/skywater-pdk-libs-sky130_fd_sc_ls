* NGSPICE file created from sky130_fd_sc_ls__a2111o_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 a_137_260# D1 a_549_392# VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=8.5e+11p ps=7.7e+06u
M1001 VGND a_137_260# X VNB nshort w=740000u l=150000u
+  ad=1.3711e+12p pd=1.359e+07u as=4.144e+11p ps=4.08e+06u
M1002 a_814_392# C1 a_549_392# VPB phighvt w=1e+06u l=150000u
+  ad=6e+11p pd=5.2e+06u as=0p ps=0u
M1003 VGND C1 a_137_260# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=7.168e+11p ps=7.36e+06u
M1004 VPWR A2 a_1013_392# VPB phighvt w=1e+06u l=150000u
+  ad=1.552e+12p pd=1.362e+07u as=1.15e+12p ps=1.03e+07u
M1005 X a_137_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1006 a_1210_74# A2 VGND VNB nshort w=640000u l=150000u
+  ad=5.184e+11p pd=5.46e+06u as=0p ps=0u
M1007 a_814_392# B1 a_1013_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B1 a_137_260# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_549_392# C1 a_814_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1013_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_137_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_137_260# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_137_260# D1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1013_392# B1 a_814_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1210_74# A1 a_137_260# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_137_260# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A1 a_1013_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_137_260# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND D1 a_137_260# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_137_260# C1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_137_260# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_137_260# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_549_392# D1 a_137_260# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_137_260# B1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A2 a_1210_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1013_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_137_260# A1 a_1210_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

