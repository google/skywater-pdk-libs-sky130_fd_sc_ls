* File: sky130_fd_sc_ls__or4bb_1.spice
* Created: Fri Aug 28 14:00:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__or4bb_1.pex.spice"
.subckt sky130_fd_sc_ls__or4bb_1  VNB VPB C_N D_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* D_N	D_N
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_C_N_M1003_g N_A_27_424#_M1003_s VNB NSHORT L=0.15 W=0.55
+ AD=0.1155 AS=0.15675 PD=0.97 PS=1.67 NRD=15.264 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1004 N_A_216_424#_M1004_d N_D_N_M1004_g N_VGND_M1003_d VNB NSHORT L=0.15
+ W=0.55 AD=0.15675 AS=0.1155 PD=1.67 PS=0.97 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75000.8 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1001 N_A_357_378#_M1001_d N_A_216_424#_M1001_g N_VGND_M1001_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.092125 AS=0.165 PD=0.885 PS=1.7 NRD=11.988 NRS=3.264 M=1
+ R=3.66667 SA=75000.2 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1013 N_VGND_M1013_d N_A_27_424#_M1013_g N_A_357_378#_M1001_d VNB NSHORT L=0.15
+ W=0.55 AD=0.114125 AS=0.092125 PD=0.965 PS=0.885 NRD=21.816 NRS=0 M=1
+ R=3.66667 SA=75000.7 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1009 N_A_357_378#_M1009_d N_B_M1009_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.55
+ AD=0.09625 AS=0.114125 PD=0.9 PS=0.965 NRD=15.264 NRS=7.632 M=1 R=3.66667
+ SA=75001.3 SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_357_378#_M1009_d VNB NSHORT L=0.15 W=0.55
+ AD=0.126948 AS=0.09625 PD=1.01899 PS=0.9 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75001.8 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1010 N_X_M1010_d N_A_357_378#_M1010_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.170802 PD=2.05 PS=1.37101 NRD=0 NRS=17.016 M=1 R=4.93333
+ SA=75001.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_C_N_M1008_g N_A_27_424#_M1008_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.147 AS=0.2478 PD=1.19 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1006 N_A_216_424#_M1006_d N_D_N_M1006_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.43785 AS=0.147 PD=2.97 PS=1.19 NRD=109.335 NRS=0 M=1 R=5.6
+ SA=75000.7 SB=75000.4 A=0.126 P=1.98 MULT=1
MM1000 A_446_378# N_A_216_424#_M1000_g N_A_357_378#_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1011 A_530_378# N_A_27_424#_M1011_g A_446_378# VPB PHIGHVT L=0.15 W=1 AD=0.165
+ AS=0.135 PD=1.33 PS=1.27 NRD=21.6503 NRS=15.7403 M=1 R=6.66667 SA=75000.6
+ SB=75001.8 A=0.15 P=2.3 MULT=1
MM1002 A_626_378# N_B_M1002_g A_530_378# VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.165 PD=1.39 PS=1.33 NRD=27.5603 NRS=21.6503 M=1 R=6.66667 SA=75001.1
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1012_d N_A_M1012_g A_626_378# VPB PHIGHVT L=0.15 W=1 AD=0.22283
+ AS=0.195 PD=1.46698 PS=1.39 NRD=19.0302 NRS=27.5603 M=1 R=6.66667 SA=75001.7
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1007 N_X_M1007_d N_A_357_378#_M1007_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.24957 PD=2.83 PS=1.64302 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002 SB=75000.2 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ls__or4bb_1.pxi.spice"
*
.ends
*
*
