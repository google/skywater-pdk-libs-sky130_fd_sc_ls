* File: sky130_fd_sc_ls__nand4bb_1.spice
* Created: Fri Aug 28 13:35:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nand4bb_1.pex.spice"
.subckt sky130_fd_sc_ls__nand4bb_1  VNB VPB A_N B_N C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B_N	B_N
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_N_M1002_g N_A_27_398#_M1002_s VNB NSHORT L=0.15 W=0.55
+ AD=0.122187 AS=0.150975 PD=1.025 PS=1.67 NRD=17.448 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1000 N_A_226_398#_M1000_d N_B_N_M1000_g N_VGND_M1002_d VNB NSHORT L=0.15
+ W=0.55 AD=0.15055 AS=0.122187 PD=1.69 PS=1.025 NRD=1.08 NRS=15.264 M=1
+ R=3.66667 SA=75000.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1005 A_435_74# N_A_27_398#_M1005_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.0888 AS=0.19585 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1001 A_513_74# N_A_226_398#_M1001_g A_435_74# VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333
+ SA=75000.6 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1010 A_627_74# N_C_M1010_g A_513_74# VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.1554 PD=1.16 PS=1.16 NRD=25.128 NRS=25.128 M=1 R=4.93333 SA=75001.1
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_D_M1003_g A_627_74# VNB NSHORT L=0.15 W=0.74 AD=0.266
+ AS=0.1554 PD=2.34 PS=1.16 NRD=23.508 NRS=25.128 M=1 R=4.93333 SA=75001.7
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1009 N_VPWR_M1009_d N_A_N_M1009_g N_A_27_398#_M1009_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.168 AS=0.2478 PD=1.24 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1007 N_A_226_398#_M1007_d N_B_N_M1007_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.168 PD=2.27 PS=1.24 NRD=2.3443 NRS=14.0658 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_VPWR_M1008_d N_A_27_398#_M1008_g N_Y_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.2464 AS=0.3304 PD=1.56 PS=2.83 NRD=18.4589 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1004_d N_A_226_398#_M1004_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.2464 PD=1.47 PS=1.56 NRD=10.5395 NRS=9.6727 M=1 R=7.46667
+ SA=75000.8 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_C_M1006_g N_Y_M1004_d VPB PHIGHVT L=0.15 W=1.12 AD=0.224
+ AS=0.196 PD=1.52 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75001.3
+ SB=75000.8 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1011_d N_D_M1011_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.224 PD=2.83 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.9 SB=75000.2 A=0.168 P=2.54 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__nand4bb_1.pxi.spice"
*
.ends
*
*
