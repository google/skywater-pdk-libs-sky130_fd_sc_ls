* File: sky130_fd_sc_ls__sdfbbp_1.pex.spice
* Created: Wed Sep  2 11:26:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%SCD 2 3 5 8 9 10 14 15 16
r28 18 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.97 $X2=0.385 $Y2=1.97
r29 14 16 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.29
+ $X2=0.407 $Y2=1.125
r30 14 15 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.29 $X2=0.385 $Y2=1.29
r31 10 19 8.27047 $w=4.23e-07 $l=3.05e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.97
r32 9 10 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.665
r33 9 15 0.135582 $w=4.23e-07 $l=5e-09 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.29
r34 8 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.52 $Y=0.805
+ $X2=0.52 $Y2=1.125
r35 3 18 56.1009 $w=3.02e-07 $l=3.20273e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.407 $Y2=1.97
r36 3 5 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.64
r37 2 18 4.79453 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.407 $Y=1.948
+ $X2=0.407 $Y2=1.97
r38 1 14 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.407 $Y=1.312
+ $X2=0.407 $Y2=1.29
r39 1 2 94.3237 $w=3.75e-07 $l=6.36e-07 $layer=POLY_cond $X=0.407 $Y=1.312
+ $X2=0.407 $Y2=1.948
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%D 3 6 7 9 10 16
c45 10 0 1.39381e-19 $X=1.68 $Y=1.665
r46 14 16 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=1.435 $Y=1.69
+ $X2=1.61 $Y2=1.69
r47 12 14 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.42 $Y=1.69
+ $X2=1.435 $Y2=1.69
r48 10 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.69 $X2=1.61 $Y2=1.69
r49 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.435 $Y=2.245
+ $X2=1.435 $Y2=2.64
r50 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.435 $Y=2.155 $X2=1.435
+ $Y2=2.245
r51 5 14 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.855
+ $X2=1.435 $Y2=1.69
r52 5 6 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=1.435 $Y=1.855 $X2=1.435
+ $Y2=2.155
r53 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.525
+ $X2=1.42 $Y2=1.69
r54 1 3 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.42 $Y=1.525 $X2=1.42
+ $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%A_341_93# 1 2 9 11 13 14 15 17 22 26 30 33
+ 34 35 38
c82 15 0 6.84835e-20 $X=1.855 $Y=1.24
r83 35 38 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=2.695 $Y=1.83
+ $X2=2.695 $Y2=1.035
r84 33 36 6.39487 $w=5.03e-07 $l=2.7e-07 $layer=LI1_cond $X=2.527 $Y=1.995
+ $X2=2.527 $Y2=2.265
r85 33 35 9.54788 $w=5.03e-07 $l=1.65e-07 $layer=LI1_cond $X=2.527 $Y=1.995
+ $X2=2.527 $Y2=1.83
r86 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.43
+ $Y=1.995 $X2=2.43 $Y2=1.995
r87 28 30 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=2.35
+ $X2=3.12 $Y2=2.465
r88 27 36 7.21919 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=2.78 $Y=2.265
+ $X2=2.527 $Y2=2.265
r89 26 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.955 $Y=2.265
+ $X2=3.12 $Y2=2.35
r90 26 27 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.955 $Y=2.265
+ $X2=2.78 $Y2=2.265
r91 20 38 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.735 $Y=0.91
+ $X2=2.735 $Y2=1.035
r92 20 22 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=2.735 $Y=0.91
+ $X2=2.735 $Y2=0.815
r93 19 34 35.5134 $w=4.15e-07 $l=2.65e-07 $layer=POLY_cond $X=2.165 $Y=2.037
+ $X2=2.43 $Y2=2.037
r94 17 19 49.3036 $w=2.29e-07 $l=2.41607e-07 $layer=POLY_cond $X=2.09 $Y=1.83
+ $X2=2.015 $Y2=2.037
r95 16 17 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=2.09 $Y=1.315
+ $X2=2.09 $Y2=1.83
r96 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.015 $Y=1.24
+ $X2=2.09 $Y2=1.315
r97 14 15 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.015 $Y=1.24
+ $X2=1.855 $Y2=1.24
r98 11 19 49.5141 $w=2.29e-07 $l=2.65149e-07 $layer=POLY_cond $X=1.885 $Y=2.245
+ $X2=2.015 $Y2=2.037
r99 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.885 $Y=2.245
+ $X2=1.885 $Y2=2.64
r100 7 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.78 $Y=1.165
+ $X2=1.855 $Y2=1.24
r101 7 9 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.78 $Y=1.165
+ $X2=1.78 $Y2=0.805
r102 2 30 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.97
+ $Y=2.32 $X2=3.12 $Y2=2.465
r103 1 22 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.595 $X2=2.695 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%SCE 4 5 7 8 9 13 14 15 17 18 20 21
c84 5 0 7.0898e-20 $X=1.015 $Y=2.245
r85 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.93 $X2=0.97 $Y2=1.93
r86 21 25 6.60335 $w=4.78e-07 $l=2.65e-07 $layer=LI1_cond $X=1.045 $Y=1.665
+ $X2=1.045 $Y2=1.93
r87 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.895 $Y=2.245
+ $X2=2.895 $Y2=2.64
r88 17 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.895 $Y=2.155
+ $X2=2.895 $Y2=2.245
r89 16 17 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=2.895 $Y=1.455
+ $X2=2.895 $Y2=2.155
r90 14 16 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.805 $Y=1.38
+ $X2=2.895 $Y2=1.455
r91 14 15 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.805 $Y=1.38
+ $X2=2.555 $Y2=1.38
r92 11 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.48 $Y=1.305
+ $X2=2.555 $Y2=1.38
r93 11 13 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.48 $Y=1.305 $X2=2.48
+ $Y2=0.805
r94 10 13 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.48 $Y=0.255
+ $X2=2.48 $Y2=0.805
r95 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.405 $Y=0.18
+ $X2=2.48 $Y2=0.255
r96 8 9 728.128 $w=1.5e-07 $l=1.42e-06 $layer=POLY_cond $X=2.405 $Y=0.18
+ $X2=0.985 $Y2=0.18
r97 5 24 64.2376 $w=2.83e-07 $l=3.36749e-07 $layer=POLY_cond $X=1.015 $Y=2.245
+ $X2=0.97 $Y2=1.93
r98 5 7 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.015 $Y=2.245
+ $X2=1.015 $Y2=2.64
r99 2 24 38.6899 $w=2.83e-07 $l=1.92678e-07 $layer=POLY_cond $X=0.91 $Y=1.765
+ $X2=0.97 $Y2=1.93
r100 2 4 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=0.91 $Y=1.765
+ $X2=0.91 $Y2=0.805
r101 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.91 $Y=0.255
+ $X2=0.985 $Y2=0.18
r102 1 4 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.91 $Y=0.255
+ $X2=0.91 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%CLK 1 3 4 6 7 11
r44 11 13 42.8138 $w=3.49e-07 $l=3.1e-07 $layer=POLY_cond $X=3.595 $Y=1.552
+ $X2=3.905 $Y2=1.552
r45 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.595
+ $Y=1.505 $X2=3.595 $Y2=1.505
r46 9 11 17.2636 $w=3.49e-07 $l=1.25e-07 $layer=POLY_cond $X=3.47 $Y=1.552
+ $X2=3.595 $Y2=1.552
r47 7 12 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.595 $Y=1.295
+ $X2=3.595 $Y2=1.505
r48 4 13 22.56 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=3.905 $Y=1.765
+ $X2=3.905 $Y2=1.552
r49 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.905 $Y=1.765
+ $X2=3.905 $Y2=2.4
r50 1 9 22.56 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=3.47 $Y=1.34 $X2=3.47
+ $Y2=1.552
r51 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.47 $Y=1.34 $X2=3.47
+ $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%A_1250_231# 1 2 9 11 12 14 15 17 18 20 22
+ 25 26 29 32 34 35 36 41 43 47 48 49 51
c159 43 0 2.56036e-20 $X=8.85 $Y=1.5
c160 41 0 2.04581e-20 $X=8.85 $Y=1.825
c161 29 0 1.67029e-19 $X=6.535 $Y=0.815
c162 18 0 3.40541e-20 $X=9.25 $Y=1.295
c163 15 0 1.14272e-19 $X=8.755 $Y=1.82
r164 46 48 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=7.985 $Y=0.777
+ $X2=8.15 $Y2=0.777
r165 46 47 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=7.985 $Y=0.777
+ $X2=7.82 $Y2=0.777
r166 44 53 32.2908 $w=3.06e-07 $l=2.05e-07 $layer=POLY_cond $X=8.84 $Y=1.5
+ $X2=8.84 $Y2=1.295
r167 43 49 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.85 $Y=1.5
+ $X2=8.85 $Y2=1.335
r168 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.85
+ $Y=1.5 $X2=8.85 $Y2=1.5
r169 41 43 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=8.85 $Y=1.825
+ $X2=8.85 $Y2=1.5
r170 38 49 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=8.77 $Y=0.9
+ $X2=8.77 $Y2=1.335
r171 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.685 $Y=0.815
+ $X2=8.77 $Y2=0.9
r172 36 48 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=8.685 $Y=0.815
+ $X2=8.15 $Y2=0.815
r173 34 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.685 $Y=1.91
+ $X2=8.85 $Y2=1.825
r174 34 35 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.685 $Y=1.91
+ $X2=7.765 $Y2=1.91
r175 30 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.6 $Y=1.995
+ $X2=7.765 $Y2=1.91
r176 30 32 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=7.6 $Y=1.995
+ $X2=7.6 $Y2=2.04
r177 29 47 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=6.535 $Y=0.815
+ $X2=7.82 $Y2=0.815
r178 26 52 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.415 $Y=1.32
+ $X2=6.415 $Y2=1.485
r179 26 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.415 $Y=1.32
+ $X2=6.415 $Y2=1.155
r180 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.415
+ $Y=1.32 $X2=6.415 $Y2=1.32
r181 23 29 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=6.415 $Y=0.9
+ $X2=6.535 $Y2=0.815
r182 23 25 20.1678 $w=2.38e-07 $l=4.2e-07 $layer=LI1_cond $X=6.415 $Y=0.9
+ $X2=6.415 $Y2=1.32
r183 20 22 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.325 $Y=1.22
+ $X2=9.325 $Y2=0.87
r184 19 53 19.4347 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=9.015 $Y=1.295
+ $X2=8.84 $Y2=1.295
r185 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.25 $Y=1.295
+ $X2=9.325 $Y2=1.22
r186 18 19 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=9.25 $Y=1.295
+ $X2=9.015 $Y2=1.295
r187 15 44 62.95 $w=3.06e-07 $l=3.6e-07 $layer=POLY_cond $X=8.755 $Y=1.82
+ $X2=8.84 $Y2=1.5
r188 15 17 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.755 $Y=1.82
+ $X2=8.755 $Y2=2.315
r189 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.45 $Y=2.02
+ $X2=6.45 $Y2=2.305
r190 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.45 $Y=1.93 $X2=6.45
+ $Y2=2.02
r191 11 52 172.976 $w=1.8e-07 $l=4.45e-07 $layer=POLY_cond $X=6.45 $Y=1.93
+ $X2=6.45 $Y2=1.485
r192 9 51 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.36 $Y=0.835
+ $X2=6.36 $Y2=1.155
r193 2 32 300 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=2 $X=7.36
+ $Y=1.895 $X2=7.6 $Y2=2.04
r194 1 46 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=7.845
+ $Y=0.595 $X2=7.985 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%SET_B 3 5 7 10 12 14 16 17 18 20 21 22 24
+ 25 26 28 31 32 34 38 39 40
c169 26 0 9.6863e-20 $X=9.025 $Y=2.99
r170 45 47 5.37107 $w=3.18e-07 $l=1.4e-07 $layer=LI1_cond $X=11.22 $Y=1.635
+ $X2=11.22 $Y2=1.775
r171 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.22
+ $Y=1.635 $X2=11.22 $Y2=1.635
r172 40 47 9.97484 $w=3.18e-07 $l=2.6e-07 $layer=LI1_cond $X=11.22 $Y=2.035
+ $X2=11.22 $Y2=1.775
r173 38 39 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=10.195 $Y=2.015
+ $X2=10.195 $Y2=2.185
r174 34 37 6.89066 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=7.21 $Y=1.535
+ $X2=7.21 $Y2=1.655
r175 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.21
+ $Y=1.535 $X2=7.21 $Y2=1.535
r176 31 47 4.40442 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.055 $Y=1.775
+ $X2=11.22 $Y2=1.775
r177 31 32 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=11.055 $Y=1.775
+ $X2=10.295 $Y2=1.775
r178 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.21 $Y=1.86
+ $X2=10.295 $Y2=1.775
r179 29 38 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=10.21 $Y=1.86
+ $X2=10.21 $Y2=2.015
r180 28 39 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=10.18 $Y=2.905
+ $X2=10.18 $Y2=2.185
r181 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.095 $Y=2.99
+ $X2=10.18 $Y2=2.905
r182 25 26 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=10.095 $Y=2.99
+ $X2=9.025 $Y2=2.99
r183 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.94 $Y=2.905
+ $X2=9.025 $Y2=2.99
r184 23 24 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.94 $Y=2.335
+ $X2=8.94 $Y2=2.905
r185 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.855 $Y=2.25
+ $X2=8.94 $Y2=2.335
r186 21 22 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=8.855 $Y=2.25
+ $X2=8.105 $Y2=2.25
r187 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.02 $Y=2.335
+ $X2=8.105 $Y2=2.25
r188 19 20 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.02 $Y=2.335
+ $X2=8.02 $Y2=2.905
r189 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.935 $Y=2.99
+ $X2=8.02 $Y2=2.905
r190 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.935 $Y=2.99
+ $X2=7.265 $Y2=2.99
r191 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.18 $Y=2.905
+ $X2=7.265 $Y2=2.99
r192 16 37 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=7.18 $Y=2.905
+ $X2=7.18 $Y2=1.655
r193 12 44 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=11.295
+ $Y=1.885 $X2=11.22 $Y2=1.635
r194 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=11.295 $Y=1.885
+ $X2=11.295 $Y2=2.46
r195 8 44 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=11.28 $Y=1.47
+ $X2=11.22 $Y2=1.635
r196 8 10 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=11.28 $Y=1.47
+ $X2=11.28 $Y2=0.74
r197 5 35 54.7705 $w=3.67e-07 $l=3.43082e-07 $layer=POLY_cond $X=7.285 $Y=1.82
+ $X2=7.157 $Y2=1.535
r198 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.285 $Y=1.82
+ $X2=7.285 $Y2=2.315
r199 1 35 39.0103 $w=3.67e-07 $l=2.25067e-07 $layer=POLY_cond $X=7.015 $Y=1.37
+ $X2=7.157 $Y2=1.535
r200 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=7.015 $Y=1.37 $X2=7.015
+ $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%A_1092_96# 1 2 9 11 12 14 15 20 22 23 26 27
+ 28 31 32 35 37 39
c119 39 0 8.70027e-20 $X=7.75 $Y=1.255
c120 37 0 3.53193e-20 $X=6.04 $Y=1.74
c121 31 0 8.34275e-20 $X=7.75 $Y=1.42
c122 27 0 7.45928e-20 $X=7.585 $Y=1.155
c123 15 0 1.28158e-19 $X=5.955 $Y=2.37
r124 32 40 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.75 $Y=1.42
+ $X2=7.75 $Y2=1.585
r125 32 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.75 $Y=1.42
+ $X2=7.75 $Y2=1.255
r126 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.75
+ $Y=1.42 $X2=7.75 $Y2=1.42
r127 29 31 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=7.75 $Y=1.24
+ $X2=7.75 $Y2=1.42
r128 27 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.585 $Y=1.155
+ $X2=7.75 $Y2=1.24
r129 27 28 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.585 $Y=1.155
+ $X2=6.875 $Y2=1.155
r130 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.79 $Y=1.24
+ $X2=6.875 $Y2=1.155
r131 25 26 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.79 $Y=1.24
+ $X2=6.79 $Y2=1.655
r132 24 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.125 $Y=1.74
+ $X2=6.04 $Y2=1.74
r133 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.705 $Y=1.74
+ $X2=6.79 $Y2=1.655
r134 23 24 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=6.705 $Y=1.74
+ $X2=6.125 $Y2=1.74
r135 21 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.04 $Y=1.825
+ $X2=6.04 $Y2=1.74
r136 21 22 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.04 $Y=1.825
+ $X2=6.04 $Y2=2.205
r137 20 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.04 $Y=1.655
+ $X2=6.04 $Y2=1.74
r138 19 35 15.6194 $w=2.89e-07 $l=4.58432e-07 $layer=LI1_cond $X=6.04 $Y=0.855
+ $X2=5.67 $Y2=0.657
r139 19 20 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=6.04 $Y=0.855
+ $X2=6.04 $Y2=1.655
r140 15 22 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.955 $Y=2.37
+ $X2=6.04 $Y2=2.205
r141 15 17 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=5.955 $Y=2.37
+ $X2=5.77 $Y2=2.37
r142 12 14 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.825 $Y=1.82
+ $X2=7.825 $Y2=2.315
r143 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.825 $Y=1.73
+ $X2=7.825 $Y2=1.82
r144 11 40 56.3629 $w=1.8e-07 $l=1.45e-07 $layer=POLY_cond $X=7.825 $Y=1.73
+ $X2=7.825 $Y2=1.585
r145 9 39 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=7.77 $Y=0.87
+ $X2=7.77 $Y2=1.255
r146 2 17 600 $w=1.7e-07 $l=3.72659e-07 $layer=licon1_PDIFF $count=1 $X=5.54
+ $Y=2.095 $X2=5.77 $Y2=2.37
r147 1 35 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=5.46
+ $Y=0.48 $X2=5.67 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%A_1625_93# 1 2 9 11 12 14 16 17 19 20 22 24
+ 26 30 32 33 36 39 40 43 47 49
c137 49 0 8.34275e-20 $X=8.29 $Y=1.255
c138 36 0 8.70027e-20 $X=8.4 $Y=1.295
c139 32 0 1.79863e-19 $X=12.575 $Y=1.295
c140 20 0 1.08742e-19 $X=12.25 $Y=1.22
c141 12 0 2.04581e-20 $X=8.245 $Y=1.82
r142 47 50 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.29 $Y=1.42
+ $X2=8.29 $Y2=1.585
r143 47 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.29 $Y=1.42
+ $X2=8.29 $Y2=1.255
r144 40 56 16.2483 $w=4.43e-07 $l=5.9e-07 $layer=LI1_cond $X=12.8 $Y=1.295
+ $X2=12.8 $Y2=1.885
r145 40 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.61
+ $Y=1.385 $X2=12.61 $Y2=1.385
r146 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=1.295
+ $X2=12.72 $Y2=1.295
r147 36 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.29
+ $Y=1.42 $X2=8.29 $Y2=1.42
r148 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.295
+ $X2=8.4 $Y2=1.295
r149 33 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.545 $Y=1.295
+ $X2=8.4 $Y2=1.295
r150 32 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.575 $Y=1.295
+ $X2=12.72 $Y2=1.295
r151 32 33 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=12.575 $Y=1.295
+ $X2=8.545 $Y2=1.295
r152 27 30 7.45698 $w=3.38e-07 $l=2.2e-07 $layer=LI1_cond $X=12.81 $Y=0.84
+ $X2=13.03 $Y2=0.84
r153 26 40 7.99268 $w=4.43e-07 $l=1.19896e-07 $layer=LI1_cond $X=12.81 $Y=1.18
+ $X2=12.8 $Y2=1.295
r154 25 27 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=12.81 $Y=1.01
+ $X2=12.81 $Y2=0.84
r155 25 26 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=12.81 $Y=1.01
+ $X2=12.81 $Y2=1.18
r156 23 43 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=12.325 $Y=1.385
+ $X2=12.61 $Y2=1.385
r157 23 24 3.90195 $w=3.3e-07 $l=1.8735e-07 $layer=POLY_cond $X=12.325 $Y=1.385
+ $X2=12.145 $Y2=1.4
r158 20 24 34.7346 $w=1.65e-07 $l=2.26495e-07 $layer=POLY_cond $X=12.25 $Y=1.22
+ $X2=12.145 $Y2=1.4
r159 20 22 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=12.25 $Y=1.22
+ $X2=12.25 $Y2=0.74
r160 17 19 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.235 $Y=1.885
+ $X2=12.235 $Y2=2.46
r161 16 17 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.235 $Y=1.795
+ $X2=12.235 $Y2=1.885
r162 15 24 34.7346 $w=1.65e-07 $l=1.89737e-07 $layer=POLY_cond $X=12.235 $Y=1.55
+ $X2=12.145 $Y2=1.4
r163 15 16 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=12.235 $Y=1.55
+ $X2=12.235 $Y2=1.795
r164 12 14 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.245 $Y=1.82
+ $X2=8.245 $Y2=2.315
r165 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.245 $Y=1.73
+ $X2=8.245 $Y2=1.82
r166 11 50 56.3629 $w=1.8e-07 $l=1.45e-07 $layer=POLY_cond $X=8.245 $Y=1.73
+ $X2=8.245 $Y2=1.585
r167 9 49 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=8.2 $Y=0.87 $X2=8.2
+ $Y2=1.255
r168 2 56 600 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=12.86
+ $Y=1.74 $X2=12.99 $Y2=1.885
r169 1 30 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=12.885
+ $Y=0.69 $X2=13.03 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%A_622_98# 1 2 7 9 10 12 13 16 18 19 20 21
+ 22 23 25 26 27 28 30 31 33 36 39 40 41 44 47 48 49 52 54 57 60 65 66 69 70 72
+ 74 78 81 82 87
c244 78 0 4.76468e-20 $X=4.4 $Y=1.505
c245 40 0 4.96599e-20 $X=4.875 $Y=1.415
c246 33 0 2.14452e-19 $X=9.315 $Y=2.025
c247 31 0 1.28158e-19 $X=9.225 $Y=3.15
c248 28 0 1.35332e-19 $X=6.03 $Y=2.59
c249 23 0 1.65947e-19 $X=5.385 $Y=0.405
r250 81 82 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=9.435 $Y=1.335
+ $X2=9.435 $Y2=1.505
r251 79 83 14.6554 $w=2.96e-07 $l=9e-08 $layer=POLY_cond $X=4.4 $Y=1.505 $X2=4.4
+ $Y2=1.415
r252 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.4
+ $Y=1.505 $X2=4.4 $Y2=1.505
r253 75 78 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.16 $Y=1.505
+ $X2=4.4 $Y2=1.505
r254 70 87 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.32 $Y=1.065
+ $X2=10.32 $Y2=0.9
r255 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.32
+ $Y=1.065 $X2=10.32 $Y2=1.065
r256 67 69 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=10.32 $Y=0.425
+ $X2=10.32 $Y2=1.065
r257 65 67 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.155 $Y=0.34
+ $X2=10.32 $Y2=0.425
r258 65 66 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=10.155 $Y=0.34
+ $X2=9.615 $Y2=0.34
r259 63 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.53 $Y=0.425
+ $X2=9.615 $Y2=0.34
r260 63 81 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=9.53 $Y=0.425
+ $X2=9.53 $Y2=1.335
r261 60 82 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=9.42 $Y=1.775
+ $X2=9.42 $Y2=1.505
r262 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.42
+ $Y=1.775 $X2=9.42 $Y2=1.775
r263 56 75 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.16 $Y=1.67
+ $X2=4.16 $Y2=1.505
r264 56 57 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.16 $Y=1.67
+ $X2=4.16 $Y2=1.84
r265 55 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.845 $Y=1.925
+ $X2=3.68 $Y2=1.925
r266 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.075 $Y=1.925
+ $X2=4.16 $Y2=1.84
r267 54 55 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.075 $Y=1.925
+ $X2=3.845 $Y2=1.925
r268 50 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=2.01
+ $X2=3.68 $Y2=1.925
r269 50 52 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=3.68 $Y=2.01
+ $X2=3.68 $Y2=2.815
r270 48 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=1.925
+ $X2=3.68 $Y2=1.925
r271 48 49 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.515 $Y=1.925
+ $X2=3.26 $Y2=1.925
r272 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.175 $Y=1.84
+ $X2=3.26 $Y2=1.925
r273 47 72 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.175 $Y=1.84
+ $X2=3.175 $Y2=1.01
r274 42 72 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.215 $Y=0.885
+ $X2=3.215 $Y2=1.01
r275 42 44 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=0.885
+ $X2=3.215 $Y2=0.8
r276 39 87 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.23 $Y=0.58
+ $X2=10.23 $Y2=0.9
r277 34 36 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.315 $Y=3.015
+ $X2=9.315 $Y2=2.52
r278 33 61 51.2457 $w=3.23e-07 $l=2.91548e-07 $layer=POLY_cond $X=9.315 $Y=2.025
+ $X2=9.405 $Y2=1.775
r279 33 36 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.315 $Y=2.025
+ $X2=9.315 $Y2=2.52
r280 32 41 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.12 $Y=3.15 $X2=6.03
+ $Y2=3.15
r281 31 34 26.9307 $w=1.5e-07 $l=1.74284e-07 $layer=POLY_cond $X=9.225 $Y=3.15
+ $X2=9.315 $Y2=3.015
r282 31 32 1592.14 $w=1.5e-07 $l=3.105e-06 $layer=POLY_cond $X=9.225 $Y=3.15
+ $X2=6.12 $Y2=3.15
r283 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.03 $Y=2.59
+ $X2=6.03 $Y2=2.305
r284 27 41 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.03 $Y=3.075
+ $X2=6.03 $Y2=3.15
r285 26 28 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.03 $Y=2.68 $X2=6.03
+ $Y2=2.59
r286 26 27 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=6.03 $Y=2.68
+ $X2=6.03 $Y2=3.075
r287 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.385 $Y=0.405
+ $X2=5.385 $Y2=0.69
r288 21 41 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.94 $Y=3.15 $X2=6.03
+ $Y2=3.15
r289 21 22 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=5.94 $Y=3.15
+ $X2=4.95 $Y2=3.15
r290 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.31 $Y=0.33
+ $X2=5.385 $Y2=0.405
r291 19 20 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=5.31 $Y=0.33
+ $X2=4.95 $Y2=0.33
r292 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.875 $Y=3.075
+ $X2=4.95 $Y2=3.15
r293 17 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.875 $Y=1.49
+ $X2=4.875 $Y2=1.415
r294 17 18 812.734 $w=1.5e-07 $l=1.585e-06 $layer=POLY_cond $X=4.875 $Y=1.49
+ $X2=4.875 $Y2=3.075
r295 16 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.875 $Y=1.34
+ $X2=4.875 $Y2=1.415
r296 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.875 $Y=0.405
+ $X2=4.95 $Y2=0.33
r297 15 16 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=4.875 $Y=0.405
+ $X2=4.875 $Y2=1.34
r298 14 83 18.6531 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.565 $Y=1.415
+ $X2=4.4 $Y2=1.415
r299 13 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.8 $Y=1.415
+ $X2=4.875 $Y2=1.415
r300 13 14 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=4.8 $Y=1.415
+ $X2=4.565 $Y2=1.415
r301 10 79 54.0414 $w=2.96e-07 $l=2.81603e-07 $layer=POLY_cond $X=4.355 $Y=1.765
+ $X2=4.4 $Y2=1.505
r302 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.355 $Y=1.765
+ $X2=4.355 $Y2=2.4
r303 7 83 23.9164 $w=2.96e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.31 $Y=1.34
+ $X2=4.4 $Y2=1.415
r304 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.31 $Y=1.34 $X2=4.31
+ $Y2=0.86
r305 2 74 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=3.535
+ $Y=1.84 $X2=3.68 $Y2=2.005
r306 2 52 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=3.535
+ $Y=1.84 $X2=3.68 $Y2=2.815
r307 1 44 182 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_NDIFF $count=1 $X=3.11
+ $Y=0.49 $X2=3.255 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%A_877_98# 1 2 7 9 10 15 16 17 21 22 24 29
+ 31 32 38 41 46 50 51 52
c150 46 0 1.3428e-19 $X=5.325 $Y=1.53
c151 32 0 3.16672e-20 $X=4.735 $Y=1.085
c152 29 0 2.56036e-20 $X=9.87 $Y=1.295
c153 15 0 2.61122e-19 $X=5.885 $Y=0.69
c154 10 0 1.35332e-19 $X=5.81 $Y=1.44
c155 7 0 1.40154e-19 $X=5.465 $Y=2.02
r156 50 51 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=2.005
+ $X2=4.66 $Y2=1.84
r157 47 53 16.0667 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.357 $Y=1.53
+ $X2=5.357 $Y2=1.44
r158 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.325
+ $Y=1.53 $X2=5.325 $Y2=1.53
r159 44 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=1.53
+ $X2=4.82 $Y2=1.53
r160 44 46 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.905 $Y=1.53
+ $X2=5.325 $Y2=1.53
r161 42 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=1.695
+ $X2=4.82 $Y2=1.53
r162 42 51 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.82 $Y=1.695
+ $X2=4.82 $Y2=1.84
r163 41 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=1.365
+ $X2=4.82 $Y2=1.53
r164 40 41 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.82 $Y=1.17
+ $X2=4.82 $Y2=1.365
r165 36 50 1.95278 $w=4.88e-07 $l=8e-08 $layer=LI1_cond $X=4.66 $Y=2.085
+ $X2=4.66 $Y2=2.005
r166 36 38 17.8191 $w=4.88e-07 $l=7.3e-07 $layer=LI1_cond $X=4.66 $Y=2.085
+ $X2=4.66 $Y2=2.815
r167 32 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.735 $Y=1.085
+ $X2=4.82 $Y2=1.17
r168 32 34 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.735 $Y=1.085
+ $X2=4.55 $Y2=1.085
r169 27 29 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=9.685 $Y=1.295
+ $X2=9.87 $Y2=1.295
r170 25 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.87 $Y=1.37
+ $X2=9.87 $Y2=1.295
r171 25 31 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=9.87 $Y=1.37
+ $X2=9.87 $Y2=2.18
r172 22 31 103.008 $w=1.8e-07 $l=2.65e-07 $layer=POLY_cond $X=9.855 $Y=2.445
+ $X2=9.855 $Y2=2.18
r173 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.855 $Y=2.445
+ $X2=9.855 $Y2=2.73
r174 19 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.685 $Y=1.22
+ $X2=9.685 $Y2=1.295
r175 19 21 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.685 $Y=1.22
+ $X2=9.685 $Y2=0.87
r176 18 21 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=9.685 $Y=0.255
+ $X2=9.685 $Y2=0.87
r177 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.61 $Y=0.18
+ $X2=9.685 $Y2=0.255
r178 16 17 1871.6 $w=1.5e-07 $l=3.65e-06 $layer=POLY_cond $X=9.61 $Y=0.18
+ $X2=5.96 $Y2=0.18
r179 13 15 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=5.885 $Y=1.365
+ $X2=5.885 $Y2=0.69
r180 12 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.885 $Y=0.255
+ $X2=5.96 $Y2=0.18
r181 12 15 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.885 $Y=0.255
+ $X2=5.885 $Y2=0.69
r182 11 53 16.5046 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=5.525 $Y=1.44
+ $X2=5.357 $Y2=1.44
r183 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.81 $Y=1.44
+ $X2=5.885 $Y2=1.365
r184 10 11 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.81 $Y=1.44
+ $X2=5.525 $Y2=1.44
r185 7 47 96.9211 $w=2.7e-07 $l=5.41313e-07 $layer=POLY_cond $X=5.465 $Y=2.02
+ $X2=5.357 $Y2=1.53
r186 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.465 $Y=2.02
+ $X2=5.465 $Y2=2.415
r187 2 50 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=4.43
+ $Y=1.84 $X2=4.58 $Y2=2.005
r188 2 38 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.43
+ $Y=1.84 $X2=4.58 $Y2=2.815
r189 1 34 182 $w=1.7e-07 $l=6.72458e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.49 $X2=4.55 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%A_2037_442# 1 2 7 9 12 14 16 17 19 20 23 24
+ 26 27 28 30 31 33 34 37 42 43 44 46 48 49 54 58 64
r182 65 70 14.9072 $w=2.91e-07 $l=9e-08 $layer=POLY_cond $X=13.75 $Y=1.385
+ $X2=13.75 $Y2=1.295
r183 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.75
+ $Y=1.385 $X2=13.75 $Y2=1.385
r184 61 64 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=13.615 $Y=1.385
+ $X2=13.75 $Y2=1.385
r185 58 60 9.98259 $w=3.43e-07 $l=2.1e-07 $layer=LI1_cond $X=12.042 $Y=0.8
+ $X2=12.042 $Y2=1.01
r186 54 56 15.3251 $w=4.06e-07 $l=5.1e-07 $layer=LI1_cond $X=11.62 $Y=2.23
+ $X2=12.13 $Y2=2.23
r187 49 69 24.4493 $w=2.76e-07 $l=1.4e-07 $layer=POLY_cond $X=10.63 $Y=2.237
+ $X2=10.77 $Y2=2.237
r188 49 67 61.9964 $w=2.76e-07 $l=3.55e-07 $layer=POLY_cond $X=10.63 $Y=2.237
+ $X2=10.275 $Y2=2.237
r189 48 51 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=10.63 $Y=2.195
+ $X2=10.63 $Y2=2.405
r190 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.63
+ $Y=2.195 $X2=10.63 $Y2=2.195
r191 45 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.615 $Y=1.55
+ $X2=13.615 $Y2=1.385
r192 45 46 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=13.615 $Y=1.55
+ $X2=13.615 $Y2=2.14
r193 44 56 6.77762 $w=4.06e-07 $l=8.74643e-08 $layer=LI1_cond $X=12.215 $Y=2.225
+ $X2=12.13 $Y2=2.23
r194 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.53 $Y=2.225
+ $X2=13.615 $Y2=2.14
r195 43 44 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=13.53 $Y=2.225
+ $X2=12.215 $Y2=2.225
r196 42 56 5.869 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=12.13 $Y=1.97
+ $X2=12.13 $Y2=2.23
r197 42 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.13 $Y=1.97
+ $X2=12.13 $Y2=1.01
r198 38 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.795 $Y=2.405
+ $X2=10.63 $Y2=2.405
r199 37 54 6.77762 $w=4.06e-07 $l=2.13307e-07 $layer=LI1_cond $X=11.535 $Y=2.405
+ $X2=11.62 $Y2=2.23
r200 37 38 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=11.535 $Y=2.405
+ $X2=10.795 $Y2=2.405
r201 34 36 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=14.23 $Y=1.07
+ $X2=14.23 $Y2=1.295
r202 31 33 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=14.835 $Y=2.045
+ $X2=14.835 $Y2=2.54
r203 28 30 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=14.765 $Y=0.995
+ $X2=14.765 $Y2=0.645
r204 26 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.76 $Y=1.97
+ $X2=14.835 $Y2=2.045
r205 26 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=14.76 $Y=1.97
+ $X2=14.305 $Y2=1.97
r206 25 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.305 $Y=1.07
+ $X2=14.23 $Y2=1.07
r207 24 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.69 $Y=1.07
+ $X2=14.765 $Y2=0.995
r208 24 25 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=14.69 $Y=1.07
+ $X2=14.305 $Y2=1.07
r209 23 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.23 $Y=1.895
+ $X2=14.305 $Y2=1.97
r210 22 36 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.23 $Y=1.37
+ $X2=14.23 $Y2=1.295
r211 22 23 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=14.23 $Y=1.37
+ $X2=14.23 $Y2=1.895
r212 21 70 18.2534 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.915 $Y=1.295
+ $X2=13.75 $Y2=1.295
r213 20 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.155 $Y=1.295
+ $X2=14.23 $Y2=1.295
r214 20 21 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=14.155 $Y=1.295
+ $X2=13.915 $Y2=1.295
r215 17 65 57.6553 $w=2.91e-07 $l=2.89828e-07 $layer=POLY_cond $X=13.73 $Y=1.665
+ $X2=13.75 $Y2=1.385
r216 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.73 $Y=1.665
+ $X2=13.73 $Y2=2.3
r217 14 70 23.6999 $w=2.91e-07 $l=8.87412e-08 $layer=POLY_cond $X=13.72 $Y=1.22
+ $X2=13.75 $Y2=1.295
r218 14 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=13.72 $Y=1.22
+ $X2=13.72 $Y2=0.74
r219 10 69 17.0164 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.77 $Y=2.03
+ $X2=10.77 $Y2=2.237
r220 10 12 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=10.77 $Y=2.03
+ $X2=10.77 $Y2=0.58
r221 7 67 17.0164 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=10.275 $Y=2.445
+ $X2=10.275 $Y2=2.237
r222 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.275 $Y=2.445
+ $X2=10.275 $Y2=2.73
r223 2 54 300 $w=1.7e-07 $l=6.27674e-07 $layer=licon1_PDIFF $count=2 $X=11.37
+ $Y=1.96 $X2=11.62 $Y2=2.475
r224 2 54 600 $w=1.7e-07 $l=3.2596e-07 $layer=licon1_PDIFF $count=1 $X=11.37
+ $Y=1.96 $X2=11.62 $Y2=2.135
r225 1 58 182 $w=1.7e-07 $l=5.4074e-07 $layer=licon1_NDIFF $count=1 $X=11.785
+ $Y=0.37 $X2=12.035 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%A_1878_420# 1 2 7 9 10 11 12 14 19 23 25 28
+ 29 33 34 35 36 40
c117 40 0 1.08742e-19 $X=11.735 $Y=1.265
c118 35 0 1.95765e-20 $X=9.885 $Y=1.435
c119 19 0 1.44776e-20 $X=9.9 $Y=0.88
r120 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.76
+ $Y=1.385 $X2=11.76 $Y2=1.385
r121 40 43 4.93904 $w=2.78e-07 $l=1.2e-07 $layer=LI1_cond $X=11.735 $Y=1.265
+ $X2=11.735 $Y2=1.385
r122 36 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=10.8 $Y=1.265
+ $X2=10.8 $Y2=1.435
r123 33 34 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=9.855 $Y=1.675
+ $X2=9.855 $Y2=1.845
r124 29 34 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.84 $Y=2.11
+ $X2=9.84 $Y2=1.845
r125 28 31 9.24242 $w=5.48e-07 $l=4.25e-07 $layer=LI1_cond $X=9.65 $Y=2.225
+ $X2=9.65 $Y2=2.65
r126 28 29 8.74464 $w=5.48e-07 $l=1.15e-07 $layer=LI1_cond $X=9.65 $Y=2.225
+ $X2=9.65 $Y2=2.11
r127 26 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.885 $Y=1.265
+ $X2=10.8 $Y2=1.265
r128 25 40 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=11.595 $Y=1.265
+ $X2=11.735 $Y2=1.265
r129 25 26 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=11.595 $Y=1.265
+ $X2=10.885 $Y2=1.265
r130 24 35 1.64875 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=9.985 $Y=1.435
+ $X2=9.885 $Y2=1.435
r131 23 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.715 $Y=1.435
+ $X2=10.8 $Y2=1.435
r132 23 24 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=10.715 $Y=1.435
+ $X2=9.985 $Y2=1.435
r133 21 35 4.81226 $w=1.85e-07 $l=9.21954e-08 $layer=LI1_cond $X=9.87 $Y=1.52
+ $X2=9.885 $Y2=1.435
r134 21 33 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=9.87 $Y=1.52
+ $X2=9.87 $Y2=1.675
r135 17 35 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=9.885 $Y=1.35
+ $X2=9.885 $Y2=1.435
r136 17 19 26.0636 $w=1.98e-07 $l=4.7e-07 $layer=LI1_cond $X=9.885 $Y=1.35
+ $X2=9.885 $Y2=0.88
r137 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=11.845 $Y=1.885
+ $X2=11.845 $Y2=2.46
r138 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.845 $Y=1.795
+ $X2=11.845 $Y2=1.885
r139 10 44 48.8089 $w=2.97e-07 $l=2.92276e-07 $layer=POLY_cond $X=11.845 $Y=1.64
+ $X2=11.765 $Y2=1.385
r140 10 11 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=11.845 $Y=1.64
+ $X2=11.845 $Y2=1.795
r141 7 44 38.5662 $w=2.97e-07 $l=1.90526e-07 $layer=POLY_cond $X=11.71 $Y=1.22
+ $X2=11.765 $Y2=1.385
r142 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.71 $Y=1.22
+ $X2=11.71 $Y2=0.74
r143 2 31 600 $w=1.7e-07 $l=6.20484e-07 $layer=licon1_PDIFF $count=1 $X=9.39
+ $Y=2.1 $X2=9.54 $Y2=2.65
r144 2 28 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=9.39
+ $Y=2.1 $X2=9.54 $Y2=2.225
r145 1 19 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=9.76
+ $Y=0.595 $X2=9.9 $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%RESET_B 1 3 4 6 7
r32 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.21
+ $Y=1.385 $X2=13.21 $Y2=1.385
r33 7 11 3.51593 $w=2.93e-07 $l=9e-08 $layer=LI1_cond $X=13.212 $Y=1.295
+ $X2=13.212 $Y2=1.385
r34 4 10 38.6072 $w=2.91e-07 $l=1.81659e-07 $layer=POLY_cond $X=13.245 $Y=1.22
+ $X2=13.21 $Y2=1.385
r35 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=13.245 $Y=1.22
+ $X2=13.245 $Y2=0.9
r36 1 10 57.6553 $w=2.91e-07 $l=2.82489e-07 $layer=POLY_cond $X=13.215 $Y=1.665
+ $X2=13.21 $Y2=1.385
r37 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=13.215 $Y=1.665
+ $X2=13.215 $Y2=2.06
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%A_2881_74# 1 2 7 11 13 15 19 23 26 30
r50 27 30 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=14.68 $Y=1.52
+ $X2=14.68 $Y2=1.43
r51 26 29 5.14086 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=14.645 $Y=1.52
+ $X2=14.645 $Y2=1.685
r52 26 28 5.97663 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=14.645 $Y=1.52
+ $X2=14.645 $Y2=1.355
r53 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.68
+ $Y=1.52 $X2=14.68 $Y2=1.52
r54 23 29 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=14.61 $Y=2.265
+ $X2=14.61 $Y2=1.685
r55 19 28 30.305 $w=2.68e-07 $l=7.1e-07 $layer=LI1_cond $X=14.58 $Y=0.645
+ $X2=14.58 $Y2=1.355
r56 13 16 93.8489 $w=1.74e-07 $l=3.35e-07 $layer=POLY_cond $X=15.345 $Y=1.765
+ $X2=15.345 $Y2=1.43
r57 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=15.345 $Y=1.765
+ $X2=15.345 $Y2=2.4
r58 9 16 21.8259 $w=1.74e-07 $l=7.5e-08 $layer=POLY_cond $X=15.345 $Y=1.355
+ $X2=15.345 $Y2=1.43
r59 9 11 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=15.345 $Y=1.355
+ $X2=15.345 $Y2=0.74
r60 8 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.845 $Y=1.43
+ $X2=14.68 $Y2=1.43
r61 7 16 6.34751 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=15.255 $Y=1.43
+ $X2=15.345 $Y2=1.43
r62 7 8 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=15.255 $Y=1.43
+ $X2=14.845 $Y2=1.43
r63 2 23 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=14.465
+ $Y=2.12 $X2=14.61 $Y2=2.265
r64 1 19 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=14.405
+ $Y=0.37 $X2=14.55 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%A_27_464# 1 2 9 12 13 14 17 20
c41 14 0 1.00461e-19 $X=1.285 $Y=2.99
r42 15 17 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.11 $Y=2.905
+ $X2=2.11 $Y2=2.75
r43 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.945 $Y=2.99
+ $X2=2.11 $Y2=2.905
r44 13 14 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.945 $Y=2.99
+ $X2=1.285 $Y2=2.99
r45 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.2 $Y=2.905
+ $X2=1.285 $Y2=2.99
r46 11 12 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.2 $Y=2.475 $X2=1.2
+ $Y2=2.905
r47 10 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.39
+ $X2=0.28 $Y2=2.39
r48 9 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.115 $Y=2.39
+ $X2=1.2 $Y2=2.475
r49 9 10 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=2.39
+ $X2=0.445 $Y2=2.39
r50 2 17 600 $w=1.7e-07 $l=4.994e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=2.32 $X2=2.11 $Y2=2.75
r51 1 20 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.47
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54
+ 58 61 62 64 65 67 68 69 71 76 84 96 121 130 131 134 137 140 143 147 153 155
r176 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r177 152 153 11.1544 $w=7.53e-07 $l=1.65e-07 $layer=LI1_cond $X=10.985 $Y=3.037
+ $X2=11.15 $Y2=3.037
r178 149 152 2.93079 $w=7.53e-07 $l=1.85e-07 $layer=LI1_cond $X=10.8 $Y=3.037
+ $X2=10.985 $Y2=3.037
r179 149 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r180 146 149 3.16842 $w=7.53e-07 $l=2e-07 $layer=LI1_cond $X=10.6 $Y=3.037
+ $X2=10.8 $Y2=3.037
r181 146 147 11.1544 $w=7.53e-07 $l=1.65e-07 $layer=LI1_cond $X=10.6 $Y=3.037
+ $X2=10.435 $Y2=3.037
r182 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r183 140 141 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r184 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r185 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r186 131 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=15.12 $Y2=3.33
r187 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r188 128 155 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=15.205 $Y=3.33
+ $X2=15.075 $Y2=3.33
r189 128 130 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=15.205 $Y=3.33
+ $X2=15.6 $Y2=3.33
r190 127 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r191 126 127 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r192 124 127 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.64 $Y2=3.33
r193 123 126 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=13.68 $Y=3.33
+ $X2=14.64 $Y2=3.33
r194 123 124 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r195 121 155 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=14.945 $Y=3.33
+ $X2=15.075 $Y2=3.33
r196 121 126 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=14.945 $Y=3.33
+ $X2=14.64 $Y2=3.33
r197 120 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r198 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r199 117 120 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=13.2 $Y2=3.33
r200 116 117 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r201 114 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r202 114 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r203 113 116 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r204 113 153 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=11.28 $Y=3.33
+ $X2=11.15 $Y2=3.33
r205 113 114 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r206 110 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r207 109 147 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=10.32 $Y=3.33
+ $X2=10.435 $Y2=3.33
r208 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r209 107 110 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r210 107 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r211 106 109 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r212 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r213 104 143 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.685 $Y=3.33
+ $X2=8.5 $Y2=3.33
r214 104 106 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.685 $Y=3.33
+ $X2=8.88 $Y2=3.33
r215 98 101 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r216 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r217 96 143 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.315 $Y=3.33
+ $X2=8.5 $Y2=3.33
r218 96 101 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.315 $Y=3.33
+ $X2=7.92 $Y2=3.33
r219 95 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r220 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r221 92 95 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r222 92 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r223 91 94 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r224 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r225 89 140 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.215 $Y=3.33
+ $X2=4.13 $Y2=3.33
r226 89 91 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.215 $Y=3.33
+ $X2=4.56 $Y2=3.33
r227 88 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r228 88 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r229 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r230 85 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.63 $Y2=3.33
r231 85 87 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=3.12 $Y2=3.33
r232 84 140 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=4.13 $Y2=3.33
r233 84 87 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=3.12 $Y2=3.33
r234 83 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r235 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r236 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r237 80 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r238 79 82 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r239 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r240 77 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r241 77 79 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r242 76 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.63 $Y2=3.33
r243 76 82 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.16 $Y2=3.33
r244 74 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r245 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r246 71 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r247 71 73 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r248 69 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r249 69 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=6.96 $Y2=3.33
r250 69 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r251 67 119 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=13.34 $Y=3.33
+ $X2=13.2 $Y2=3.33
r252 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.34 $Y=3.33
+ $X2=13.505 $Y2=3.33
r253 66 123 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=13.67 $Y=3.33
+ $X2=13.68 $Y2=3.33
r254 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.67 $Y=3.33
+ $X2=13.505 $Y2=3.33
r255 64 116 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=12.295 $Y=3.33
+ $X2=12.24 $Y2=3.33
r256 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.295 $Y=3.33
+ $X2=12.46 $Y2=3.33
r257 63 119 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=12.625 $Y=3.33
+ $X2=13.2 $Y2=3.33
r258 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.625 $Y=3.33
+ $X2=12.46 $Y2=3.33
r259 61 94 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.595 $Y=3.33
+ $X2=6.48 $Y2=3.33
r260 61 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.595 $Y=3.33
+ $X2=6.76 $Y2=3.33
r261 60 98 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.925 $Y=3.33
+ $X2=6.96 $Y2=3.33
r262 60 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.925 $Y=3.33
+ $X2=6.76 $Y2=3.33
r263 56 155 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=15.075 $Y=3.245
+ $X2=15.075 $Y2=3.33
r264 56 58 42.7734 $w=2.58e-07 $l=9.65e-07 $layer=LI1_cond $X=15.075 $Y=3.245
+ $X2=15.075 $Y2=2.28
r265 52 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.505 $Y=3.245
+ $X2=13.505 $Y2=3.33
r266 52 54 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=13.505 $Y=3.245
+ $X2=13.505 $Y2=2.645
r267 48 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.46 $Y=3.245
+ $X2=12.46 $Y2=3.33
r268 48 50 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=12.46 $Y=3.245
+ $X2=12.46 $Y2=2.645
r269 44 143 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.5 $Y=3.245
+ $X2=8.5 $Y2=3.33
r270 44 46 20.4014 $w=3.68e-07 $l=6.55e-07 $layer=LI1_cond $X=8.5 $Y=3.245
+ $X2=8.5 $Y2=2.59
r271 40 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.76 $Y=3.245
+ $X2=6.76 $Y2=3.33
r272 40 42 35.0971 $w=3.28e-07 $l=1.005e-06 $layer=LI1_cond $X=6.76 $Y=3.245
+ $X2=6.76 $Y2=2.24
r273 36 140 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=3.245
+ $X2=4.13 $Y2=3.33
r274 36 38 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=4.13 $Y=3.245
+ $X2=4.13 $Y2=2.345
r275 32 137 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=3.245
+ $X2=2.63 $Y2=3.33
r276 32 34 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.63 $Y=3.245
+ $X2=2.63 $Y2=2.75
r277 28 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r278 28 30 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.77
r279 9 58 300 $w=1.7e-07 $l=2.73542e-07 $layer=licon1_PDIFF $count=2 $X=14.91
+ $Y=2.12 $X2=15.115 $Y2=2.28
r280 8 54 600 $w=1.7e-07 $l=1.00678e-06 $layer=licon1_PDIFF $count=1 $X=13.29
+ $Y=1.74 $X2=13.505 $Y2=2.645
r281 7 50 600 $w=1.7e-07 $l=7.5629e-07 $layer=licon1_PDIFF $count=1 $X=12.31
+ $Y=1.96 $X2=12.46 $Y2=2.645
r282 6 152 600 $w=1.7e-07 $l=7.72593e-07 $layer=licon1_PDIFF $count=1 $X=10.35
+ $Y=2.52 $X2=10.985 $Y2=2.825
r283 6 146 600 $w=1.7e-07 $l=4.1143e-07 $layer=licon1_PDIFF $count=1 $X=10.35
+ $Y=2.52 $X2=10.6 $Y2=2.825
r284 5 46 600 $w=1.7e-07 $l=7.79824e-07 $layer=licon1_PDIFF $count=1 $X=8.32
+ $Y=1.895 $X2=8.5 $Y2=2.59
r285 4 42 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=6.525
+ $Y=2.095 $X2=6.76 $Y2=2.24
r286 3 38 300 $w=1.7e-07 $l=5.7513e-07 $layer=licon1_PDIFF $count=2 $X=3.98
+ $Y=1.84 $X2=4.13 $Y2=2.345
r287 2 34 600 $w=1.7e-07 $l=4.97242e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=2.32 $X2=2.67 $Y2=2.75
r288 1 30 600 $w=1.7e-07 $l=5.40833e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.32 $X2=0.78 $Y2=2.77
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%A_197_119# 1 2 3 4 15 17 18 21 23 24 26 28
+ 29 30 32 34 37 40 41 42 43 44 46 48 52 53
c172 53 0 1.86601e-19 $X=5.25 $Y=0.645
c173 46 0 4.96599e-20 $X=5.7 $Y=1.865
r174 51 53 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=5.17 $Y=0.645
+ $X2=5.25 $Y2=0.645
r175 51 52 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.17 $Y=0.645
+ $X2=5.005 $Y2=0.645
r176 47 48 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.02 $Y=1.27
+ $X2=2.335 $Y2=1.27
r177 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.7 $Y=1.195
+ $X2=5.7 $Y2=1.865
r178 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.615 $Y=1.95
+ $X2=5.7 $Y2=1.865
r179 43 44 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.615 $Y=1.95
+ $X2=5.405 $Y2=1.95
r180 41 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.615 $Y=1.11
+ $X2=5.7 $Y2=1.195
r181 41 42 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.615 $Y=1.11
+ $X2=5.335 $Y2=1.11
r182 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.25 $Y=1.025
+ $X2=5.335 $Y2=1.11
r183 39 53 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.25 $Y=0.83
+ $X2=5.25 $Y2=0.645
r184 39 40 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.25 $Y=0.83
+ $X2=5.25 $Y2=1.025
r185 35 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.24 $Y=2.035
+ $X2=5.405 $Y2=1.95
r186 35 37 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=5.24 $Y=2.035
+ $X2=5.24 $Y2=2.24
r187 34 52 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=3.68 $Y=0.745
+ $X2=5.005 $Y2=0.745
r188 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.595 $Y=0.66
+ $X2=3.68 $Y2=0.745
r189 31 32 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.595 $Y=0.425
+ $X2=3.595 $Y2=0.66
r190 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.51 $Y=0.34
+ $X2=3.595 $Y2=0.425
r191 29 30 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=3.51 $Y=0.34
+ $X2=2.42 $Y2=0.34
r192 28 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.335 $Y=1.185
+ $X2=2.335 $Y2=1.27
r193 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.335 $Y=0.425
+ $X2=2.42 $Y2=0.34
r194 27 28 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.335 $Y=0.425
+ $X2=2.335 $Y2=1.185
r195 25 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=1.355
+ $X2=2.02 $Y2=1.27
r196 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.02 $Y=1.355
+ $X2=2.02 $Y2=2.025
r197 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.935 $Y=2.11
+ $X2=2.02 $Y2=2.025
r198 23 24 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.935 $Y=2.11
+ $X2=1.745 $Y2=2.11
r199 19 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.62 $Y=2.195
+ $X2=1.745 $Y2=2.11
r200 19 21 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=1.62 $Y=2.195
+ $X2=1.62 $Y2=2.515
r201 17 47 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.935 $Y=1.27
+ $X2=2.02 $Y2=1.27
r202 17 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.935 $Y=1.27
+ $X2=1.37 $Y2=1.27
r203 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.205 $Y=1.185
+ $X2=1.37 $Y2=1.27
r204 13 15 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.205 $Y=1.185
+ $X2=1.205 $Y2=0.805
r205 4 37 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.095
+ $Y=2.095 $X2=5.24 $Y2=2.24
r206 3 21 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=2.32 $X2=1.66 $Y2=2.515
r207 2 51 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=5.025
+ $Y=0.48 $X2=5.17 $Y2=0.645
r208 1 15 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.595 $X2=1.205 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%Q_N 1 2 10 15 16 17 18 19
r37 19 28 1.70732 $w=4.03e-07 $l=6e-08 $layer=LI1_cond $X=14.072 $Y=2.775
+ $X2=14.072 $Y2=2.715
r38 18 28 8.82117 $w=4.03e-07 $l=3.1e-07 $layer=LI1_cond $X=14.072 $Y=2.405
+ $X2=14.072 $Y2=2.715
r39 17 18 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=14.072 $Y=2.035
+ $X2=14.072 $Y2=2.405
r40 15 16 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=14.072 $Y=1.885
+ $X2=14.072 $Y2=1.72
r41 13 17 3.21546 $w=4.03e-07 $l=1.13e-07 $layer=LI1_cond $X=14.072 $Y=1.922
+ $X2=14.072 $Y2=2.035
r42 13 15 1.05285 $w=4.03e-07 $l=3.7e-08 $layer=LI1_cond $X=14.072 $Y=1.922
+ $X2=14.072 $Y2=1.885
r43 12 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.19 $Y=1.05
+ $X2=14.19 $Y2=1.72
r44 10 12 18.3112 $w=5.03e-07 $l=5.35e-07 $layer=LI1_cond $X=14.022 $Y=0.515
+ $X2=14.022 $Y2=1.05
r45 2 28 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.805
+ $Y=1.74 $X2=13.955 $Y2=2.715
r46 2 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.805
+ $Y=1.74 $X2=13.955 $Y2=1.885
r47 1 10 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.795
+ $Y=0.37 $X2=13.935 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%Q 1 2 7 8 9 10 11 12 13
r16 12 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=15.565 $Y=2.405
+ $X2=15.565 $Y2=2.775
r17 11 12 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=15.565 $Y=1.985
+ $X2=15.565 $Y2=2.405
r18 10 11 10.8465 $w=3.38e-07 $l=3.2e-07 $layer=LI1_cond $X=15.565 $Y=1.665
+ $X2=15.565 $Y2=1.985
r19 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=15.565 $Y=1.295
+ $X2=15.565 $Y2=1.665
r20 8 9 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=15.565 $Y=0.925
+ $X2=15.565 $Y2=1.295
r21 7 8 13.8971 $w=3.38e-07 $l=4.1e-07 $layer=LI1_cond $X=15.565 $Y=0.515
+ $X2=15.565 $Y2=0.925
r22 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=15.42
+ $Y=1.84 $X2=15.57 $Y2=2.815
r23 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=15.42
+ $Y=1.84 $X2=15.57 $Y2=1.985
r24 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.42
+ $Y=0.37 $X2=15.56 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%VGND 1 2 3 4 5 6 7 8 25 27 31 35 39 43 47
+ 53 57 62 63 65 66 68 69 71 72 74 75 76 85 117 126 127 133 136
c169 43 0 3.45888e-20 $X=9.11 $Y=0.845
c170 4 0 7.45928e-20 $X=6.435 $Y=0.625
r171 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r172 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r173 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r174 127 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=15.12 $Y2=0
r175 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r176 124 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.225 $Y=0
+ $X2=15.06 $Y2=0
r177 124 126 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=15.225 $Y=0
+ $X2=15.6 $Y2=0
r178 123 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.12 $Y2=0
r179 122 123 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r180 120 123 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.64 $Y2=0
r181 119 122 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=13.68 $Y=0
+ $X2=14.64 $Y2=0
r182 119 120 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r183 117 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.895 $Y=0
+ $X2=15.06 $Y2=0
r184 117 122 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=14.895 $Y=0
+ $X2=14.64 $Y2=0
r185 116 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r186 115 116 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r187 113 116 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=13.2 $Y2=0
r188 112 115 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=11.28 $Y=0
+ $X2=13.2 $Y2=0
r189 112 113 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r190 110 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r191 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r192 107 110 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=10.8 $Y2=0
r193 106 109 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=10.8 $Y2=0
r194 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r195 104 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r196 103 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r197 100 103 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.96 $Y=0
+ $X2=8.88 $Y2=0
r198 100 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r199 98 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r200 97 98 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r201 95 98 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=6.48 $Y2=0
r202 95 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=4.08 $Y2=0
r203 94 97 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r204 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r205 92 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.18 $Y=0
+ $X2=4.015 $Y2=0
r206 92 94 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.18 $Y=0 $X2=4.56
+ $Y2=0
r207 91 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r208 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r209 88 91 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r210 87 90 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r211 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r212 85 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.85 $Y=0
+ $X2=4.015 $Y2=0
r213 85 90 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.85 $Y=0 $X2=3.6
+ $Y2=0
r214 84 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r215 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r216 81 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r217 81 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r218 80 83 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r219 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r220 78 130 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=0
+ $X2=0.235 $Y2=0
r221 78 80 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.72
+ $Y2=0
r222 76 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.88 $Y2=0
r223 76 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=6.96 $Y2=0
r224 74 115 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=13.295 $Y=0
+ $X2=13.2 $Y2=0
r225 74 75 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=13.295 $Y=0
+ $X2=13.442 $Y2=0
r226 73 119 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=13.59 $Y=0 $X2=13.68
+ $Y2=0
r227 73 75 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=13.59 $Y=0
+ $X2=13.442 $Y2=0
r228 71 109 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=10.9 $Y=0 $X2=10.8
+ $Y2=0
r229 71 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.9 $Y=0
+ $X2=11.025 $Y2=0
r230 70 112 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=11.15 $Y=0
+ $X2=11.28 $Y2=0
r231 70 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.15 $Y=0
+ $X2=11.025 $Y2=0
r232 68 103 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=9.025 $Y=0
+ $X2=8.88 $Y2=0
r233 68 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.025 $Y=0 $X2=9.15
+ $Y2=0
r234 67 106 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=9.275 $Y=0
+ $X2=9.36 $Y2=0
r235 67 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.275 $Y=0 $X2=9.15
+ $Y2=0
r236 65 97 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=6.49 $Y=0 $X2=6.48
+ $Y2=0
r237 65 66 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=6.49 $Y=0 $X2=6.687
+ $Y2=0
r238 64 100 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.885 $Y=0
+ $X2=6.96 $Y2=0
r239 64 66 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=6.885 $Y=0
+ $X2=6.687 $Y2=0
r240 62 83 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=1.68
+ $Y2=0
r241 62 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=1.955
+ $Y2=0
r242 61 87 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.08 $Y=0 $X2=2.16
+ $Y2=0
r243 61 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.08 $Y=0 $X2=1.955
+ $Y2=0
r244 57 59 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=15.06 $Y=0.495
+ $X2=15.06 $Y2=0.855
r245 55 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.06 $Y=0.085
+ $X2=15.06 $Y2=0
r246 55 57 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=15.06 $Y=0.085
+ $X2=15.06 $Y2=0.495
r247 51 75 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=13.442 $Y=0.085
+ $X2=13.442 $Y2=0
r248 51 53 29.2994 $w=2.93e-07 $l=7.5e-07 $layer=LI1_cond $X=13.442 $Y=0.085
+ $X2=13.442 $Y2=0.835
r249 47 49 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=11.025 $Y=0.505
+ $X2=11.025 $Y2=0.845
r250 45 72 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.025 $Y=0.085
+ $X2=11.025 $Y2=0
r251 45 47 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=11.025 $Y=0.085
+ $X2=11.025 $Y2=0.505
r252 41 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.15 $Y=0.085
+ $X2=9.15 $Y2=0
r253 41 43 35.0343 $w=2.48e-07 $l=7.6e-07 $layer=LI1_cond $X=9.15 $Y=0.085
+ $X2=9.15 $Y2=0.845
r254 37 66 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.687 $Y=0.085
+ $X2=6.687 $Y2=0
r255 37 39 11.3786 $w=3.93e-07 $l=3.9e-07 $layer=LI1_cond $X=6.687 $Y=0.085
+ $X2=6.687 $Y2=0.475
r256 33 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.015 $Y=0.085
+ $X2=4.015 $Y2=0
r257 33 35 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.015 $Y=0.085
+ $X2=4.015 $Y2=0.325
r258 29 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=0.085
+ $X2=1.955 $Y2=0
r259 29 31 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=1.955 $Y=0.085
+ $X2=1.955 $Y2=0.795
r260 25 130 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.305 $Y=0.085
+ $X2=0.235 $Y2=0
r261 25 27 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.305 $Y=0.085
+ $X2=0.305 $Y2=0.765
r262 8 59 182 $w=1.7e-07 $l=5.84744e-07 $layer=licon1_NDIFF $count=1 $X=14.84
+ $Y=0.37 $X2=15.06 $Y2=0.855
r263 8 57 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=14.84
+ $Y=0.37 $X2=15.06 $Y2=0.495
r264 7 53 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=13.32
+ $Y=0.69 $X2=13.48 $Y2=0.835
r265 6 49 182 $w=1.7e-07 $l=5.74565e-07 $layer=licon1_NDIFF $count=1 $X=10.845
+ $Y=0.37 $X2=11.065 $Y2=0.845
r266 6 47 182 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=1 $X=10.845
+ $Y=0.37 $X2=11.065 $Y2=0.505
r267 5 43 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=8.965
+ $Y=0.595 $X2=9.11 $Y2=0.845
r268 4 39 182 $w=1.7e-07 $l=3.16228e-07 $layer=licon1_NDIFF $count=1 $X=6.435
+ $Y=0.625 $X2=6.685 $Y2=0.475
r269 3 35 182 $w=1.7e-07 $l=5.46306e-07 $layer=licon1_NDIFF $count=1 $X=3.545
+ $Y=0.49 $X2=4.015 $Y2=0.325
r270 2 31 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1.855
+ $Y=0.595 $X2=1.995 $Y2=0.795
r271 1 27 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.595 $X2=0.305 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%A_1418_125# 1 2 7 13 15 16
c24 15 0 1.14272e-19 $X=8.52 $Y=0.475
r25 15 16 9.94572 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=8.52 $Y=0.435
+ $X2=8.33 $Y2=0.435
r26 13 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.64 $Y=0.395
+ $X2=8.33 $Y2=0.395
r27 7 13 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=7.515 $Y=0.435
+ $X2=7.64 $Y2=0.435
r28 7 9 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=7.515 $Y=0.435
+ $X2=7.39 $Y2=0.435
r29 2 15 182 $w=1.7e-07 $l=2.9904e-07 $layer=licon1_NDIFF $count=1 $X=8.275
+ $Y=0.595 $X2=8.52 $Y2=0.475
r30 1 9 182 $w=1.7e-07 $l=3.67423e-07 $layer=licon1_NDIFF $count=1 $X=7.09
+ $Y=0.625 $X2=7.39 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_LS__SDFBBP_1%A_2271_74# 1 2 9 11 12 15
r26 13 15 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=12.47 $Y=0.425
+ $X2=12.47 $Y2=0.505
r27 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.385 $Y=0.34
+ $X2=12.47 $Y2=0.425
r28 11 12 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=12.385 $Y=0.34
+ $X2=11.66 $Y2=0.34
r29 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.495 $Y=0.425
+ $X2=11.66 $Y2=0.34
r30 7 9 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=11.495 $Y=0.425
+ $X2=11.495 $Y2=0.505
r31 2 15 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=12.325
+ $Y=0.37 $X2=12.47 $Y2=0.505
r32 1 9 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=11.355
+ $Y=0.37 $X2=11.495 $Y2=0.505
.ends

