* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 X a_187_338# VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=1.34918e+12p ps=1.097e+07u
M1001 VPWR A1 a_596_392# VPB phighvt w=1e+06u l=150000u
+  ad=1.642e+12p pd=1.38e+07u as=1.15e+12p ps=1.03e+07u
M1002 VPWR a_187_338# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.72e+11p ps=5.68e+06u
M1003 VGND a_187_338# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND B1_N a_29_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1005 a_864_123# A1 a_187_338# VNB nshort w=640000u l=150000u
+  ad=3.968e+11p pd=3.8e+06u as=3.584e+11p ps=3.68e+06u
M1006 X a_187_338# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_864_123# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_187_338# a_29_392# a_596_392# VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1009 a_596_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_187_338# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_187_338# A1 a_864_123# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_187_338# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_596_392# a_29_392# a_187_338# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_29_392# a_187_338# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_187_338# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A2 a_596_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_864_123# A2 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_187_338# a_29_392# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR B1_N a_29_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1020 X a_187_338# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_596_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
