* File: sky130_fd_sc_ls__a222o_1.pex.spice
* Created: Fri Aug 28 12:54:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A222O_1%C1 2 3 5 8 9 10 14 15 16
c30 15 0 1.41241e-19 $X=0.385 $Y=1.285
r31 14 17 39.5669 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.285
+ $X2=0.407 $Y2=1.45
r32 14 16 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.285
+ $X2=0.407 $Y2=1.12
r33 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.285 $X2=0.385 $Y2=1.285
r34 9 10 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.665
r35 9 15 0.271163 $w=4.23e-07 $l=1e-08 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.285
r36 8 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.52 $Y=0.69 $X2=0.52
+ $Y2=1.12
r37 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.875
+ $X2=0.505 $Y2=2.45
r38 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.785 $X2=0.505
+ $Y2=1.875
r39 2 17 130.218 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=0.505 $Y=1.785
+ $X2=0.505 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LS__A222O_1%C2 1 3 5 6 8 9 12
c43 12 0 1.41241e-19 $X=1.11 $Y=1.285
r44 12 14 20.5296 $w=2.7e-07 $l=1.15e-07 $layer=POLY_cond $X=1.11 $Y=1.285
+ $X2=1.225 $Y2=1.285
r45 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.225
+ $Y=1.285 $X2=1.225 $Y2=1.285
r46 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.11 $Y=1.875
+ $X2=1.11 $Y2=2.45
r47 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.11 $Y=1.785 $X2=1.11
+ $Y2=1.875
r48 4 12 12.2893 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.11 $Y=1.45
+ $X2=1.11 $Y2=1.285
r49 4 5 130.218 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=1.11 $Y=1.45 $X2=1.11
+ $Y2=1.785
r50 1 12 35.7037 $w=2.7e-07 $l=2.70185e-07 $layer=POLY_cond $X=0.91 $Y=1.12
+ $X2=1.11 $Y2=1.285
r51 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.91 $Y=1.12 $X2=0.91
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__A222O_1%B2 1 3 5 8 10 12 15
c49 10 0 1.60193e-19 $X=1.61 $Y=1.782
c50 1 0 1.93956e-19 $X=1.61 $Y=1.875
r51 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.345
+ $X2=1.765 $Y2=1.51
r52 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.345
+ $X2=1.765 $Y2=1.18
r53 12 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.765
+ $Y=1.345 $X2=1.765 $Y2=1.345
r54 10 11 17.7006 $w=1.77e-07 $l=6.5e-08 $layer=POLY_cond $X=1.61 $Y=1.782
+ $X2=1.675 $Y2=1.782
r55 8 17 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.855 $Y=0.69
+ $X2=1.855 $Y2=1.18
r56 5 11 6.7465 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=1.675 $Y=1.69
+ $X2=1.675 $Y2=1.782
r57 5 18 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.675 $Y=1.69
+ $X2=1.675 $Y2=1.51
r58 1 10 6.7465 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=1.61 $Y=1.875 $X2=1.61
+ $Y2=1.782
r59 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.61 $Y=1.875
+ $X2=1.61 $Y2=2.45
.ends

.subckt PM_SKY130_FD_SC_LS__A222O_1%B1 3 8 9 10 11 12 16 17 18
c42 17 0 1.60193e-19 $X=2.385 $Y=1.285
r43 16 19 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.345 $Y=1.285
+ $X2=2.345 $Y2=1.45
r44 16 18 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.345 $Y=1.285
+ $X2=2.345 $Y2=1.12
r45 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.385
+ $Y=1.285 $X2=2.385 $Y2=1.285
r46 11 12 8.27194 $w=5.33e-07 $l=3.7e-07 $layer=LI1_cond $X=2.487 $Y=1.295
+ $X2=2.487 $Y2=1.665
r47 11 17 0.223566 $w=5.33e-07 $l=1e-08 $layer=LI1_cond $X=2.487 $Y=1.295
+ $X2=2.487 $Y2=1.285
r48 9 10 37.0276 $w=1.65e-07 $l=8.5e-08 $layer=POLY_cond $X=2.207 $Y=1.79
+ $X2=2.207 $Y2=1.875
r49 9 19 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.215 $Y=1.79
+ $X2=2.215 $Y2=1.45
r50 8 18 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.245 $Y=0.69
+ $X2=2.245 $Y2=1.12
r51 3 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.2 $Y=2.45 $X2=2.2
+ $Y2=1.875
.ends

.subckt PM_SKY130_FD_SC_LS__A222O_1%A1 3 5 6 8 11 13 16 18
c38 13 0 7.1933e-20 $X=3.12 $Y=1.295
r39 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.285
+ $X2=3.09 $Y2=1.45
r40 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.285
+ $X2=3.09 $Y2=1.12
r41 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.285 $X2=3.09 $Y2=1.285
r42 9 11 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=3.18 $Y=1.765 $X2=3.26
+ $Y2=1.765
r43 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.26 $Y=1.84 $X2=3.26
+ $Y2=1.765
r44 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.26 $Y=1.84 $X2=3.26
+ $Y2=2.415
r45 5 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.18 $Y=1.69 $X2=3.18
+ $Y2=1.765
r46 5 19 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.18 $Y=1.69 $X2=3.18
+ $Y2=1.45
r47 3 18 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.18 $Y=0.69 $X2=3.18
+ $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LS__A222O_1%A2 3 5 6 8 9 12 14
c41 5 0 7.1933e-20 $X=3.71 $Y=1.75
r42 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.66 $Y=1.285
+ $X2=3.66 $Y2=1.45
r43 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.66 $Y=1.285
+ $X2=3.66 $Y2=1.12
r44 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.66
+ $Y=1.285 $X2=3.66 $Y2=1.285
r45 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.71 $Y=1.84 $X2=3.71
+ $Y2=2.415
r46 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.71 $Y=1.75 $X2=3.71
+ $Y2=1.84
r47 5 15 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=3.71 $Y=1.75 $X2=3.71
+ $Y2=1.45
r48 3 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.57 $Y=0.69 $X2=3.57
+ $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LS__A222O_1%A_32_74# 1 2 3 10 12 15 19 21 22 27 31 34 35
+ 36 39 40 44
c103 27 0 1.93956e-19 $X=0.885 $Y=2.095
r104 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.205
+ $Y=1.465 $X2=4.205 $Y2=1.465
r105 41 44 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=4.1 $Y=1.465
+ $X2=4.205 $Y2=1.465
r106 38 40 10.2865 $w=6.18e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=0.64
+ $X2=3.13 $Y2=0.64
r107 38 39 20.0288 $w=6.18e-07 $l=6.7e-07 $layer=LI1_cond $X=2.965 $Y=0.64
+ $X2=2.295 $Y2=0.64
r108 34 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.1 $Y=1.3 $X2=4.1
+ $Y2=1.465
r109 33 34 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.1 $Y=0.95 $X2=4.1
+ $Y2=1.3
r110 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.015 $Y=0.865
+ $X2=4.1 $Y2=0.95
r111 31 40 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=4.015 $Y=0.865
+ $X2=3.13 $Y2=0.865
r112 30 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=0.865
+ $X2=0.805 $Y2=0.865
r113 30 39 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=0.89 $Y=0.865
+ $X2=2.295 $Y2=0.865
r114 27 36 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=2.095
+ $X2=0.885 $Y2=1.93
r115 23 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0.95
+ $X2=0.805 $Y2=0.865
r116 23 36 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=0.805 $Y=0.95
+ $X2=0.805 $Y2=1.93
r117 21 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.865
+ $X2=0.805 $Y2=0.865
r118 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.72 $Y=0.865
+ $X2=0.47 $Y2=0.865
r119 17 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.305 $Y=0.78
+ $X2=0.47 $Y2=0.865
r120 17 19 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.305 $Y=0.78
+ $X2=0.305 $Y2=0.515
r121 13 45 38.5662 $w=2.97e-07 $l=2.06325e-07 $layer=POLY_cond $X=4.305 $Y=1.3
+ $X2=4.212 $Y2=1.465
r122 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.305 $Y=1.3
+ $X2=4.305 $Y2=0.74
r123 10 45 60.4753 $w=2.97e-07 $l=3.38969e-07 $layer=POLY_cond $X=4.295 $Y=1.765
+ $X2=4.212 $Y2=1.465
r124 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.295 $Y=1.765
+ $X2=4.295 $Y2=2.4
r125 3 27 300 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.95 $X2=0.885 $Y2=2.095
r126 2 38 45.5 $w=1.7e-07 $l=7.04734e-07 $layer=licon1_NDIFF $count=4 $X=2.32
+ $Y=0.37 $X2=2.965 $Y2=0.495
r127 1 19 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.37 $X2=0.305 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A222O_1%A_27_390# 1 2 3 12 16 17 20 24 28 30
r45 26 28 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.425 $Y=2.905
+ $X2=2.425 $Y2=2.465
r46 25 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=2.99
+ $X2=1.385 $Y2=2.99
r47 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.26 $Y=2.99
+ $X2=2.425 $Y2=2.905
r48 24 25 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.26 $Y=2.99
+ $X2=1.55 $Y2=2.99
r49 20 23 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.385 $Y=2.095
+ $X2=1.385 $Y2=2.805
r50 18 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.385 $Y=2.905
+ $X2=1.385 $Y2=2.99
r51 18 23 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.385 $Y=2.905
+ $X2=1.385 $Y2=2.805
r52 16 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.22 $Y=2.99
+ $X2=1.385 $Y2=2.99
r53 16 17 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.22 $Y=2.99
+ $X2=0.445 $Y2=2.99
r54 12 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.28 $Y=2.125
+ $X2=0.28 $Y2=2.805
r55 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r56 10 15 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=0.28 $Y=2.905 $X2=0.28
+ $Y2=2.805
r57 3 28 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=2.275
+ $Y=1.95 $X2=2.425 $Y2=2.465
r58 2 23 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=1.185
+ $Y=1.95 $X2=1.385 $Y2=2.805
r59 2 20 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=1.185
+ $Y=1.95 $X2=1.385 $Y2=2.095
r60 1 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.95 $X2=0.28 $Y2=2.805
r61 1 12 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.95 $X2=0.28 $Y2=2.125
.ends

.subckt PM_SKY130_FD_SC_LS__A222O_1%A_337_390# 1 2 9 11 13 16
r36 11 18 2.90003 $w=3.3e-07 $l=1.18e-07 $layer=LI1_cond $X=3.485 $Y=2.13
+ $X2=3.485 $Y2=2.012
r37 11 13 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=3.485 $Y=2.13
+ $X2=3.485 $Y2=2.77
r38 10 16 4.99254 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.05 $Y=2.045
+ $X2=1.885 $Y2=2.03
r39 9 18 4.86615 $w=1.7e-07 $l=1.80748e-07 $layer=LI1_cond $X=3.32 $Y=2.045
+ $X2=3.485 $Y2=2.012
r40 9 10 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=3.32 $Y=2.045
+ $X2=2.05 $Y2=2.045
r41 2 18 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.335
+ $Y=1.915 $X2=3.485 $Y2=2.06
r42 2 13 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.335
+ $Y=1.915 $X2=3.485 $Y2=2.77
r43 1 16 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=1.685
+ $Y=1.95 $X2=1.885 $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_LS__A222O_1%VPWR 1 2 9 13 18 19 20 29 35 36 39
r48 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r49 36 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r50 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r51 33 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.02 $Y2=3.33
r52 33 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.56 $Y2=3.33
r53 32 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r54 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r55 29 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=4.02 $Y2=3.33
r56 29 31 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=3.6 $Y2=3.33
r57 28 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 23 27 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 23 24 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 20 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r62 20 24 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 18 27 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.82 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.82 $Y=3.33
+ $X2=2.985 $Y2=3.33
r65 17 31 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.15 $Y=3.33 $X2=3.6
+ $Y2=3.33
r66 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=3.33
+ $X2=2.985 $Y2=3.33
r67 13 16 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=4.02 $Y=2.06
+ $X2=4.02 $Y2=2.815
r68 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=3.245
+ $X2=4.02 $Y2=3.33
r69 11 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.02 $Y=3.245
+ $X2=4.02 $Y2=2.815
r70 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=3.245
+ $X2=2.985 $Y2=3.33
r71 7 9 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=2.985 $Y=3.245
+ $X2=2.985 $Y2=2.385
r72 2 16 400 $w=1.7e-07 $l=1.01069e-06 $layer=licon1_PDIFF $count=1 $X=3.785
+ $Y=1.915 $X2=4.02 $Y2=2.815
r73 2 13 400 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=3.785
+ $Y=1.915 $X2=4.02 $Y2=2.06
r74 1 9 300 $w=1.7e-07 $l=5.37634e-07 $layer=licon1_PDIFF $count=2 $X=2.84
+ $Y=1.915 $X2=2.985 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_LS__A222O_1%X 1 2 9 13 14 15 16 23 32
r25 21 23 1.2336 $w=3.53e-07 $l=3.8e-08 $layer=LI1_cond $X=4.532 $Y=1.997
+ $X2=4.532 $Y2=2.035
r26 15 16 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=4.532 $Y=2.405
+ $X2=4.532 $Y2=2.775
r27 14 21 0.779116 $w=3.53e-07 $l=2.4e-08 $layer=LI1_cond $X=4.532 $Y=1.973
+ $X2=4.532 $Y2=1.997
r28 14 32 8.1095 $w=3.53e-07 $l=1.53e-07 $layer=LI1_cond $X=4.532 $Y=1.973
+ $X2=4.532 $Y2=1.82
r29 14 15 11.2647 $w=3.53e-07 $l=3.47e-07 $layer=LI1_cond $X=4.532 $Y=2.058
+ $X2=4.532 $Y2=2.405
r30 14 23 0.746653 $w=3.53e-07 $l=2.3e-08 $layer=LI1_cond $X=4.532 $Y=2.058
+ $X2=4.532 $Y2=2.035
r31 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.625 $Y=1.13
+ $X2=4.625 $Y2=1.82
r32 7 13 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=4.532 $Y=0.953
+ $X2=4.532 $Y2=1.13
r33 7 9 14.2189 $w=3.53e-07 $l=4.38e-07 $layer=LI1_cond $X=4.532 $Y=0.953
+ $X2=4.532 $Y2=0.515
r34 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=1.84 $X2=4.52 $Y2=1.985
r35 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=1.84 $X2=4.52 $Y2=2.815
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.38
+ $Y=0.37 $X2=4.52 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A222O_1%VGND 1 2 7 14 24 25 30 36
r43 34 36 10.0102 $w=6.83e-07 $l=1.25e-07 $layer=LI1_cond $X=1.68 $Y=0.257
+ $X2=1.805 $Y2=0.257
r44 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r45 32 34 0.69844 $w=6.83e-07 $l=4e-08 $layer=LI1_cond $X=1.64 $Y=0.257 $X2=1.68
+ $Y2=0.257
r46 29 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r47 28 32 7.68284 $w=6.83e-07 $l=4.4e-07 $layer=LI1_cond $X=1.2 $Y=0.257
+ $X2=1.64 $Y2=0.257
r48 28 30 12.0182 $w=6.83e-07 $l=2.4e-07 $layer=LI1_cond $X=1.2 $Y=0.257
+ $X2=0.96 $Y2=0.257
r49 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r50 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r51 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r52 22 24 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.56
+ $Y2=0
r53 21 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r54 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 18 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r56 17 20 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r57 17 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=1.805
+ $Y2=0
r58 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r59 14 42 10.9023 $w=5.63e-07 $l=5.15e-07 $layer=LI1_cond $X=3.902 $Y=0
+ $X2=3.902 $Y2=0.515
r60 14 22 7.93092 $w=1.7e-07 $l=2.83e-07 $layer=LI1_cond $X=3.902 $Y=0 $X2=4.185
+ $Y2=0
r61 14 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r62 14 20 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.62 $Y=0 $X2=3.6
+ $Y2=0
r63 12 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r64 11 30 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=0.96
+ $Y2=0
r65 11 12 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r66 7 21 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.6
+ $Y2=0
r67 7 18 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r68 2 42 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=3.645
+ $Y=0.37 $X2=3.9 $Y2=0.515
r69 1 32 91 $w=1.7e-07 $l=7.23878e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.37 $X2=1.64 $Y2=0.515
.ends

