# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__inv_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.232000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.350000 2.250000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.172800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 0.350000 0.810000 1.010000 ;
        RECT 0.560000 1.010000 2.680000 1.140000 ;
        RECT 0.560000 1.140000 4.195000 1.180000 ;
        RECT 0.565000 1.950000 2.665000 2.120000 ;
        RECT 0.565000 2.120000 0.815000 2.980000 ;
        RECT 1.500000 0.350000 1.670000 1.010000 ;
        RECT 1.515000 2.120000 1.845000 2.980000 ;
        RECT 2.350000 0.350000 2.680000 1.010000 ;
        RECT 2.420000 1.180000 4.195000 1.310000 ;
        RECT 2.495000 1.310000 4.195000 1.620000 ;
        RECT 2.495000 1.620000 2.665000 1.950000 ;
        RECT 2.495000 2.120000 2.665000 2.980000 ;
        RECT 3.350000 0.350000 3.610000 1.140000 ;
        RECT 3.365000 1.620000 3.695000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.130000  0.085000 0.380000 1.130000 ;
      RECT 0.990000  0.085000 1.320000 0.840000 ;
      RECT 1.015000  2.290000 1.345000 3.245000 ;
      RECT 1.850000  0.085000 2.180000 0.840000 ;
      RECT 2.045000  2.290000 2.295000 3.245000 ;
      RECT 2.850000  0.085000 3.180000 0.970000 ;
      RECT 2.865000  1.820000 3.195000 3.245000 ;
      RECT 3.780000  0.085000 4.110000 0.970000 ;
      RECT 3.865000  1.820000 4.195000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_ls__inv_8
