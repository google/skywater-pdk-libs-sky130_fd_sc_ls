* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__edfxbp_1 CLK D DE VGND VNB VPB VPWR Q Q_N
M1000 VPWR a_575_48# a_2206_443# VPB phighvt w=420000u l=150000u
+  ad=2.56525e+12p pd=2.156e+07u as=1.386e+11p ps=1.5e+06u
M1001 a_1423_508# a_818_74# a_1198_97# VPB phighvt w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=1.26e+11p ps=1.44e+06u
M1002 a_1807_74# a_1419_71# VGND VNB nshort w=740000u l=150000u
+  ad=1.554e+11p pd=1.9e+06u as=1.908e+12p ps=1.641e+07u
M1003 a_1008_74# a_818_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1004 VPWR a_1419_71# a_1423_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_2008_392# a_1419_71# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1006 a_1879_74# a_1008_74# a_1807_74# VNB nshort w=740000u l=150000u
+  ad=7.478e+11p pd=4.66e+06u as=0p ps=0u
M1007 a_27_74# a_575_48# a_556_504# VPB phighvt w=420000u l=150000u
+  ad=4.538e+11p pd=4.78e+06u as=1.008e+11p ps=1.32e+06u
M1008 a_818_74# CLK VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1009 VGND a_575_48# a_2227_118# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1010 a_1198_97# a_1008_74# a_27_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_1879_74# Q VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1012 a_1334_97# a_1008_74# a_1198_97# VNB nshort w=420000u l=150000u
+  ad=1.785e+11p pd=1.69e+06u as=2.226e+11p ps=1.9e+06u
M1013 a_1419_71# a_1198_97# VGND VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1014 a_575_48# a_1879_74# VGND VNB nshort w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1015 VGND a_1879_74# Q VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1016 a_1419_71# a_1198_97# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1017 VGND DE a_145_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1018 a_2206_443# a_1008_74# a_1879_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=3.475e+11p ps=2.84e+06u
M1019 VGND a_1419_71# a_1334_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Q_N a_575_48# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1021 a_1879_74# a_818_74# a_2008_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Q_N a_575_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1023 a_575_48# a_1879_74# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1024 a_116_508# D a_27_74# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1025 a_2227_118# a_818_74# a_1879_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND DE a_161_446# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.281e+11p ps=1.45e+06u
M1027 a_818_74# CLK VGND VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1028 a_1008_74# a_818_74# VGND VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1029 VPWR a_161_446# a_116_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_556_504# DE VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_145_74# D a_27_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=4.158e+11p ps=4.5e+06u
M1032 VPWR DE a_161_446# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1033 a_1198_97# a_818_74# a_27_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_527_74# a_161_446# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1035 a_27_74# a_575_48# a_527_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
