* File: sky130_fd_sc_ls__xnor2_4.pex.spice
* Created: Wed Sep  2 11:30:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__XNOR2_4%A 3 5 7 8 10 13 17 19 21 24 26 28 31 33 35
+ 36 38 40 42 48 50 51 54 57 63 73 86
c180 54 0 1.77085e-19 $X=1.2 $Y=1.665
c181 51 0 2.2033e-19 $X=1.345 $Y=1.665
c182 40 0 9.55446e-20 $X=6.815 $Y=1.765
c183 38 0 3.01101e-20 $X=6.55 $Y=0.74
c184 31 0 3.01101e-20 $X=5.96 $Y=0.74
c185 24 0 3.01105e-20 $X=5.53 $Y=0.74
c186 3 0 7.39126e-20 $X=0.495 $Y=0.69
r187 75 76 37.3828 $w=3.03e-07 $l=2.35e-07 $layer=POLY_cond $X=5.96 $Y=1.557
+ $X2=6.195 $Y2=1.557
r188 74 75 34.2013 $w=3.03e-07 $l=2.15e-07 $layer=POLY_cond $X=5.745 $Y=1.557
+ $X2=5.96 $Y2=1.557
r189 72 74 11.9307 $w=3.03e-07 $l=7.5e-08 $layer=POLY_cond $X=5.67 $Y=1.557
+ $X2=5.745 $Y2=1.557
r190 72 73 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.67
+ $Y=1.515 $X2=5.67 $Y2=1.515
r191 70 72 22.2706 $w=3.03e-07 $l=1.4e-07 $layer=POLY_cond $X=5.53 $Y=1.557
+ $X2=5.67 $Y2=1.557
r192 69 70 65.2211 $w=3.03e-07 $l=4.1e-07 $layer=POLY_cond $X=5.12 $Y=1.557
+ $X2=5.53 $Y2=1.557
r193 68 73 18.4391 $w=4.23e-07 $l=6.8e-07 $layer=LI1_cond $X=4.99 $Y=1.562
+ $X2=5.67 $Y2=1.562
r194 67 69 20.6799 $w=3.03e-07 $l=1.3e-07 $layer=POLY_cond $X=4.99 $Y=1.557
+ $X2=5.12 $Y2=1.557
r195 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.99
+ $Y=1.515 $X2=4.99 $Y2=1.515
r196 65 67 7.9538 $w=3.03e-07 $l=5e-08 $layer=POLY_cond $X=4.94 $Y=1.557
+ $X2=4.99 $Y2=1.557
r197 63 64 4.99482 $w=3.86e-07 $l=4e-08 $layer=POLY_cond $X=0.955 $Y=1.542
+ $X2=0.995 $Y2=1.542
r198 60 61 1.2487 $w=3.86e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.542
+ $X2=0.505 $Y2=1.542
r199 54 86 3.96409 $w=4.58e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.55
+ $X2=1.085 $Y2=1.55
r200 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.665
r201 51 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=1.665
+ $X2=1.2 $Y2=1.665
r202 50 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.415 $Y=1.665
+ $X2=4.56 $Y2=1.665
r203 50 51 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=4.415 $Y=1.665
+ $X2=1.345 $Y2=1.665
r204 48 68 11.66 $w=4.23e-07 $l=4.3e-07 $layer=LI1_cond $X=4.56 $Y=1.562
+ $X2=4.99 $Y2=1.562
r205 48 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=1.665
+ $X2=4.56 $Y2=1.665
r206 46 63 30.5933 $w=3.86e-07 $l=2.45e-07 $layer=POLY_cond $X=0.71 $Y=1.542
+ $X2=0.955 $Y2=1.542
r207 46 61 25.5984 $w=3.86e-07 $l=2.05e-07 $layer=POLY_cond $X=0.71 $Y=1.542
+ $X2=0.505 $Y2=1.542
r208 45 86 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=0.71 $Y=1.485
+ $X2=1.085 $Y2=1.485
r209 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.71
+ $Y=1.485 $X2=0.71 $Y2=1.485
r210 40 42 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.815 $Y=1.765
+ $X2=6.815 $Y2=2.4
r211 36 40 42.1551 $w=3.03e-07 $l=3.54041e-07 $layer=POLY_cond $X=6.55 $Y=1.557
+ $X2=6.815 $Y2=1.765
r212 36 76 56.4719 $w=3.03e-07 $l=3.55e-07 $layer=POLY_cond $X=6.55 $Y=1.557
+ $X2=6.195 $Y2=1.557
r213 36 38 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=6.55 $Y=1.425
+ $X2=6.55 $Y2=0.74
r214 33 76 19.2026 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.195 $Y=1.765
+ $X2=6.195 $Y2=1.557
r215 33 35 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.195 $Y=1.765
+ $X2=6.195 $Y2=2.4
r216 29 75 19.2026 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.96 $Y=1.35
+ $X2=5.96 $Y2=1.557
r217 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.96 $Y=1.35
+ $X2=5.96 $Y2=0.74
r218 26 74 19.2026 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.745 $Y=1.765
+ $X2=5.745 $Y2=1.557
r219 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.745 $Y=1.765
+ $X2=5.745 $Y2=2.4
r220 22 70 19.2026 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.53 $Y=1.35
+ $X2=5.53 $Y2=1.557
r221 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.53 $Y=1.35
+ $X2=5.53 $Y2=0.74
r222 19 69 19.2026 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.12 $Y=1.765
+ $X2=5.12 $Y2=1.557
r223 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.12 $Y=1.765
+ $X2=5.12 $Y2=2.4
r224 15 65 19.2026 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.94 $Y=1.35
+ $X2=4.94 $Y2=1.557
r225 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.94 $Y=1.35
+ $X2=4.94 $Y2=0.74
r226 11 64 24.9932 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.995 $Y=1.32
+ $X2=0.995 $Y2=1.542
r227 11 13 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.995 $Y=1.32
+ $X2=0.995 $Y2=0.69
r228 8 63 24.9932 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.542
r229 8 10 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.26
r230 5 61 24.9932 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.542
r231 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.26
r232 1 60 24.9932 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=1.542
r233 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_4%B 1 3 6 8 10 13 15 17 18 20 23 25 27 30 32
+ 34 35 36 38 39 41 44 46 49 50 51 52 53 54 56 58 59 60 61 70 81
c200 49 0 8.76351e-20 $X=2.07 $Y=1.68
c201 30 0 3.01101e-20 $X=8.035 $Y=0.74
c202 23 0 3.01105e-20 $X=7.605 $Y=0.74
c203 15 0 3.01105e-20 $X=6.98 $Y=1.185
c204 13 0 1.04341e-19 $X=1.925 $Y=0.69
c205 8 0 6.28755e-20 $X=1.855 $Y=1.765
c206 1 0 1.77085e-19 $X=1.405 $Y=1.765
r207 80 81 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.99
+ $Y=1.515 $X2=7.99 $Y2=1.515
r208 78 80 37.8714 $w=3.5e-07 $l=2.75e-07 $layer=POLY_cond $X=7.715 $Y=1.475
+ $X2=7.99 $Y2=1.475
r209 75 76 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.31
+ $Y=1.515 $X2=7.31 $Y2=1.515
r210 73 75 6.19714 $w=3.5e-07 $l=4.5e-08 $layer=POLY_cond $X=7.265 $Y=1.475
+ $X2=7.31 $Y2=1.475
r211 69 70 9.21858 $w=3.66e-07 $l=7e-08 $layer=POLY_cond $X=1.855 $Y=1.557
+ $X2=1.925 $Y2=1.557
r212 68 69 56.6284 $w=3.66e-07 $l=4.3e-07 $layer=POLY_cond $X=1.425 $Y=1.557
+ $X2=1.855 $Y2=1.557
r213 67 68 2.63388 $w=3.66e-07 $l=2e-08 $layer=POLY_cond $X=1.405 $Y=1.557
+ $X2=1.425 $Y2=1.557
r214 61 81 1.94388 $w=4.13e-07 $l=7e-08 $layer=LI1_cond $X=7.92 $Y=1.557
+ $X2=7.99 $Y2=1.557
r215 60 61 13.3295 $w=4.13e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.557
+ $X2=7.92 $Y2=1.557
r216 60 76 3.61006 $w=4.13e-07 $l=1.3e-07 $layer=LI1_cond $X=7.44 $Y=1.557
+ $X2=7.31 $Y2=1.557
r217 59 76 9.7194 $w=4.13e-07 $l=3.5e-07 $layer=LI1_cond $X=6.96 $Y=1.557
+ $X2=7.31 $Y2=1.557
r218 58 84 2.46632 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=6.45 $Y=1.557
+ $X2=6.535 $Y2=1.557
r219 58 59 11.3856 $w=4.13e-07 $l=4.1e-07 $layer=LI1_cond $X=6.55 $Y=1.557
+ $X2=6.96 $Y2=1.557
r220 58 84 0.416546 $w=4.13e-07 $l=1.5e-08 $layer=LI1_cond $X=6.55 $Y=1.557
+ $X2=6.535 $Y2=1.557
r221 57 70 8.56011 $w=3.66e-07 $l=6.5e-08 $layer=POLY_cond $X=1.99 $Y=1.557
+ $X2=1.925 $Y2=1.557
r222 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.99
+ $Y=1.515 $X2=1.99 $Y2=1.515
r223 53 58 6.03523 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=6.45 $Y=1.765
+ $X2=6.45 $Y2=1.557
r224 53 54 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.45 $Y=1.765
+ $X2=6.45 $Y2=1.945
r225 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.365 $Y=2.03
+ $X2=6.45 $Y2=1.945
r226 51 52 274.663 $w=1.68e-07 $l=4.21e-06 $layer=LI1_cond $X=6.365 $Y=2.03
+ $X2=2.155 $Y2=2.03
r227 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.07 $Y=1.945
+ $X2=2.155 $Y2=2.03
r228 49 56 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=1.68
+ $X2=2.07 $Y2=1.515
r229 49 50 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.07 $Y=1.68
+ $X2=2.07 $Y2=1.945
r230 42 46 18.8402 $w=1.65e-07 $l=7.98436e-08 $layer=POLY_cond $X=8.625 $Y=1.35
+ $X2=8.615 $Y2=1.425
r231 42 44 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.625 $Y=1.35
+ $X2=8.625 $Y2=0.74
r232 39 41 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.615 $Y=1.765
+ $X2=8.615 $Y2=2.4
r233 38 39 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.615 $Y=1.675
+ $X2=8.615 $Y2=1.765
r234 37 46 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=8.615 $Y=1.5
+ $X2=8.615 $Y2=1.425
r235 37 38 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=8.615 $Y=1.5
+ $X2=8.615 $Y2=1.675
r236 36 83 28.4554 $w=3.5e-07 $l=1.1225e-07 $layer=POLY_cond $X=8.255 $Y=1.425
+ $X2=8.165 $Y2=1.475
r237 35 46 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.525 $Y=1.425
+ $X2=8.615 $Y2=1.425
r238 35 36 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.525 $Y=1.425
+ $X2=8.255 $Y2=1.425
r239 32 83 22.6286 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.165 $Y=1.765
+ $X2=8.165 $Y2=1.475
r240 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.165 $Y=1.765
+ $X2=8.165 $Y2=2.4
r241 28 83 17.9029 $w=3.5e-07 $l=1.3e-07 $layer=POLY_cond $X=8.035 $Y=1.475
+ $X2=8.165 $Y2=1.475
r242 28 80 6.19714 $w=3.5e-07 $l=4.5e-08 $layer=POLY_cond $X=8.035 $Y=1.475
+ $X2=7.99 $Y2=1.475
r243 28 30 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.035 $Y=1.35
+ $X2=8.035 $Y2=0.74
r244 25 78 22.6286 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.715 $Y=1.765
+ $X2=7.715 $Y2=1.475
r245 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.715 $Y=1.765
+ $X2=7.715 $Y2=2.4
r246 21 78 15.1486 $w=3.5e-07 $l=1.1e-07 $layer=POLY_cond $X=7.605 $Y=1.475
+ $X2=7.715 $Y2=1.475
r247 21 75 40.6257 $w=3.5e-07 $l=2.95e-07 $layer=POLY_cond $X=7.605 $Y=1.475
+ $X2=7.31 $Y2=1.475
r248 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.605 $Y=1.35
+ $X2=7.605 $Y2=0.74
r249 18 73 22.6286 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.265 $Y=1.765
+ $X2=7.265 $Y2=1.475
r250 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.265 $Y=1.765
+ $X2=7.265 $Y2=2.4
r251 15 73 39.2486 $w=3.5e-07 $l=4.0835e-07 $layer=POLY_cond $X=6.98 $Y=1.185
+ $X2=7.265 $Y2=1.475
r252 15 17 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.98 $Y=1.185
+ $X2=6.98 $Y2=0.74
r253 11 70 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=1.557
r254 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=0.69
r255 8 69 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.557
r256 8 10 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.26
r257 4 68 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=1.557
r258 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=0.69
r259 1 67 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.557
r260 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_4%A_116_368# 1 2 3 10 12 15 17 19 22 26 29 30
+ 34 36 37 39 40 43 45 46 48 49 52 55 58 60 61 64 68 78 81
c172 55 0 1.20688e-19 $X=3.92 $Y=1.515
c173 52 0 9.22535e-20 $X=2.48 $Y=1.35
r174 88 89 64.8067 $w=3.57e-07 $l=4.8e-07 $layer=POLY_cond $X=2.935 $Y=1.557
+ $X2=3.415 $Y2=1.557
r175 87 88 2.70028 $w=3.57e-07 $l=2e-08 $layer=POLY_cond $X=2.915 $Y=1.557
+ $X2=2.935 $Y2=1.557
r176 81 89 10.4808 $w=3.57e-07 $l=9.3675e-08 $layer=POLY_cond $X=3.49 $Y=1.515
+ $X2=3.415 $Y2=1.557
r177 76 78 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=2.79
+ $X2=3.58 $Y2=2.79
r178 76 77 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.745
+ $Y=2.79 $X2=3.745 $Y2=2.79
r179 74 87 47.93 $w=3.57e-07 $l=3.55e-07 $layer=POLY_cond $X=2.56 $Y=1.557
+ $X2=2.915 $Y2=1.557
r180 74 85 10.126 $w=3.57e-07 $l=7.5e-08 $layer=POLY_cond $X=2.56 $Y=1.557
+ $X2=2.485 $Y2=1.557
r181 73 74 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.56
+ $Y=1.515 $X2=2.56 $Y2=1.515
r182 68 70 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.71 $Y=0.86
+ $X2=1.71 $Y2=1.095
r183 60 61 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.425
+ $Y=2.79 $X2=4.425 $Y2=2.79
r184 58 76 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.91 $Y=2.79
+ $X2=3.745 $Y2=2.79
r185 58 60 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=3.91 $Y=2.79
+ $X2=4.425 $Y2=2.79
r186 56 81 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.92 $Y=1.515
+ $X2=3.49 $Y2=1.515
r187 55 56 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.92
+ $Y=1.515 $X2=3.92 $Y2=1.515
r188 53 73 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=1.515
+ $X2=2.48 $Y2=1.515
r189 53 55 47.32 $w=3.28e-07 $l=1.355e-06 $layer=LI1_cond $X=2.565 $Y=1.515
+ $X2=3.92 $Y2=1.515
r190 52 73 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=1.35
+ $X2=2.48 $Y2=1.515
r191 51 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.48 $Y=1.18
+ $X2=2.48 $Y2=1.35
r192 50 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=1.095
+ $X2=1.71 $Y2=1.095
r193 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.395 $Y=1.095
+ $X2=2.48 $Y2=1.18
r194 49 50 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.395 $Y=1.095
+ $X2=1.875 $Y2=1.095
r195 48 78 116.455 $w=1.68e-07 $l=1.785e-06 $layer=LI1_cond $X=1.795 $Y=2.71
+ $X2=3.58 $Y2=2.71
r196 46 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.63 $Y=2.625
+ $X2=1.795 $Y2=2.71
r197 45 66 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=2.12 $X2=1.63
+ $Y2=2.035
r198 45 46 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=1.63 $Y=2.12
+ $X2=1.63 $Y2=2.625
r199 44 64 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=0.895 $Y=2.035
+ $X2=0.73 $Y2=1.97
r200 43 66 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=1.63 $Y2=2.035
r201 43 44 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=0.895 $Y2=2.035
r202 39 77 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.935 $Y=2.79
+ $X2=3.745 $Y2=2.79
r203 39 40 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.935 $Y=2.79
+ $X2=4.01 $Y2=2.79
r204 38 61 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.085 $Y=2.79
+ $X2=4.425 $Y2=2.79
r205 38 40 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.085 $Y=2.79
+ $X2=4.01 $Y2=2.79
r206 36 56 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.935 $Y=1.515
+ $X2=3.92 $Y2=1.515
r207 36 37 6.91837 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.935 $Y=1.515
+ $X2=4.01 $Y2=1.515
r208 32 34 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.44 $Y=1.35
+ $X2=4.44 $Y2=0.74
r209 31 37 6.91837 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.085 $Y=1.425
+ $X2=4.01 $Y2=1.515
r210 30 32 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.365 $Y=1.425
+ $X2=4.44 $Y2=1.35
r211 30 31 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.365 $Y=1.425
+ $X2=4.085 $Y2=1.425
r212 29 40 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.01 $Y=2.625
+ $X2=4.01 $Y2=2.79
r213 28 37 18.1359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.01 $Y=1.68
+ $X2=4.01 $Y2=1.515
r214 28 29 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=4.01 $Y=1.68
+ $X2=4.01 $Y2=2.625
r215 24 37 18.1359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.01 $Y=1.35
+ $X2=4.01 $Y2=1.515
r216 24 26 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.01 $Y=1.35
+ $X2=4.01 $Y2=0.74
r217 20 89 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.415 $Y=1.35
+ $X2=3.415 $Y2=1.557
r218 20 22 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.415 $Y=1.35
+ $X2=3.415 $Y2=0.74
r219 17 88 23.1043 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.935 $Y=1.765
+ $X2=2.935 $Y2=1.557
r220 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.935 $Y=1.765
+ $X2=2.935 $Y2=2.4
r221 13 87 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.915 $Y=1.35
+ $X2=2.915 $Y2=1.557
r222 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.915 $Y=1.35
+ $X2=2.915 $Y2=0.74
r223 10 85 23.1043 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.485 $Y=1.765
+ $X2=2.485 $Y2=1.557
r224 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.485 $Y=1.765
+ $X2=2.485 $Y2=2.4
r225 3 66 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.115
r226 2 64 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r227 1 68 182 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.71 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_4%VPWR 1 2 3 4 5 6 19 21 25 27 30 31 33 36 39
+ 45 56 65 66 72 79 86
r112 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r113 86 89 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.505 $Y=3.05
+ $X2=6.505 $Y2=3.33
r114 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r115 79 82 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.245 $Y=3.05
+ $X2=3.245 $Y2=3.33
r116 76 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r117 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r118 72 75 9.49071 $w=3.38e-07 $l=2.8e-07 $layer=LI1_cond $X=2.17 $Y=3.05
+ $X2=2.17 $Y2=3.33
r119 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r120 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r121 63 66 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r122 63 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r123 62 65 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r124 62 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r125 60 89 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.67 $Y=3.33
+ $X2=6.505 $Y2=3.33
r126 60 62 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.67 $Y=3.33
+ $X2=6.96 $Y2=3.33
r127 59 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r128 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r129 56 89 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.34 $Y=3.33
+ $X2=6.505 $Y2=3.33
r130 56 58 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.34 $Y=3.33 $X2=6
+ $Y2=3.33
r131 55 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r132 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r133 52 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r134 51 54 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r135 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r136 49 82 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.41 $Y=3.33
+ $X2=3.245 $Y2=3.33
r137 49 51 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.41 $Y=3.33
+ $X2=3.6 $Y2=3.33
r138 48 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r139 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r140 45 75 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2 $Y=3.33 $X2=2.17
+ $Y2=3.33
r141 45 47 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2 $Y=3.33 $X2=1.68
+ $Y2=3.33
r142 44 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r143 44 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r144 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r145 41 69 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r146 41 43 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r147 39 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r148 39 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.6 $Y2=3.33
r149 37 58 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.6 $Y=3.33 $X2=6
+ $Y2=3.33
r150 36 54 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.265 $Y=3.33
+ $X2=5.04 $Y2=3.33
r151 36 37 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=5.432 $Y=3.33
+ $X2=5.6 $Y2=3.33
r152 33 36 9.63236 $w=3.33e-07 $l=2.8e-07 $layer=LI1_cond $X=5.432 $Y=3.05
+ $X2=5.432 $Y2=3.33
r153 30 43 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r154 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.18 $Y2=3.33
r155 29 47 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r156 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.18 $Y2=3.33
r157 28 75 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.34 $Y=3.33
+ $X2=2.17 $Y2=3.33
r158 27 82 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=3.33
+ $X2=3.245 $Y2=3.33
r159 27 28 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.08 $Y=3.33
+ $X2=2.34 $Y2=3.33
r160 23 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r161 23 25 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.495
r162 19 69 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r163 19 21 58.0831 $w=2.48e-07 $l=1.26e-06 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=1.985
r164 6 86 600 $w=1.7e-07 $l=1.32229e-06 $layer=licon1_PDIFF $count=1 $X=6.27
+ $Y=1.84 $X2=6.505 $Y2=3.05
r165 5 33 600 $w=1.7e-07 $l=1.32229e-06 $layer=licon1_PDIFF $count=1 $X=5.195
+ $Y=1.84 $X2=5.43 $Y2=3.05
r166 4 79 600 $w=1.7e-07 $l=1.32229e-06 $layer=licon1_PDIFF $count=1 $X=3.01
+ $Y=1.84 $X2=3.245 $Y2=3.05
r167 3 72 600 $w=1.7e-07 $l=1.32458e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.17 $Y2=3.05
r168 2 25 600 $w=1.7e-07 $l=7.26137e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.495
r169 1 21 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_4%Y 1 2 3 4 5 16 22 24 25 28 30 32 37 38 41 42
+ 45
r133 42 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.49 $Y=2.02 $X2=7.49
+ $Y2=2.105
r134 42 45 0.244458 $w=3.28e-07 $l=7e-09 $layer=LI1_cond $X=7.49 $Y=2.112
+ $X2=7.49 $Y2=2.105
r135 39 42 6.04159 $w=3.28e-07 $l=1.73e-07 $layer=LI1_cond $X=7.49 $Y=2.285
+ $X2=7.49 $Y2=2.112
r136 37 41 3.70735 $w=2.5e-07 $l=9.44722e-08 $layer=LI1_cond $X=8.41 $Y=1.935
+ $X2=8.39 $Y2=2.02
r137 36 37 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=8.41 $Y=1.18
+ $X2=8.41 $Y2=1.935
r138 33 42 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.655 $Y=2.02
+ $X2=7.49 $Y2=2.02
r139 32 41 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.225 $Y=2.02
+ $X2=8.39 $Y2=2.02
r140 32 33 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.225 $Y=2.02
+ $X2=7.655 $Y2=2.02
r141 31 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.39 $Y=1.095
+ $X2=4.225 $Y2=1.095
r142 30 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.325 $Y=1.095
+ $X2=8.41 $Y2=1.18
r143 30 31 256.722 $w=1.68e-07 $l=3.935e-06 $layer=LI1_cond $X=8.325 $Y=1.095
+ $X2=4.39 $Y2=1.095
r144 26 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=1.01
+ $X2=4.225 $Y2=1.095
r145 26 28 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.225 $Y=1.01
+ $X2=4.225 $Y2=0.86
r146 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=1.095
+ $X2=4.225 $Y2=1.095
r147 24 25 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.06 $Y=1.095
+ $X2=3.365 $Y2=1.095
r148 20 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.2 $Y=1.01
+ $X2=3.365 $Y2=1.095
r149 20 22 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.2 $Y=1.01 $X2=3.2
+ $Y2=0.86
r150 16 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.325 $Y=2.37
+ $X2=7.49 $Y2=2.285
r151 16 18 301.086 $w=1.68e-07 $l=4.615e-06 $layer=LI1_cond $X=7.325 $Y=2.37
+ $X2=2.71 $Y2=2.37
r152 5 41 300 $w=1.7e-07 $l=3.26497e-07 $layer=licon1_PDIFF $count=2 $X=8.24
+ $Y=1.84 $X2=8.39 $Y2=2.1
r153 4 42 300 $w=1.7e-07 $l=3.26497e-07 $layer=licon1_PDIFF $count=2 $X=7.34
+ $Y=1.84 $X2=7.49 $Y2=2.1
r154 3 18 600 $w=1.7e-07 $l=6.00333e-07 $layer=licon1_PDIFF $count=1 $X=2.56
+ $Y=1.84 $X2=2.71 $Y2=2.37
r155 2 28 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=4.085
+ $Y=0.37 $X2=4.225 $Y2=0.86
r156 1 22 182 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=1 $X=2.99
+ $Y=0.37 $X2=3.2 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_4%A_950_368# 1 2 3 4 5 18 20 24 26 30 34 41 42
+ 43 49
c70 20 0 9.55446e-20 $X=7.855 $Y=2.99
r71 46 47 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=7 $Y=2.8 $X2=7
+ $Y2=2.99
r72 43 46 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=7 $Y=2.71 $X2=7
+ $Y2=2.8
r73 40 42 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=5.97 $Y=2.802
+ $X2=6.135 $Y2=2.802
r74 40 41 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=5.97 $Y=2.802
+ $X2=5.805 $Y2=2.802
r75 34 37 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.935 $Y=2.71
+ $X2=4.935 $Y2=2.8
r76 30 33 32.9599 $w=2.48e-07 $l=7.15e-07 $layer=LI1_cond $X=8.88 $Y=2.1
+ $X2=8.88 $Y2=2.815
r77 28 33 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=8.88 $Y=2.905 $X2=8.88
+ $Y2=2.815
r78 27 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.025 $Y=2.99
+ $X2=7.94 $Y2=2.99
r79 26 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.755 $Y=2.99
+ $X2=8.88 $Y2=2.905
r80 26 27 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=8.755 $Y=2.99
+ $X2=8.025 $Y2=2.99
r81 22 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.94 $Y=2.905
+ $X2=7.94 $Y2=2.99
r82 22 24 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=7.94 $Y=2.905
+ $X2=7.94 $Y2=2.44
r83 21 47 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.125 $Y=2.99 $X2=7
+ $Y2=2.99
r84 20 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.855 $Y=2.99
+ $X2=7.94 $Y2=2.99
r85 20 21 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.855 $Y=2.99
+ $X2=7.125 $Y2=2.99
r86 18 43 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.875 $Y=2.71 $X2=7
+ $Y2=2.71
r87 18 42 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.875 $Y=2.71
+ $X2=6.135 $Y2=2.71
r88 17 34 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.06 $Y=2.71
+ $X2=4.935 $Y2=2.71
r89 17 41 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=5.06 $Y=2.71
+ $X2=5.805 $Y2=2.71
r90 5 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.69
+ $Y=1.84 $X2=8.84 $Y2=2.815
r91 5 30 400 $w=1.7e-07 $l=3.26497e-07 $layer=licon1_PDIFF $count=1 $X=8.69
+ $Y=1.84 $X2=8.84 $Y2=2.1
r92 4 24 300 $w=1.7e-07 $l=6.7082e-07 $layer=licon1_PDIFF $count=2 $X=7.79
+ $Y=1.84 $X2=7.94 $Y2=2.44
r93 3 46 600 $w=1.7e-07 $l=1.03228e-06 $layer=licon1_PDIFF $count=1 $X=6.89
+ $Y=1.84 $X2=7.04 $Y2=2.8
r94 2 40 600 $w=1.7e-07 $l=1.03228e-06 $layer=licon1_PDIFF $count=1 $X=5.82
+ $Y=1.84 $X2=5.97 $Y2=2.8
r95 1 37 600 $w=1.7e-07 $l=1.02995e-06 $layer=licon1_PDIFF $count=1 $X=4.75
+ $Y=1.84 $X2=4.895 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_4%A_27_74# 1 2 3 12 14 15 16 17 20
c40 16 0 7.39126e-20 $X=1.21 $Y=0.6
c41 14 0 1.04341e-19 $X=1.045 $Y=1.065
r42 18 23 3.97509 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.475
+ $X2=1.21 $Y2=0.475
r43 18 20 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=1.375 $Y=0.475
+ $X2=2.14 $Y2=0.475
r44 16 23 3.01144 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=1.21 $Y=0.6 $X2=1.21
+ $Y2=0.475
r45 16 17 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.21 $Y=0.6 $X2=1.21
+ $Y2=0.98
r46 14 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.045 $Y=1.065
+ $X2=1.21 $Y2=0.98
r47 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=1.065
+ $X2=0.365 $Y2=1.065
r48 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.98
+ $X2=0.365 $Y2=1.065
r49 10 12 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=0.24 $Y=0.98
+ $X2=0.24 $Y2=0.515
r50 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2 $Y=0.37
+ $X2=2.14 $Y2=0.515
r51 2 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.515
r52 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_4%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41 43
+ 44 45 47 65 71 72 75 78
r117 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r118 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r119 72 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r120 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r121 69 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.495 $Y=0 $X2=8.33
+ $Y2=0
r122 69 71 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.495 $Y=0
+ $X2=8.88 $Y2=0
r123 68 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r124 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r125 65 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.165 $Y=0 $X2=8.33
+ $Y2=0
r126 65 67 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=8.165 $Y=0 $X2=7.92
+ $Y2=0
r127 64 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r128 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r129 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r130 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r131 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r132 57 58 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r133 55 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r134 54 57 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=5.04
+ $Y2=0
r135 54 55 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r136 52 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r137 52 54 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r138 50 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r139 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r140 47 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r141 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r142 45 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r143 45 55 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=1.2
+ $Y2=0
r144 43 63 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.11 $Y=0 $X2=6.96
+ $Y2=0
r145 43 44 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=7.11 $Y=0 $X2=7.292
+ $Y2=0
r146 42 67 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=7.475 $Y=0
+ $X2=7.92 $Y2=0
r147 42 44 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=7.475 $Y=0
+ $X2=7.292 $Y2=0
r148 40 60 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.09 $Y=0 $X2=6 $Y2=0
r149 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.09 $Y=0 $X2=6.255
+ $Y2=0
r150 39 63 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=6.42 $Y=0 $X2=6.96
+ $Y2=0
r151 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.42 $Y=0 $X2=6.255
+ $Y2=0
r152 37 57 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=5.07 $Y=0 $X2=5.04
+ $Y2=0
r153 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.07 $Y=0 $X2=5.235
+ $Y2=0
r154 36 60 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.4 $Y=0 $X2=6 $Y2=0
r155 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.4 $Y=0 $X2=5.235
+ $Y2=0
r156 32 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.33 $Y=0.085
+ $X2=8.33 $Y2=0
r157 32 34 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=8.33 $Y=0.085
+ $X2=8.33 $Y2=0.335
r158 28 44 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=7.292 $Y=0.085
+ $X2=7.292 $Y2=0
r159 28 30 7.89345 $w=3.63e-07 $l=2.5e-07 $layer=LI1_cond $X=7.292 $Y=0.085
+ $X2=7.292 $Y2=0.335
r160 24 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.255 $Y=0.085
+ $X2=6.255 $Y2=0
r161 24 26 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6.255 $Y=0.085
+ $X2=6.255 $Y2=0.335
r162 20 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.235 $Y=0.085
+ $X2=5.235 $Y2=0
r163 20 22 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=5.235 $Y=0.085
+ $X2=5.235 $Y2=0.335
r164 16 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r165 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.58
r166 5 34 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=8.11
+ $Y=0.37 $X2=8.33 $Y2=0.335
r167 4 30 182 $w=1.7e-07 $l=2.51893e-07 $layer=licon1_NDIFF $count=1 $X=7.055
+ $Y=0.37 $X2=7.29 $Y2=0.335
r168 3 26 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=6.035
+ $Y=0.37 $X2=6.255 $Y2=0.335
r169 2 22 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=5.015
+ $Y=0.37 $X2=5.235 $Y2=0.335
r170 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__XNOR2_4%A_511_74# 1 2 3 4 5 6 7 24 26 27 30 32 37 38
+ 39 40 42 44 46 48 53 58 63
c121 44 0 3.01105e-20 $X=8.675 $Y=0.755
c122 42 0 6.02202e-20 $X=7.655 $Y=0.755
c123 40 0 6.0221e-20 $X=6.6 $Y=0.755
c124 38 0 3.01101e-20 $X=5.58 $Y=0.755
r125 63 65 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=8.84 $Y=0.515
+ $X2=8.84 $Y2=0.755
r126 58 60 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=7.82 $Y=0.595
+ $X2=7.82 $Y2=0.755
r127 53 55 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=6.765 $Y=0.595
+ $X2=6.765 $Y2=0.755
r128 48 50 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=5.745 $Y=0.595
+ $X2=5.745 $Y2=0.755
r129 45 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.985 $Y=0.755
+ $X2=7.82 $Y2=0.755
r130 44 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.675 $Y=0.755
+ $X2=8.84 $Y2=0.755
r131 44 45 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.675 $Y=0.755
+ $X2=7.985 $Y2=0.755
r132 43 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.93 $Y=0.755
+ $X2=6.765 $Y2=0.755
r133 42 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.655 $Y=0.755
+ $X2=7.82 $Y2=0.755
r134 42 43 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.655 $Y=0.755
+ $X2=6.93 $Y2=0.755
r135 41 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.91 $Y=0.755
+ $X2=5.745 $Y2=0.755
r136 40 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.6 $Y=0.755
+ $X2=6.765 $Y2=0.755
r137 40 41 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.6 $Y=0.755
+ $X2=5.91 $Y2=0.755
r138 38 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.58 $Y=0.755
+ $X2=5.745 $Y2=0.755
r139 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.58 $Y=0.755
+ $X2=4.89 $Y2=0.755
r140 35 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.725 $Y=0.67
+ $X2=4.89 $Y2=0.755
r141 35 37 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=4.725 $Y=0.67
+ $X2=4.725 $Y2=0.595
r142 34 37 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.725 $Y=0.425
+ $X2=4.725 $Y2=0.595
r143 33 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.865 $Y=0.34
+ $X2=3.7 $Y2=0.34
r144 32 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.56 $Y=0.34
+ $X2=4.725 $Y2=0.425
r145 32 33 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.56 $Y=0.34
+ $X2=3.865 $Y2=0.34
r146 28 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.425 $X2=3.7
+ $Y2=0.34
r147 28 30 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.7 $Y=0.425
+ $X2=3.7 $Y2=0.595
r148 26 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.535 $Y=0.34
+ $X2=3.7 $Y2=0.34
r149 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.535 $Y=0.34
+ $X2=2.865 $Y2=0.34
r150 22 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.7 $Y=0.425
+ $X2=2.865 $Y2=0.34
r151 22 24 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.7 $Y=0.425
+ $X2=2.7 $Y2=0.595
r152 7 63 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.37 $X2=8.84 $Y2=0.515
r153 6 58 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=7.68
+ $Y=0.37 $X2=7.82 $Y2=0.595
r154 5 53 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=6.625
+ $Y=0.37 $X2=6.765 $Y2=0.595
r155 4 48 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=5.605
+ $Y=0.37 $X2=5.745 $Y2=0.595
r156 3 37 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=4.515
+ $Y=0.37 $X2=4.725 $Y2=0.595
r157 2 30 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=3.49
+ $Y=0.37 $X2=3.7 $Y2=0.595
r158 1 24 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.37 $X2=2.7 $Y2=0.595
.ends

