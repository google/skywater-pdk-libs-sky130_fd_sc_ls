* File: sky130_fd_sc_ls__dlygate4sd1_1.spice
* Created: Wed Sep  2 11:05:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dlygate4sd1_1.pex.spice"
.subckt sky130_fd_sc_ls__dlygate4sd1_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_28_74#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.15435 AS=0.1113 PD=1.155 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_A_286_392#_M1007_d N_A_28_74#_M1007_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.15435 PD=1.37 PS=1.155 NRD=0 NRS=114.276 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_286_392#_M1001_g N_A_405_138#_M1001_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0831672 AS=0.2562 PD=0.78569 PS=2.06 NRD=40.86 NRS=41.424
+ M=1 R=2.8 SA=75000.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_405_138#_M1006_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.146533 PD=2.01 PS=1.38431 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_28_74#_M1002_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.188556 AS=0.1176 PD=1.01155 PS=1.4 NRD=14.0658 NRS=7.0329 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_A_286_392#_M1000_d N_A_28_74#_M1000_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=1 AD=0.275 AS=0.448944 PD=2.55 PS=2.40845 NRD=1.9503 NRS=78.7803 M=1
+ R=6.66667 SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A_286_392#_M1004_g N_A_405_138#_M1004_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.190094 AS=0.595 PD=1.40566 PS=3.19 NRD=16.2328 NRS=65.01 M=1
+ R=6.66667 SA=75000.5 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1003 N_X_M1003_d N_A_405_138#_M1003_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3136 AS=0.212906 PD=2.8 PS=1.57434 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75000.9 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ls__dlygate4sd1_1.pxi.spice"
*
.ends
*
*
