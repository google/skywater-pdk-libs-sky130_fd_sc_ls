* File: sky130_fd_sc_ls__or2_1.pxi.spice
* Created: Wed Sep  2 11:24:04 2020
* 
x_PM_SKY130_FD_SC_LS__OR2_1%B N_B_c_41_n N_B_c_45_n N_B_M1000_g N_B_M1004_g B
+ N_B_c_42_n N_B_c_43_n PM_SKY130_FD_SC_LS__OR2_1%B
x_PM_SKY130_FD_SC_LS__OR2_1%A N_A_c_68_n N_A_M1005_g N_A_M1003_g A N_A_c_70_n
+ PM_SKY130_FD_SC_LS__OR2_1%A
x_PM_SKY130_FD_SC_LS__OR2_1%A_63_368# N_A_63_368#_M1004_d N_A_63_368#_M1000_s
+ N_A_63_368#_c_104_n N_A_63_368#_M1002_g N_A_63_368#_M1001_g
+ N_A_63_368#_c_114_n N_A_63_368#_c_106_n N_A_63_368#_c_107_n
+ N_A_63_368#_c_108_n N_A_63_368#_c_109_n N_A_63_368#_c_110_n
+ N_A_63_368#_c_113_n PM_SKY130_FD_SC_LS__OR2_1%A_63_368#
x_PM_SKY130_FD_SC_LS__OR2_1%VPWR N_VPWR_M1005_d N_VPWR_c_173_n VPWR
+ N_VPWR_c_174_n N_VPWR_c_175_n N_VPWR_c_172_n N_VPWR_c_177_n
+ PM_SKY130_FD_SC_LS__OR2_1%VPWR
x_PM_SKY130_FD_SC_LS__OR2_1%X N_X_M1001_d N_X_M1002_d N_X_c_196_n N_X_c_197_n X
+ X X X N_X_c_198_n PM_SKY130_FD_SC_LS__OR2_1%X
x_PM_SKY130_FD_SC_LS__OR2_1%VGND N_VGND_M1004_s N_VGND_M1003_d N_VGND_c_221_n
+ N_VGND_c_222_n N_VGND_c_223_n N_VGND_c_224_n VGND N_VGND_c_225_n
+ N_VGND_c_226_n N_VGND_c_227_n N_VGND_c_228_n PM_SKY130_FD_SC_LS__OR2_1%VGND
cc_1 VNB N_B_c_41_n 0.0794593f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.385
cc_2 VNB N_B_c_42_n 0.0221254f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.22
cc_3 VNB N_B_c_43_n 0.0293162f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_4 VNB N_A_c_68_n 0.0302615f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.385
cc_5 VNB N_A_M1003_g 0.027266f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_6 VNB N_A_c_70_n 0.00189714f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.22
cc_7 VNB N_A_63_368#_c_104_n 0.0360092f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.835
cc_8 VNB N_A_63_368#_M1001_g 0.0286452f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.22
cc_9 VNB N_A_63_368#_c_106_n 0.0038832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_63_368#_c_107_n 0.00741821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_63_368#_c_108_n 0.00541617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_63_368#_c_109_n 0.00770034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_63_368#_c_110_n 4.1382e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_172_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.365
cc_15 VNB N_X_c_196_n 0.0265168f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB N_X_c_197_n 0.0133911f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_17 VNB N_X_c_198_n 0.0246503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_221_n 0.0267471f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_19 VNB N_VGND_c_222_n 0.0168543f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_20 VNB N_VGND_c_223_n 0.0115308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_224_n 0.00682834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_225_n 0.0239783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_226_n 0.0189562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_227_n 0.177517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_228_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VPB N_B_c_41_n 0.00964707f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.385
cc_27 VPB N_B_c_45_n 0.0206185f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=1.765
cc_28 VPB N_A_c_68_n 0.0301014f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.385
cc_29 VPB N_A_c_70_n 0.00259191f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=1.22
cc_30 VPB N_A_63_368#_c_104_n 0.0301784f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=0.835
cc_31 VPB N_A_63_368#_c_110_n 0.00318732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_A_63_368#_c_113_n 0.0406471f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_173_n 0.022626f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.22
cc_34 VPB N_VPWR_c_174_n 0.0377411f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_175_n 0.0189562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_172_n 0.0756276f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.365
cc_37 VPB N_VPWR_c_177_n 0.0118997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB X 0.0135031f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_39 VPB X 0.0415177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_X_c_198_n 0.00755527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 N_B_c_41_n N_A_c_68_n 0.0215463f $X=0.595 $Y=1.385 $X2=-0.19 $Y2=-0.245
cc_42 N_B_c_45_n N_A_c_68_n 0.0476034f $X=0.685 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_43 N_B_c_43_n N_A_c_68_n 7.73509e-19 $X=0.61 $Y=1.385 $X2=-0.19 $Y2=-0.245
cc_44 N_B_c_42_n N_A_M1003_g 0.0135545f $X=0.685 $Y=1.22 $X2=0 $Y2=0
cc_45 N_B_c_43_n N_A_M1003_g 9.09937e-19 $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_46 N_B_c_41_n N_A_c_70_n 0.00158099f $X=0.595 $Y=1.385 $X2=0 $Y2=0
cc_47 N_B_c_43_n N_A_c_70_n 0.0109438f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_48 N_B_c_45_n N_A_63_368#_c_114_n 0.0128795f $X=0.685 $Y=1.765 $X2=0 $Y2=0
cc_49 N_B_c_43_n N_A_63_368#_c_114_n 0.00515375f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_50 N_B_c_42_n N_A_63_368#_c_106_n 0.00461704f $X=0.685 $Y=1.22 $X2=0 $Y2=0
cc_51 N_B_c_42_n N_A_63_368#_c_108_n 0.00500991f $X=0.685 $Y=1.22 $X2=0 $Y2=0
cc_52 N_B_c_41_n N_A_63_368#_c_113_n 0.00706476f $X=0.595 $Y=1.385 $X2=0 $Y2=0
cc_53 N_B_c_45_n N_A_63_368#_c_113_n 0.0169085f $X=0.685 $Y=1.765 $X2=0 $Y2=0
cc_54 N_B_c_43_n N_A_63_368#_c_113_n 0.0197713f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_55 N_B_c_45_n N_VPWR_c_173_n 0.00170182f $X=0.685 $Y=1.765 $X2=0 $Y2=0
cc_56 N_B_c_45_n N_VPWR_c_174_n 0.00393873f $X=0.685 $Y=1.765 $X2=0 $Y2=0
cc_57 N_B_c_45_n N_VPWR_c_172_n 0.00462577f $X=0.685 $Y=1.765 $X2=0 $Y2=0
cc_58 N_B_c_41_n N_VGND_c_221_n 0.00215345f $X=0.595 $Y=1.385 $X2=0 $Y2=0
cc_59 N_B_c_42_n N_VGND_c_221_n 0.0135644f $X=0.685 $Y=1.22 $X2=0 $Y2=0
cc_60 N_B_c_43_n N_VGND_c_221_n 0.0264066f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_61 N_B_c_42_n N_VGND_c_225_n 0.00375057f $X=0.685 $Y=1.22 $X2=0 $Y2=0
cc_62 N_B_c_42_n N_VGND_c_227_n 0.00409726f $X=0.685 $Y=1.22 $X2=0 $Y2=0
cc_63 N_A_c_68_n N_A_63_368#_c_104_n 0.00972422f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_64 N_A_M1003_g N_A_63_368#_c_104_n 0.0174761f $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_65 N_A_c_70_n N_A_63_368#_c_104_n 3.285e-19 $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_66 N_A_M1003_g N_A_63_368#_M1001_g 0.0176009f $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_67 N_A_c_68_n N_A_63_368#_c_114_n 0.0180645f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_68 N_A_c_70_n N_A_63_368#_c_114_n 0.0232724f $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_69 N_A_M1003_g N_A_63_368#_c_106_n 6.93808e-19 $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_70 N_A_M1003_g N_A_63_368#_c_107_n 0.0162525f $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_71 N_A_c_70_n N_A_63_368#_c_107_n 0.00982684f $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_72 N_A_c_68_n N_A_63_368#_c_108_n 0.00262205f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A_c_70_n N_A_63_368#_c_108_n 0.0166608f $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_74 N_A_M1003_g N_A_63_368#_c_109_n 0.00546476f $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_75 N_A_c_70_n N_A_63_368#_c_109_n 0.0172973f $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_76 N_A_c_68_n N_A_63_368#_c_110_n 0.00360163f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_77 N_A_c_70_n N_A_63_368#_c_110_n 0.00910638f $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_78 N_A_c_68_n N_A_63_368#_c_113_n 0.00262311f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_79 N_A_c_68_n N_VPWR_c_173_n 0.0141899f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A_c_68_n N_VPWR_c_174_n 0.00361294f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A_c_68_n N_VPWR_c_172_n 0.00419404f $X=1.105 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_M1003_g N_X_c_196_n 8.51118e-19 $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_83 N_A_M1003_g N_VGND_c_221_n 6.19635e-19 $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_84 N_A_M1003_g N_VGND_c_222_n 0.00508306f $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_85 N_A_M1003_g N_VGND_c_225_n 0.00451272f $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_86 N_A_M1003_g N_VGND_c_227_n 0.00487769f $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_87 N_A_63_368#_c_114_n A_152_368# 0.0119045f $X=1.615 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_88 N_A_63_368#_c_114_n N_VPWR_M1005_d 0.0190678f $X=1.615 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_89 N_A_63_368#_c_110_n N_VPWR_M1005_d 0.00247124f $X=1.7 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_90 N_A_63_368#_c_104_n N_VPWR_c_173_n 0.00595709f $X=1.895 $Y=1.765 $X2=0
+ $Y2=0
cc_91 N_A_63_368#_c_114_n N_VPWR_c_173_n 0.0450402f $X=1.615 $Y=2.035 $X2=0
+ $Y2=0
cc_92 N_A_63_368#_c_113_n N_VPWR_c_173_n 0.0125263f $X=0.46 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A_63_368#_c_113_n N_VPWR_c_174_n 0.0066794f $X=0.46 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A_63_368#_c_104_n N_VPWR_c_175_n 0.00445602f $X=1.895 $Y=1.765 $X2=0
+ $Y2=0
cc_95 N_A_63_368#_c_104_n N_VPWR_c_172_n 0.00865213f $X=1.895 $Y=1.765 $X2=0
+ $Y2=0
cc_96 N_A_63_368#_c_113_n N_VPWR_c_172_n 0.00997343f $X=0.46 $Y=1.985 $X2=0
+ $Y2=0
cc_97 N_A_63_368#_M1001_g N_X_c_196_n 0.00926861f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_98 N_A_63_368#_c_104_n N_X_c_197_n 2.30445e-19 $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_63_368#_M1001_g N_X_c_197_n 0.00349857f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A_63_368#_c_109_n N_X_c_197_n 0.00658407f $X=1.7 $Y=1.63 $X2=0 $Y2=0
cc_101 N_A_63_368#_c_104_n X 0.00318178f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_63_368#_c_109_n X 0.00102654f $X=1.7 $Y=1.63 $X2=0 $Y2=0
cc_103 N_A_63_368#_c_110_n X 0.00564758f $X=1.7 $Y=1.95 $X2=0 $Y2=0
cc_104 N_A_63_368#_c_104_n X 0.01695f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A_63_368#_c_104_n N_X_c_198_n 0.0106907f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_106 N_A_63_368#_M1001_g N_X_c_198_n 0.00255066f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_63_368#_c_109_n N_X_c_198_n 0.0304892f $X=1.7 $Y=1.63 $X2=0 $Y2=0
cc_108 N_A_63_368#_c_110_n N_X_c_198_n 0.00628995f $X=1.7 $Y=1.95 $X2=0 $Y2=0
cc_109 N_A_63_368#_c_107_n N_VGND_M1003_d 0.00185525f $X=1.615 $Y=1.095 $X2=0
+ $Y2=0
cc_110 N_A_63_368#_c_109_n N_VGND_M1003_d 0.002623f $X=1.7 $Y=1.63 $X2=0 $Y2=0
cc_111 N_A_63_368#_c_106_n N_VGND_c_221_n 0.0231039f $X=1.075 $Y=0.82 $X2=0
+ $Y2=0
cc_112 N_A_63_368#_c_104_n N_VGND_c_222_n 5.87857e-19 $X=1.895 $Y=1.765 $X2=0
+ $Y2=0
cc_113 N_A_63_368#_M1001_g N_VGND_c_222_n 0.00879154f $X=1.905 $Y=0.74 $X2=0
+ $Y2=0
cc_114 N_A_63_368#_c_106_n N_VGND_c_222_n 0.00132933f $X=1.075 $Y=0.82 $X2=0
+ $Y2=0
cc_115 N_A_63_368#_c_107_n N_VGND_c_222_n 0.0128182f $X=1.615 $Y=1.095 $X2=0
+ $Y2=0
cc_116 N_A_63_368#_c_109_n N_VGND_c_222_n 0.0142456f $X=1.7 $Y=1.63 $X2=0 $Y2=0
cc_117 N_A_63_368#_c_106_n N_VGND_c_225_n 0.00729875f $X=1.075 $Y=0.82 $X2=0
+ $Y2=0
cc_118 N_A_63_368#_M1001_g N_VGND_c_226_n 0.00434272f $X=1.905 $Y=0.74 $X2=0
+ $Y2=0
cc_119 N_A_63_368#_M1001_g N_VGND_c_227_n 0.00828717f $X=1.905 $Y=0.74 $X2=0
+ $Y2=0
cc_120 N_A_63_368#_c_106_n N_VGND_c_227_n 0.00950289f $X=1.075 $Y=0.82 $X2=0
+ $Y2=0
cc_121 N_VPWR_c_173_n X 0.0270509f $X=1.67 $Y=2.455 $X2=0 $Y2=0
cc_122 N_VPWR_c_175_n X 0.0157093f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_123 N_VPWR_c_172_n X 0.0129699f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_124 N_X_c_196_n N_VGND_c_222_n 0.0193831f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_125 N_X_c_196_n N_VGND_c_226_n 0.0156794f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_126 N_X_c_196_n N_VGND_c_227_n 0.0129217f $X=2.12 $Y=0.515 $X2=0 $Y2=0
