* NGSPICE file created from sky130_fd_sc_ls__or4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
M1000 a_446_378# a_216_424# a_357_378# VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=2.95e+11p ps=2.59e+06u
M1001 a_357_378# a_216_424# VGND VNB nshort w=550000u l=150000u
+  ad=3.7675e+11p pd=3.57e+06u as=9.22e+11p ps=7.96e+06u
M1002 a_626_378# B a_530_378# VPB phighvt w=1e+06u l=150000u
+  ad=3.9e+11p pd=2.78e+06u as=3.3e+11p ps=2.66e+06u
M1003 VGND C_N a_27_424# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1004 a_216_424# D_N VGND VNB nshort w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1005 VGND A a_357_378# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_216_424# D_N VPWR VPB phighvt w=840000u l=150000u
+  ad=4.3785e+11p pd=2.97e+06u as=7.664e+11p ps=5.49e+06u
M1007 X a_357_378# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1008 VPWR C_N a_27_424# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1009 a_357_378# B VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_357_378# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1011 a_530_378# a_27_424# a_446_378# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A a_626_378# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_27_424# a_357_378# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

