* File: sky130_fd_sc_ls__a2111o_4.spice
* Created: Wed Sep  2 10:46:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a2111o_4.pex.spice"
.subckt sky130_fd_sc_ls__a2111o_4  VNB VPB D1 C1 B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_137_260#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.8 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_137_260#_M1012_g N_X_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1012_d N_A_137_260#_M1018_g N_X_M1018_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1021_d N_A_137_260#_M1021_g N_X_M1018_s VNB NSHORT L=0.15 W=0.74
+ AD=0.124942 AS=0.1036 PD=1.14217 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1013 N_A_137_260#_M1013_d N_D1_M1013_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.108058 PD=0.92 PS=0.987826 NRD=0 NRS=8.436 M=1 R=4.26667
+ SA=75002 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1019 N_A_137_260#_M1013_d N_D1_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0928 PD=0.92 PS=0.93 NRD=0 NRS=0.936 M=1 R=4.26667 SA=75002.4
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1019_s N_C1_M1003_g N_A_137_260#_M1003_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0928 AS=0.0896 PD=0.93 PS=0.92 NRD=0.936 NRS=0 M=1 R=4.26667 SA=75002.8
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1020 N_VGND_M1020_d N_C1_M1020_g N_A_137_260#_M1003_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0928 AS=0.0896 PD=0.93 PS=0.92 NRD=0.936 NRS=0 M=1 R=4.26667 SA=75003.3
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1020_d N_B1_M1008_g N_A_137_260#_M1008_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0928 AS=0.0896 PD=0.93 PS=0.92 NRD=0.936 NRS=0 M=1 R=4.26667 SA=75003.7
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1024 N_VGND_M1024_d N_B1_M1024_g N_A_137_260#_M1008_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75004.1
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1015 N_A_1210_74#_M1015_d N_A1_M1015_g N_A_137_260#_M1015_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1027 N_A_1210_74#_M1027_d N_A1_M1027_g N_A_137_260#_M1015_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1006 N_A_1210_74#_M1027_d N_A2_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1025 N_A_1210_74#_M1025_d N_A2_M1025_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_X_M1005_d N_A_137_260#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1011 N_X_M1005_d N_A_137_260#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1016 N_X_M1016_d N_A_137_260#_M1016_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1022 N_X_M1016_d N_A_137_260#_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_A_137_260#_M1000_d N_D1_M1000_g N_A_549_392#_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1023 N_A_137_260#_M1000_d N_D1_M1023_g N_A_549_392#_M1023_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.6 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1002 N_A_814_392#_M1002_d N_C1_M1002_g N_A_549_392#_M1023_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1009 N_A_814_392#_M1002_d N_C1_M1009_g N_A_549_392#_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.5 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1007 N_A_814_392#_M1007_d N_B1_M1007_g N_A_1013_392#_M1007_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1014 N_A_814_392#_M1007_d N_B1_M1014_g N_A_1013_392#_M1014_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.6 SB=75002 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1017_d N_A1_M1017_g N_A_1013_392#_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1026 N_VPWR_M1017_d N_A1_M1026_g N_A_1013_392#_M1026_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.5
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A2_M1004_g N_A_1013_392#_M1026_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75002
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1004_d N_A2_M1010_g N_A_1013_392#_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75002.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.8844 P=20.8
c_84 VNB 0 1.80394e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__a2111o_4.pxi.spice"
*
.ends
*
*
