* File: sky130_fd_sc_ls__clkbuf_8.pxi.spice
* Created: Wed Sep  2 10:57:50 2020
* 
x_PM_SKY130_FD_SC_LS__CLKBUF_8%A N_A_c_116_n N_A_M1011_g N_A_M1008_g N_A_M1009_g
+ N_A_c_117_n N_A_M1014_g A A N_A_c_114_n N_A_c_115_n
+ PM_SKY130_FD_SC_LS__CLKBUF_8%A
x_PM_SKY130_FD_SC_LS__CLKBUF_8%A_125_368# N_A_125_368#_M1008_d
+ N_A_125_368#_M1011_s N_A_125_368#_M1000_g N_A_125_368#_c_165_n
+ N_A_125_368#_c_188_n N_A_125_368#_M1001_g N_A_125_368#_c_166_n
+ N_A_125_368#_M1003_g N_A_125_368#_c_190_n N_A_125_368#_M1002_g
+ N_A_125_368#_c_168_n N_A_125_368#_c_192_n N_A_125_368#_M1005_g
+ N_A_125_368#_M1004_g N_A_125_368#_c_170_n N_A_125_368#_c_194_n
+ N_A_125_368#_M1010_g N_A_125_368#_M1006_g N_A_125_368#_c_172_n
+ N_A_125_368#_c_196_n N_A_125_368#_M1012_g N_A_125_368#_M1007_g
+ N_A_125_368#_c_174_n N_A_125_368#_c_198_n N_A_125_368#_M1015_g
+ N_A_125_368#_M1013_g N_A_125_368#_c_176_n N_A_125_368#_c_200_n
+ N_A_125_368#_M1017_g N_A_125_368#_M1016_g N_A_125_368#_c_178_n
+ N_A_125_368#_c_202_n N_A_125_368#_M1019_g N_A_125_368#_M1018_g
+ N_A_125_368#_c_180_n N_A_125_368#_c_209_n N_A_125_368#_c_203_n
+ N_A_125_368#_c_181_n N_A_125_368#_c_182_n N_A_125_368#_c_222_n
+ N_A_125_368#_c_183_n N_A_125_368#_c_184_n N_A_125_368#_c_185_n
+ N_A_125_368#_c_186_n PM_SKY130_FD_SC_LS__CLKBUF_8%A_125_368#
x_PM_SKY130_FD_SC_LS__CLKBUF_8%VPWR N_VPWR_M1011_d N_VPWR_M1014_d N_VPWR_M1002_d
+ N_VPWR_M1010_d N_VPWR_M1015_d N_VPWR_M1019_d N_VPWR_c_382_n N_VPWR_c_383_n
+ N_VPWR_c_384_n N_VPWR_c_385_n N_VPWR_c_386_n N_VPWR_c_387_n N_VPWR_c_388_n
+ N_VPWR_c_389_n N_VPWR_c_390_n VPWR N_VPWR_c_391_n N_VPWR_c_392_n
+ N_VPWR_c_393_n N_VPWR_c_394_n N_VPWR_c_395_n N_VPWR_c_396_n N_VPWR_c_397_n
+ N_VPWR_c_398_n N_VPWR_c_381_n PM_SKY130_FD_SC_LS__CLKBUF_8%VPWR
x_PM_SKY130_FD_SC_LS__CLKBUF_8%X N_X_M1000_s N_X_M1004_s N_X_M1007_s N_X_M1016_s
+ N_X_M1001_s N_X_M1005_s N_X_M1012_s N_X_M1017_s N_X_c_466_n N_X_c_480_n
+ N_X_c_481_n N_X_c_482_n N_X_c_467_n N_X_c_468_n N_X_c_483_n N_X_c_469_n
+ N_X_c_484_n N_X_c_470_n N_X_c_485_n N_X_c_471_n N_X_c_486_n N_X_c_472_n
+ N_X_c_487_n N_X_c_473_n N_X_c_488_n N_X_c_474_n N_X_c_489_n N_X_c_475_n
+ N_X_c_476_n X X X N_X_c_479_n PM_SKY130_FD_SC_LS__CLKBUF_8%X
x_PM_SKY130_FD_SC_LS__CLKBUF_8%VGND N_VGND_M1008_s N_VGND_M1009_s N_VGND_M1003_d
+ N_VGND_M1006_d N_VGND_M1013_d N_VGND_M1018_d N_VGND_c_620_n N_VGND_c_621_n
+ N_VGND_c_622_n N_VGND_c_623_n N_VGND_c_624_n N_VGND_c_625_n N_VGND_c_626_n
+ N_VGND_c_627_n N_VGND_c_628_n N_VGND_c_629_n VGND N_VGND_c_630_n
+ N_VGND_c_631_n N_VGND_c_632_n N_VGND_c_633_n N_VGND_c_634_n N_VGND_c_635_n
+ N_VGND_c_636_n N_VGND_c_637_n PM_SKY130_FD_SC_LS__CLKBUF_8%VGND
cc_1 VNB N_A_M1008_g 0.0550721f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.58
cc_2 VNB N_A_M1009_g 0.0412328f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.58
cc_3 VNB N_A_c_114_n 0.0207044f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.515
cc_4 VNB N_A_c_115_n 0.0421198f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.557
cc_5 VNB N_A_125_368#_M1000_g 0.0345089f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.58
cc_6 VNB N_A_125_368#_c_165_n 0.00807233f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.765
cc_7 VNB N_A_125_368#_c_166_n 0.00738979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_125_368#_M1003_g 0.0332967f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.557
cc_9 VNB N_A_125_368#_c_168_n 0.00739582f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_10 VNB N_A_125_368#_M1004_g 0.0327708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_125_368#_c_170_n 0.00739582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_125_368#_M1006_g 0.029788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_125_368#_c_172_n 0.00739582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_125_368#_M1007_g 0.0297851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_125_368#_c_174_n 0.00767771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_125_368#_M1013_g 0.0312147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_125_368#_c_176_n 0.00774612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_125_368#_M1016_g 0.0311717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_125_368#_c_178_n 0.00909136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_125_368#_M1018_g 0.0380131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_125_368#_c_180_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_125_368#_c_181_n 0.00948747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_125_368#_c_182_n 0.00244471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_125_368#_c_183_n 0.00215284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_125_368#_c_184_n 0.00141621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_125_368#_c_185_n 0.00727321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_125_368#_c_186_n 0.17485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_381_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_466_n 0.00356116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_467_n 0.00791479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_468_n 0.00319211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_469_n 0.00261846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_470_n 0.0075697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_471_n 0.00284218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_472_n 0.00860164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_473_n 0.00325795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_474_n 0.00177795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_475_n 0.00125222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_476_n 0.0111242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB X 0.0135769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB X 0.0110186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_X_c_479_n 0.00551646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_620_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.557
cc_44 VNB N_VGND_c_621_n 0.0348648f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.557
cc_45 VNB N_VGND_c_622_n 0.0118552f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.557
cc_46 VNB N_VGND_c_623_n 0.018682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_624_n 0.00817312f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.565
cc_48 VNB N_VGND_c_625_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_626_n 0.002601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_627_n 0.00250542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_628_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_629_n 0.021573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_630_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_631_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_632_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_633_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_634_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_635_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_636_n 0.00732404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_637_n 0.286414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VPB N_A_c_116_n 0.0180026f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=1.765
cc_62 VPB N_A_c_117_n 0.0164958f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_63 VPB N_A_c_114_n 0.0133503f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.515
cc_64 VPB N_A_c_115_n 0.0222109f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.557
cc_65 VPB N_A_125_368#_c_165_n 8.1304e-19 $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_66 VPB N_A_125_368#_c_188_n 0.0224062f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_67 VPB N_A_125_368#_c_166_n 7.44295e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_125_368#_c_190_n 0.0194687f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.515
cc_69 VPB N_A_125_368#_c_168_n 7.44903e-19 $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_70 VPB N_A_125_368#_c_192_n 0.0194706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_125_368#_c_170_n 7.44903e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_125_368#_c_194_n 0.0199761f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_125_368#_c_172_n 7.44903e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_125_368#_c_196_n 0.0199759f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_125_368#_c_174_n 7.73294e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_125_368#_c_198_n 0.020027f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_125_368#_c_176_n 7.80184e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_125_368#_c_200_n 0.0206087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_125_368#_c_178_n 9.15677e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_125_368#_c_202_n 0.023905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_125_368#_c_203_n 0.00261637f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_125_368#_c_183_n 0.00329058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_382_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=1.557
cc_84 VPB N_VPWR_c_383_n 0.0513909f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.557
cc_85 VPB N_VPWR_c_384_n 0.00820985f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_385_n 0.0027821f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.565
cc_87 VPB N_VPWR_c_386_n 0.0184472f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_387_n 0.00670059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_388_n 0.00524329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_389_n 0.0121701f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_390_n 0.0449489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_391_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_392_n 0.0174535f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_393_n 0.0184081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_394_n 0.0179698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_395_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_396_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_397_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_398_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_381_n 0.0745543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_X_c_480_n 0.00230039f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.565
cc_102 VPB N_X_c_481_n 0.0028649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_X_c_482_n 0.0019142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_X_c_483_n 0.00225498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_X_c_484_n 0.00219429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_X_c_485_n 0.00230039f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_X_c_486_n 0.00280702f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_X_c_487_n 0.00262951f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_X_c_488_n 0.00186725f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_X_c_489_n 0.0019142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB X 0.0136246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 N_A_M1009_g N_A_125_368#_M1000_g 0.0215792f $X=0.995 $Y=0.58 $X2=0 $Y2=0
cc_113 N_A_c_117_n N_A_125_368#_c_188_n 0.0289517f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_114 N_A_M1008_g N_A_125_368#_c_180_n 0.0153383f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_115 N_A_M1009_g N_A_125_368#_c_180_n 0.0112601f $X=0.995 $Y=0.58 $X2=0 $Y2=0
cc_116 N_A_c_116_n N_A_125_368#_c_209_n 0.00177269f $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A_c_117_n N_A_125_368#_c_209_n 4.27055e-19 $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_118 N_A_c_114_n N_A_125_368#_c_209_n 0.0237949f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_119 N_A_c_115_n N_A_125_368#_c_209_n 0.00147208f $X=0.995 $Y=1.557 $X2=0
+ $Y2=0
cc_120 N_A_c_116_n N_A_125_368#_c_203_n 0.00859489f $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A_c_117_n N_A_125_368#_c_203_n 0.0103171f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A_M1009_g N_A_125_368#_c_181_n 0.0116275f $X=0.995 $Y=0.58 $X2=0 $Y2=0
cc_123 N_A_c_114_n N_A_125_368#_c_181_n 0.00967513f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_124 N_A_c_115_n N_A_125_368#_c_181_n 6.03517e-19 $X=0.995 $Y=1.557 $X2=0
+ $Y2=0
cc_125 N_A_M1008_g N_A_125_368#_c_182_n 0.010444f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_126 N_A_M1009_g N_A_125_368#_c_182_n 0.0028254f $X=0.995 $Y=0.58 $X2=0 $Y2=0
cc_127 N_A_c_114_n N_A_125_368#_c_182_n 0.024859f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A_c_115_n N_A_125_368#_c_182_n 0.00229418f $X=0.995 $Y=1.557 $X2=0
+ $Y2=0
cc_129 N_A_c_117_n N_A_125_368#_c_222_n 0.012208f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A_c_114_n N_A_125_368#_c_222_n 0.0104662f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_131 N_A_c_117_n N_A_125_368#_c_183_n 0.0036594f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_132 N_A_c_114_n N_A_125_368#_c_183_n 0.0198451f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A_c_115_n N_A_125_368#_c_183_n 8.37278e-19 $X=0.995 $Y=1.557 $X2=0
+ $Y2=0
cc_134 N_A_M1009_g N_A_125_368#_c_185_n 0.00523978f $X=0.995 $Y=0.58 $X2=0 $Y2=0
cc_135 N_A_c_114_n N_A_125_368#_c_185_n 0.0144263f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A_c_115_n N_A_125_368#_c_185_n 7.26037e-19 $X=0.995 $Y=1.557 $X2=0
+ $Y2=0
cc_137 N_A_c_114_n N_A_125_368#_c_186_n 2.4102e-19 $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A_c_115_n N_A_125_368#_c_186_n 0.0120816f $X=0.995 $Y=1.557 $X2=0 $Y2=0
cc_139 N_A_c_116_n N_VPWR_c_383_n 0.00378733f $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A_c_114_n N_VPWR_c_383_n 0.0270496f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A_c_117_n N_VPWR_c_384_n 0.00598632f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A_c_116_n N_VPWR_c_391_n 0.00451267f $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A_c_117_n N_VPWR_c_391_n 0.00445602f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A_c_116_n N_VPWR_c_381_n 0.00878831f $X=0.55 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A_c_117_n N_VPWR_c_381_n 0.00857873f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A_c_117_n N_X_c_480_n 7.99369e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A_M1009_g N_X_c_468_n 4.16027e-19 $X=0.995 $Y=0.58 $X2=0 $Y2=0
cc_148 N_A_M1008_g N_VGND_c_621_n 0.0122932f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_149 N_A_c_114_n N_VGND_c_621_n 0.0127936f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_150 N_A_c_115_n N_VGND_c_621_n 3.45262e-19 $X=0.995 $Y=1.557 $X2=0 $Y2=0
cc_151 N_A_M1009_g N_VGND_c_622_n 0.00455328f $X=0.995 $Y=0.58 $X2=0 $Y2=0
cc_152 N_A_M1008_g N_VGND_c_630_n 0.00434272f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_153 N_A_M1009_g N_VGND_c_630_n 0.00434272f $X=0.995 $Y=0.58 $X2=0 $Y2=0
cc_154 N_A_M1008_g N_VGND_c_637_n 0.00823934f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_155 N_A_M1009_g N_VGND_c_637_n 0.00821127f $X=0.995 $Y=0.58 $X2=0 $Y2=0
cc_156 N_A_125_368#_c_222_n N_VPWR_M1014_d 0.00983318f $X=1.275 $Y=2.035 $X2=0
+ $Y2=0
cc_157 N_A_125_368#_c_183_n N_VPWR_M1014_d 0.00217326f $X=1.36 $Y=1.95 $X2=0
+ $Y2=0
cc_158 N_A_125_368#_c_203_n N_VPWR_c_383_n 0.0330222f $X=0.78 $Y=2.815 $X2=0
+ $Y2=0
cc_159 N_A_125_368#_c_188_n N_VPWR_c_384_n 0.00592199f $X=1.555 $Y=1.765 $X2=0
+ $Y2=0
cc_160 N_A_125_368#_c_203_n N_VPWR_c_384_n 0.0266809f $X=0.78 $Y=2.815 $X2=0
+ $Y2=0
cc_161 N_A_125_368#_c_222_n N_VPWR_c_384_n 0.0244899f $X=1.275 $Y=2.035 $X2=0
+ $Y2=0
cc_162 N_A_125_368#_c_188_n N_VPWR_c_385_n 6.32513e-19 $X=1.555 $Y=1.765 $X2=0
+ $Y2=0
cc_163 N_A_125_368#_c_190_n N_VPWR_c_385_n 0.0134177f $X=2.005 $Y=1.765 $X2=0
+ $Y2=0
cc_164 N_A_125_368#_c_192_n N_VPWR_c_385_n 0.0135755f $X=2.455 $Y=1.765 $X2=0
+ $Y2=0
cc_165 N_A_125_368#_c_194_n N_VPWR_c_385_n 6.43035e-19 $X=2.905 $Y=1.765 $X2=0
+ $Y2=0
cc_166 N_A_125_368#_c_192_n N_VPWR_c_386_n 0.00413917f $X=2.455 $Y=1.765 $X2=0
+ $Y2=0
cc_167 N_A_125_368#_c_194_n N_VPWR_c_386_n 0.00445602f $X=2.905 $Y=1.765 $X2=0
+ $Y2=0
cc_168 N_A_125_368#_c_194_n N_VPWR_c_387_n 0.00549464f $X=2.905 $Y=1.765 $X2=0
+ $Y2=0
cc_169 N_A_125_368#_c_196_n N_VPWR_c_387_n 0.00549464f $X=3.355 $Y=1.765 $X2=0
+ $Y2=0
cc_170 N_A_125_368#_c_196_n N_VPWR_c_388_n 6.36276e-19 $X=3.355 $Y=1.765 $X2=0
+ $Y2=0
cc_171 N_A_125_368#_c_198_n N_VPWR_c_388_n 0.0134008f $X=3.805 $Y=1.765 $X2=0
+ $Y2=0
cc_172 N_A_125_368#_c_200_n N_VPWR_c_388_n 0.00682709f $X=4.305 $Y=1.765 $X2=0
+ $Y2=0
cc_173 N_A_125_368#_c_200_n N_VPWR_c_390_n 5.93605e-19 $X=4.305 $Y=1.765 $X2=0
+ $Y2=0
cc_174 N_A_125_368#_c_202_n N_VPWR_c_390_n 0.0144671f $X=4.77 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_A_125_368#_c_203_n N_VPWR_c_391_n 0.0145669f $X=0.78 $Y=2.815 $X2=0
+ $Y2=0
cc_176 N_A_125_368#_c_188_n N_VPWR_c_392_n 0.00445602f $X=1.555 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_A_125_368#_c_190_n N_VPWR_c_392_n 0.00413917f $X=2.005 $Y=1.765 $X2=0
+ $Y2=0
cc_178 N_A_125_368#_c_196_n N_VPWR_c_393_n 0.00445602f $X=3.355 $Y=1.765 $X2=0
+ $Y2=0
cc_179 N_A_125_368#_c_198_n N_VPWR_c_393_n 0.00413917f $X=3.805 $Y=1.765 $X2=0
+ $Y2=0
cc_180 N_A_125_368#_c_200_n N_VPWR_c_394_n 0.00461464f $X=4.305 $Y=1.765 $X2=0
+ $Y2=0
cc_181 N_A_125_368#_c_202_n N_VPWR_c_394_n 0.00413917f $X=4.77 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A_125_368#_c_188_n N_VPWR_c_381_n 0.00857825f $X=1.555 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A_125_368#_c_190_n N_VPWR_c_381_n 0.00817726f $X=2.005 $Y=1.765 $X2=0
+ $Y2=0
cc_184 N_A_125_368#_c_192_n N_VPWR_c_381_n 0.00817726f $X=2.455 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A_125_368#_c_194_n N_VPWR_c_381_n 0.00857589f $X=2.905 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_A_125_368#_c_196_n N_VPWR_c_381_n 0.00857589f $X=3.355 $Y=1.765 $X2=0
+ $Y2=0
cc_187 N_A_125_368#_c_198_n N_VPWR_c_381_n 0.00817726f $X=3.805 $Y=1.765 $X2=0
+ $Y2=0
cc_188 N_A_125_368#_c_200_n N_VPWR_c_381_n 0.00908883f $X=4.305 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_A_125_368#_c_202_n N_VPWR_c_381_n 0.00817869f $X=4.77 $Y=1.765 $X2=0
+ $Y2=0
cc_190 N_A_125_368#_c_203_n N_VPWR_c_381_n 0.0120032f $X=0.78 $Y=2.815 $X2=0
+ $Y2=0
cc_191 N_A_125_368#_M1000_g N_X_c_466_n 0.00114369f $X=1.54 $Y=0.58 $X2=0 $Y2=0
cc_192 N_A_125_368#_M1003_g N_X_c_466_n 0.00829498f $X=1.995 $Y=0.58 $X2=0 $Y2=0
cc_193 N_A_125_368#_M1004_g N_X_c_466_n 5.97046e-19 $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_194 N_A_125_368#_c_180_n N_X_c_466_n 0.00108577f $X=0.78 $Y=0.58 $X2=0 $Y2=0
cc_195 N_A_125_368#_c_188_n N_X_c_480_n 0.0132531f $X=1.555 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A_125_368#_c_190_n N_X_c_480_n 3.80067e-19 $X=2.005 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_A_125_368#_c_203_n N_X_c_480_n 0.00397297f $X=0.78 $Y=2.815 $X2=0 $Y2=0
cc_198 N_A_125_368#_c_190_n N_X_c_481_n 0.015489f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A_125_368#_c_192_n N_X_c_481_n 0.015489f $X=2.455 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A_125_368#_c_184_n N_X_c_481_n 0.0515664f $X=4.35 $Y=1.355 $X2=0 $Y2=0
cc_201 N_A_125_368#_c_186_n N_X_c_481_n 0.00201785f $X=4.785 $Y=1.355 $X2=0
+ $Y2=0
cc_202 N_A_125_368#_c_188_n N_X_c_482_n 0.00437905f $X=1.555 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_A_125_368#_c_183_n N_X_c_482_n 0.0127483f $X=1.36 $Y=1.95 $X2=0 $Y2=0
cc_204 N_A_125_368#_c_184_n N_X_c_482_n 0.022216f $X=4.35 $Y=1.355 $X2=0 $Y2=0
cc_205 N_A_125_368#_c_186_n N_X_c_482_n 0.00209661f $X=4.785 $Y=1.355 $X2=0
+ $Y2=0
cc_206 N_A_125_368#_M1003_g N_X_c_467_n 0.00927712f $X=1.995 $Y=0.58 $X2=0 $Y2=0
cc_207 N_A_125_368#_M1004_g N_X_c_467_n 0.00927712f $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_208 N_A_125_368#_c_184_n N_X_c_467_n 0.0493541f $X=4.35 $Y=1.355 $X2=0 $Y2=0
cc_209 N_A_125_368#_c_186_n N_X_c_467_n 0.00595379f $X=4.785 $Y=1.355 $X2=0
+ $Y2=0
cc_210 N_A_125_368#_M1000_g N_X_c_468_n 0.002818f $X=1.54 $Y=0.58 $X2=0 $Y2=0
cc_211 N_A_125_368#_M1003_g N_X_c_468_n 0.00287638f $X=1.995 $Y=0.58 $X2=0 $Y2=0
cc_212 N_A_125_368#_c_180_n N_X_c_468_n 0.00327297f $X=0.78 $Y=0.58 $X2=0 $Y2=0
cc_213 N_A_125_368#_c_184_n N_X_c_468_n 0.027687f $X=4.35 $Y=1.355 $X2=0 $Y2=0
cc_214 N_A_125_368#_c_185_n N_X_c_468_n 0.00356562f $X=1.36 $Y=1.25 $X2=0 $Y2=0
cc_215 N_A_125_368#_c_186_n N_X_c_468_n 0.0030438f $X=4.785 $Y=1.355 $X2=0 $Y2=0
cc_216 N_A_125_368#_c_192_n N_X_c_483_n 3.77415e-19 $X=2.455 $Y=1.765 $X2=0
+ $Y2=0
cc_217 N_A_125_368#_c_194_n N_X_c_483_n 0.0134289f $X=2.905 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A_125_368#_c_196_n N_X_c_483_n 7.27152e-19 $X=3.355 $Y=1.765 $X2=0
+ $Y2=0
cc_219 N_A_125_368#_M1003_g N_X_c_469_n 5.98311e-19 $X=1.995 $Y=0.58 $X2=0 $Y2=0
cc_220 N_A_125_368#_M1004_g N_X_c_469_n 0.00807849f $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_221 N_A_125_368#_M1006_g N_X_c_469_n 0.00176975f $X=2.995 $Y=0.58 $X2=0 $Y2=0
cc_222 N_A_125_368#_c_194_n N_X_c_484_n 0.0124531f $X=2.905 $Y=1.765 $X2=0 $Y2=0
cc_223 N_A_125_368#_c_196_n N_X_c_484_n 0.0124531f $X=3.355 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A_125_368#_c_184_n N_X_c_484_n 0.0416512f $X=4.35 $Y=1.355 $X2=0 $Y2=0
cc_225 N_A_125_368#_c_186_n N_X_c_484_n 0.00231334f $X=4.785 $Y=1.355 $X2=0
+ $Y2=0
cc_226 N_A_125_368#_M1006_g N_X_c_470_n 0.0117051f $X=2.995 $Y=0.58 $X2=0 $Y2=0
cc_227 N_A_125_368#_M1007_g N_X_c_470_n 0.0117051f $X=3.425 $Y=0.58 $X2=0 $Y2=0
cc_228 N_A_125_368#_c_184_n N_X_c_470_n 0.0506643f $X=4.35 $Y=1.355 $X2=0 $Y2=0
cc_229 N_A_125_368#_c_186_n N_X_c_470_n 0.00257695f $X=4.785 $Y=1.355 $X2=0
+ $Y2=0
cc_230 N_A_125_368#_c_194_n N_X_c_485_n 7.2695e-19 $X=2.905 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A_125_368#_c_196_n N_X_c_485_n 0.0134353f $X=3.355 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A_125_368#_c_198_n N_X_c_485_n 3.80067e-19 $X=3.805 $Y=1.765 $X2=0
+ $Y2=0
cc_233 N_A_125_368#_M1007_g N_X_c_471_n 0.00165866f $X=3.425 $Y=0.58 $X2=0 $Y2=0
cc_234 N_A_125_368#_M1013_g N_X_c_471_n 0.00165866f $X=3.855 $Y=0.58 $X2=0 $Y2=0
cc_235 N_A_125_368#_c_198_n N_X_c_486_n 0.0157707f $X=3.805 $Y=1.765 $X2=0 $Y2=0
cc_236 N_A_125_368#_c_200_n N_X_c_486_n 0.0149111f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A_125_368#_c_184_n N_X_c_486_n 0.0613413f $X=4.35 $Y=1.355 $X2=0 $Y2=0
cc_238 N_A_125_368#_c_186_n N_X_c_486_n 0.00327677f $X=4.785 $Y=1.355 $X2=0
+ $Y2=0
cc_239 N_A_125_368#_M1013_g N_X_c_472_n 0.0120984f $X=3.855 $Y=0.58 $X2=0 $Y2=0
cc_240 N_A_125_368#_M1016_g N_X_c_472_n 0.0120518f $X=4.355 $Y=0.58 $X2=0 $Y2=0
cc_241 N_A_125_368#_c_184_n N_X_c_472_n 0.0581804f $X=4.35 $Y=1.355 $X2=0 $Y2=0
cc_242 N_A_125_368#_c_186_n N_X_c_472_n 0.00406759f $X=4.785 $Y=1.355 $X2=0
+ $Y2=0
cc_243 N_A_125_368#_c_200_n N_X_c_487_n 4.34097e-19 $X=4.305 $Y=1.765 $X2=0
+ $Y2=0
cc_244 N_A_125_368#_c_202_n N_X_c_487_n 3.93489e-19 $X=4.77 $Y=1.765 $X2=0 $Y2=0
cc_245 N_A_125_368#_M1016_g N_X_c_473_n 0.00167832f $X=4.355 $Y=0.58 $X2=0 $Y2=0
cc_246 N_A_125_368#_M1018_g N_X_c_473_n 0.00167832f $X=4.785 $Y=0.58 $X2=0 $Y2=0
cc_247 N_A_125_368#_c_194_n N_X_c_488_n 0.00294438f $X=2.905 $Y=1.765 $X2=0
+ $Y2=0
cc_248 N_A_125_368#_c_184_n N_X_c_488_n 0.0217942f $X=4.35 $Y=1.355 $X2=0 $Y2=0
cc_249 N_A_125_368#_c_186_n N_X_c_488_n 0.00245159f $X=4.785 $Y=1.355 $X2=0
+ $Y2=0
cc_250 N_A_125_368#_M1004_g N_X_c_474_n 0.00277836f $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_251 N_A_125_368#_c_184_n N_X_c_474_n 0.0209476f $X=4.35 $Y=1.355 $X2=0 $Y2=0
cc_252 N_A_125_368#_c_186_n N_X_c_474_n 0.00270087f $X=4.785 $Y=1.355 $X2=0
+ $Y2=0
cc_253 N_A_125_368#_c_196_n N_X_c_489_n 0.00294667f $X=3.355 $Y=1.765 $X2=0
+ $Y2=0
cc_254 N_A_125_368#_c_184_n N_X_c_489_n 0.022216f $X=4.35 $Y=1.355 $X2=0 $Y2=0
cc_255 N_A_125_368#_c_186_n N_X_c_489_n 0.00231354f $X=4.785 $Y=1.355 $X2=0
+ $Y2=0
cc_256 N_A_125_368#_c_184_n N_X_c_475_n 0.0143206f $X=4.35 $Y=1.355 $X2=0 $Y2=0
cc_257 N_A_125_368#_c_186_n N_X_c_475_n 0.00258098f $X=4.785 $Y=1.355 $X2=0
+ $Y2=0
cc_258 N_A_125_368#_M1018_g N_X_c_476_n 0.0105097f $X=4.785 $Y=0.58 $X2=0 $Y2=0
cc_259 N_A_125_368#_c_186_n N_X_c_476_n 0.00285269f $X=4.785 $Y=1.355 $X2=0
+ $Y2=0
cc_260 N_A_125_368#_M1018_g X 4.35224e-19 $X=4.785 $Y=0.58 $X2=0 $Y2=0
cc_261 N_A_125_368#_c_184_n X 0.0239264f $X=4.35 $Y=1.355 $X2=0 $Y2=0
cc_262 N_A_125_368#_c_186_n X 0.0104476f $X=4.785 $Y=1.355 $X2=0 $Y2=0
cc_263 N_A_125_368#_c_176_n X 9.98591e-19 $X=4.305 $Y=1.675 $X2=0 $Y2=0
cc_264 N_A_125_368#_c_200_n X 0.00124882f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_265 N_A_125_368#_c_178_n X 0.00749165f $X=4.77 $Y=1.675 $X2=0 $Y2=0
cc_266 N_A_125_368#_c_202_n X 0.0169947f $X=4.77 $Y=1.765 $X2=0 $Y2=0
cc_267 N_A_125_368#_c_186_n X 0.00862043f $X=4.785 $Y=1.355 $X2=0 $Y2=0
cc_268 N_A_125_368#_M1016_g N_X_c_479_n 0.00106492f $X=4.355 $Y=0.58 $X2=0 $Y2=0
cc_269 N_A_125_368#_M1018_g N_X_c_479_n 0.00699065f $X=4.785 $Y=0.58 $X2=0 $Y2=0
cc_270 N_A_125_368#_c_180_n N_VGND_c_621_n 0.0188413f $X=0.78 $Y=0.58 $X2=0
+ $Y2=0
cc_271 N_A_125_368#_M1000_g N_VGND_c_622_n 0.00242063f $X=1.54 $Y=0.58 $X2=0
+ $Y2=0
cc_272 N_A_125_368#_c_180_n N_VGND_c_622_n 0.0188413f $X=0.78 $Y=0.58 $X2=0
+ $Y2=0
cc_273 N_A_125_368#_c_181_n N_VGND_c_622_n 0.0133914f $X=1.275 $Y=1.065 $X2=0
+ $Y2=0
cc_274 N_A_125_368#_c_185_n N_VGND_c_622_n 0.0158349f $X=1.36 $Y=1.25 $X2=0
+ $Y2=0
cc_275 N_A_125_368#_M1000_g N_VGND_c_623_n 0.00461464f $X=1.54 $Y=0.58 $X2=0
+ $Y2=0
cc_276 N_A_125_368#_M1003_g N_VGND_c_623_n 0.00434272f $X=1.995 $Y=0.58 $X2=0
+ $Y2=0
cc_277 N_A_125_368#_M1003_g N_VGND_c_624_n 0.00387235f $X=1.995 $Y=0.58 $X2=0
+ $Y2=0
cc_278 N_A_125_368#_M1004_g N_VGND_c_624_n 0.0037829f $X=2.565 $Y=0.58 $X2=0
+ $Y2=0
cc_279 N_A_125_368#_M1004_g N_VGND_c_625_n 0.00434272f $X=2.565 $Y=0.58 $X2=0
+ $Y2=0
cc_280 N_A_125_368#_M1006_g N_VGND_c_625_n 0.00383152f $X=2.995 $Y=0.58 $X2=0
+ $Y2=0
cc_281 N_A_125_368#_M1004_g N_VGND_c_626_n 4.49641e-19 $X=2.565 $Y=0.58 $X2=0
+ $Y2=0
cc_282 N_A_125_368#_M1006_g N_VGND_c_626_n 0.00780668f $X=2.995 $Y=0.58 $X2=0
+ $Y2=0
cc_283 N_A_125_368#_M1007_g N_VGND_c_626_n 0.00768587f $X=3.425 $Y=0.58 $X2=0
+ $Y2=0
cc_284 N_A_125_368#_M1013_g N_VGND_c_626_n 4.2389e-19 $X=3.855 $Y=0.58 $X2=0
+ $Y2=0
cc_285 N_A_125_368#_M1007_g N_VGND_c_627_n 4.23177e-19 $X=3.425 $Y=0.58 $X2=0
+ $Y2=0
cc_286 N_A_125_368#_M1013_g N_VGND_c_627_n 0.00798783f $X=3.855 $Y=0.58 $X2=0
+ $Y2=0
cc_287 N_A_125_368#_M1016_g N_VGND_c_627_n 0.00798783f $X=4.355 $Y=0.58 $X2=0
+ $Y2=0
cc_288 N_A_125_368#_M1018_g N_VGND_c_627_n 4.23177e-19 $X=4.785 $Y=0.58 $X2=0
+ $Y2=0
cc_289 N_A_125_368#_M1016_g N_VGND_c_629_n 4.2389e-19 $X=4.355 $Y=0.58 $X2=0
+ $Y2=0
cc_290 N_A_125_368#_M1018_g N_VGND_c_629_n 0.00874936f $X=4.785 $Y=0.58 $X2=0
+ $Y2=0
cc_291 N_A_125_368#_c_180_n N_VGND_c_630_n 0.0144922f $X=0.78 $Y=0.58 $X2=0
+ $Y2=0
cc_292 N_A_125_368#_M1007_g N_VGND_c_631_n 0.00383152f $X=3.425 $Y=0.58 $X2=0
+ $Y2=0
cc_293 N_A_125_368#_M1013_g N_VGND_c_631_n 0.00383152f $X=3.855 $Y=0.58 $X2=0
+ $Y2=0
cc_294 N_A_125_368#_M1016_g N_VGND_c_632_n 0.00383152f $X=4.355 $Y=0.58 $X2=0
+ $Y2=0
cc_295 N_A_125_368#_M1018_g N_VGND_c_632_n 0.00383152f $X=4.785 $Y=0.58 $X2=0
+ $Y2=0
cc_296 N_A_125_368#_M1000_g N_VGND_c_637_n 0.00908861f $X=1.54 $Y=0.58 $X2=0
+ $Y2=0
cc_297 N_A_125_368#_M1003_g N_VGND_c_637_n 0.0044839f $X=1.995 $Y=0.58 $X2=0
+ $Y2=0
cc_298 N_A_125_368#_M1004_g N_VGND_c_637_n 0.00448145f $X=2.565 $Y=0.58 $X2=0
+ $Y2=0
cc_299 N_A_125_368#_M1006_g N_VGND_c_637_n 0.00386058f $X=2.995 $Y=0.58 $X2=0
+ $Y2=0
cc_300 N_A_125_368#_M1007_g N_VGND_c_637_n 0.00386058f $X=3.425 $Y=0.58 $X2=0
+ $Y2=0
cc_301 N_A_125_368#_M1013_g N_VGND_c_637_n 0.00386058f $X=3.855 $Y=0.58 $X2=0
+ $Y2=0
cc_302 N_A_125_368#_M1016_g N_VGND_c_637_n 0.00386058f $X=4.355 $Y=0.58 $X2=0
+ $Y2=0
cc_303 N_A_125_368#_M1018_g N_VGND_c_637_n 0.00386058f $X=4.785 $Y=0.58 $X2=0
+ $Y2=0
cc_304 N_A_125_368#_c_180_n N_VGND_c_637_n 0.0118826f $X=0.78 $Y=0.58 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_384_n N_X_c_480_n 0.0258252f $X=1.28 $Y=2.455 $X2=0 $Y2=0
cc_306 N_VPWR_c_385_n N_X_c_480_n 0.0340309f $X=2.23 $Y=2.115 $X2=0 $Y2=0
cc_307 N_VPWR_c_392_n N_X_c_480_n 0.0116935f $X=2.065 $Y=3.33 $X2=0 $Y2=0
cc_308 N_VPWR_c_381_n N_X_c_480_n 0.00964594f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_309 N_VPWR_M1002_d N_X_c_481_n 0.00197722f $X=2.08 $Y=1.84 $X2=0 $Y2=0
cc_310 N_VPWR_c_385_n N_X_c_481_n 0.0171813f $X=2.23 $Y=2.115 $X2=0 $Y2=0
cc_311 N_VPWR_c_385_n N_X_c_483_n 0.0333124f $X=2.23 $Y=2.115 $X2=0 $Y2=0
cc_312 N_VPWR_c_386_n N_X_c_483_n 0.0114703f $X=3.045 $Y=3.33 $X2=0 $Y2=0
cc_313 N_VPWR_c_387_n N_X_c_483_n 0.0607847f $X=3.13 $Y=2.195 $X2=0 $Y2=0
cc_314 N_VPWR_c_381_n N_X_c_483_n 0.00946127f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_315 N_VPWR_M1010_d N_X_c_484_n 0.00247267f $X=2.98 $Y=1.84 $X2=0 $Y2=0
cc_316 N_VPWR_c_387_n N_X_c_484_n 0.0136682f $X=3.13 $Y=2.195 $X2=0 $Y2=0
cc_317 N_VPWR_c_387_n N_X_c_485_n 0.0608729f $X=3.13 $Y=2.195 $X2=0 $Y2=0
cc_318 N_VPWR_c_388_n N_X_c_485_n 0.0340309f $X=4.03 $Y=2.115 $X2=0 $Y2=0
cc_319 N_VPWR_c_393_n N_X_c_485_n 0.0116935f $X=3.865 $Y=3.33 $X2=0 $Y2=0
cc_320 N_VPWR_c_381_n N_X_c_485_n 0.00964594f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_321 N_VPWR_M1015_d N_X_c_486_n 0.00250873f $X=3.88 $Y=1.84 $X2=0 $Y2=0
cc_322 N_VPWR_c_388_n N_X_c_486_n 0.0202249f $X=4.03 $Y=2.115 $X2=0 $Y2=0
cc_323 N_VPWR_c_388_n N_X_c_487_n 0.00143579f $X=4.03 $Y=2.115 $X2=0 $Y2=0
cc_324 N_VPWR_c_390_n N_X_c_487_n 0.0340288f $X=4.995 $Y=2.115 $X2=0 $Y2=0
cc_325 N_VPWR_c_394_n N_X_c_487_n 0.0115122f $X=4.83 $Y=3.33 $X2=0 $Y2=0
cc_326 N_VPWR_c_381_n N_X_c_487_n 0.0095288f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_327 N_VPWR_M1019_d X 0.00263515f $X=4.845 $Y=1.84 $X2=0 $Y2=0
cc_328 N_VPWR_c_390_n X 0.0216168f $X=4.995 $Y=2.115 $X2=0 $Y2=0
cc_329 N_X_c_466_n N_VGND_c_622_n 0.0193875f $X=1.78 $Y=0.58 $X2=0 $Y2=0
cc_330 N_X_c_466_n N_VGND_c_623_n 0.0145482f $X=1.78 $Y=0.58 $X2=0 $Y2=0
cc_331 N_X_c_466_n N_VGND_c_624_n 0.0131729f $X=1.78 $Y=0.58 $X2=0 $Y2=0
cc_332 N_X_c_467_n N_VGND_c_624_n 0.0255516f $X=2.615 $Y=0.935 $X2=0 $Y2=0
cc_333 N_X_c_469_n N_VGND_c_624_n 0.0126571f $X=2.78 $Y=0.58 $X2=0 $Y2=0
cc_334 N_X_c_469_n N_VGND_c_625_n 0.0109824f $X=2.78 $Y=0.58 $X2=0 $Y2=0
cc_335 N_X_c_469_n N_VGND_c_626_n 0.0125556f $X=2.78 $Y=0.58 $X2=0 $Y2=0
cc_336 N_X_c_470_n N_VGND_c_626_n 0.021034f $X=3.555 $Y=0.935 $X2=0 $Y2=0
cc_337 N_X_c_471_n N_VGND_c_626_n 0.0125142f $X=3.64 $Y=0.58 $X2=0 $Y2=0
cc_338 N_X_c_471_n N_VGND_c_627_n 0.0128675f $X=3.64 $Y=0.58 $X2=0 $Y2=0
cc_339 N_X_c_472_n N_VGND_c_627_n 0.0266978f $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_340 N_X_c_473_n N_VGND_c_627_n 0.0128675f $X=4.57 $Y=0.58 $X2=0 $Y2=0
cc_341 N_X_c_473_n N_VGND_c_629_n 0.0125142f $X=4.57 $Y=0.58 $X2=0 $Y2=0
cc_342 N_X_c_476_n N_VGND_c_629_n 0.00246824f $X=4.795 $Y=0.935 $X2=0 $Y2=0
cc_343 X N_VGND_c_629_n 0.0105914f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_344 N_X_c_471_n N_VGND_c_631_n 0.0074882f $X=3.64 $Y=0.58 $X2=0 $Y2=0
cc_345 N_X_c_473_n N_VGND_c_632_n 0.00733159f $X=4.57 $Y=0.58 $X2=0 $Y2=0
cc_346 N_X_c_466_n N_VGND_c_637_n 0.0119922f $X=1.78 $Y=0.58 $X2=0 $Y2=0
cc_347 N_X_c_467_n N_VGND_c_637_n 0.0109408f $X=2.615 $Y=0.935 $X2=0 $Y2=0
cc_348 N_X_c_469_n N_VGND_c_637_n 0.00903908f $X=2.78 $Y=0.58 $X2=0 $Y2=0
cc_349 N_X_c_470_n N_VGND_c_637_n 0.0115904f $X=3.555 $Y=0.935 $X2=0 $Y2=0
cc_350 N_X_c_471_n N_VGND_c_637_n 0.00620166f $X=3.64 $Y=0.58 $X2=0 $Y2=0
cc_351 N_X_c_472_n N_VGND_c_637_n 0.0171812f $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_352 N_X_c_473_n N_VGND_c_637_n 0.00614141f $X=4.57 $Y=0.58 $X2=0 $Y2=0
