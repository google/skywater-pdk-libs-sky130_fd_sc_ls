* NGSPICE file created from sky130_fd_sc_ls__nor4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
M1000 a_498_368# C a_229_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=9.968e+11p ps=8.5e+06u
M1001 Y B VGND VNB nshort w=740000u l=150000u
+  ad=9.879e+11p pd=8.59e+06u as=1.7479e+12p ps=1.217e+07u
M1002 a_229_368# C a_498_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_27_392# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_498_368# B a_701_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=9.968e+11p ps=8.5e+06u
M1006 Y a_27_392# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND C Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y a_27_392# a_229_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1009 VGND B Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_701_368# B a_498_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_701_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.422e+11p ps=5.45e+06u
M1013 VPWR D_N a_27_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1014 a_229_368# a_27_392# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A a_701_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y C VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND D_N a_27_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
.ends

