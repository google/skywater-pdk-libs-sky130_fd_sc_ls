* File: sky130_fd_sc_ls__ha_4.pex.spice
* Created: Fri Aug 28 13:27:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__HA_4%A_435_99# 1 2 3 10 12 13 14 15 17 18 20 21 23
+ 24 26 29 31 33 36 38 40 43 45 47 50 52 55 59 63 66 68 69 74 78 81 94
c192 68 0 1.09796e-19 $X=5.965 $Y=1.82
c193 10 0 1.8401e-19 $X=2.25 $Y=1.34
r194 94 95 9.82337 $w=3.68e-07 $l=7.5e-08 $layer=POLY_cond $X=7.515 $Y=1.542
+ $X2=7.59 $Y2=1.542
r195 93 94 46.4973 $w=3.68e-07 $l=3.55e-07 $layer=POLY_cond $X=7.16 $Y=1.542
+ $X2=7.515 $Y2=1.542
r196 92 93 12.4429 $w=3.68e-07 $l=9.5e-08 $layer=POLY_cond $X=7.065 $Y=1.542
+ $X2=7.16 $Y2=1.542
r197 89 90 15.0625 $w=3.68e-07 $l=1.15e-07 $layer=POLY_cond $X=6.615 $Y=1.542
+ $X2=6.73 $Y2=1.542
r198 88 89 41.2582 $w=3.68e-07 $l=3.15e-07 $layer=POLY_cond $X=6.3 $Y=1.542
+ $X2=6.615 $Y2=1.542
r199 78 80 0.122819 $w=2.98e-07 $l=3e-09 $layer=LI1_cond $X=4.07 $Y=1.907
+ $X2=4.07 $Y2=1.91
r200 77 78 13.7966 $w=2.98e-07 $l=3.37e-07 $layer=LI1_cond $X=4.07 $Y=1.57
+ $X2=4.07 $Y2=1.907
r201 75 92 36.019 $w=3.68e-07 $l=2.75e-07 $layer=POLY_cond $X=6.79 $Y=1.542
+ $X2=7.065 $Y2=1.542
r202 75 90 7.8587 $w=3.68e-07 $l=6e-08 $layer=POLY_cond $X=6.79 $Y=1.542
+ $X2=6.73 $Y2=1.542
r203 74 75 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.79
+ $Y=1.485 $X2=6.79 $Y2=1.485
r204 72 88 24.8859 $w=3.68e-07 $l=1.9e-07 $layer=POLY_cond $X=6.11 $Y=1.542
+ $X2=6.3 $Y2=1.542
r205 72 86 13.7527 $w=3.68e-07 $l=1.05e-07 $layer=POLY_cond $X=6.11 $Y=1.542
+ $X2=6.005 $Y2=1.542
r206 71 74 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.11 $Y=1.485
+ $X2=6.79 $Y2=1.485
r207 71 72 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.11
+ $Y=1.485 $X2=6.11 $Y2=1.485
r208 69 71 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=6.05 $Y=1.485
+ $X2=6.11 $Y2=1.485
r209 67 69 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.965 $Y=1.65
+ $X2=6.05 $Y2=1.485
r210 67 68 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.965 $Y=1.65
+ $X2=5.965 $Y2=1.82
r211 66 81 8.29065 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.12 $Y=1.985
+ $X2=4.955 $Y2=1.985
r212 63 68 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.88 $Y=1.985
+ $X2=5.965 $Y2=1.82
r213 63 66 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=5.88 $Y=1.985
+ $X2=5.12 $Y2=1.985
r214 62 78 3.87205 $w=1.75e-07 $l=1.6e-07 $layer=LI1_cond $X=4.23 $Y=1.907
+ $X2=4.07 $Y2=1.907
r215 62 81 45.9481 $w=1.73e-07 $l=7.25e-07 $layer=LI1_cond $X=4.23 $Y=1.907
+ $X2=4.955 $Y2=1.907
r216 57 77 6.24057 $w=3.3e-07 $l=1.86145e-07 $layer=LI1_cond $X=4.115 $Y=1.405
+ $X2=4.07 $Y2=1.57
r217 57 59 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=4.115 $Y=1.405
+ $X2=4.115 $Y2=0.74
r218 55 85 9.19847 $w=3.93e-07 $l=7.5e-08 $layer=POLY_cond $X=3.24 $Y=1.58
+ $X2=3.315 $Y2=1.58
r219 55 83 45.9924 $w=3.93e-07 $l=3.75e-07 $layer=POLY_cond $X=3.24 $Y=1.58
+ $X2=2.865 $Y2=1.58
r220 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.24
+ $Y=1.57 $X2=3.24 $Y2=1.57
r221 52 77 0.0845041 $w=3.3e-07 $l=1.7e-07 $layer=LI1_cond $X=3.9 $Y=1.57
+ $X2=4.07 $Y2=1.57
r222 52 54 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=3.9 $Y=1.57
+ $X2=3.24 $Y2=1.57
r223 48 95 23.8357 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=7.59 $Y=1.32
+ $X2=7.59 $Y2=1.542
r224 48 50 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.59 $Y=1.32
+ $X2=7.59 $Y2=0.74
r225 45 94 23.8357 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.515 $Y=1.765
+ $X2=7.515 $Y2=1.542
r226 45 47 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.515 $Y=1.765
+ $X2=7.515 $Y2=2.4
r227 41 93 23.8357 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=7.16 $Y=1.32
+ $X2=7.16 $Y2=1.542
r228 41 43 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.16 $Y=1.32
+ $X2=7.16 $Y2=0.74
r229 38 92 23.8357 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.065 $Y=1.765
+ $X2=7.065 $Y2=1.542
r230 38 40 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.065 $Y=1.765
+ $X2=7.065 $Y2=2.4
r231 34 90 23.8357 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.73 $Y=1.32
+ $X2=6.73 $Y2=1.542
r232 34 36 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.73 $Y=1.32
+ $X2=6.73 $Y2=0.74
r233 31 89 23.8357 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.615 $Y=1.765
+ $X2=6.615 $Y2=1.542
r234 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.615 $Y=1.765
+ $X2=6.615 $Y2=2.4
r235 27 88 23.8357 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.3 $Y=1.32
+ $X2=6.3 $Y2=1.542
r236 27 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.3 $Y=1.32 $X2=6.3
+ $Y2=0.74
r237 24 86 23.8357 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.005 $Y=1.765
+ $X2=6.005 $Y2=1.542
r238 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.005 $Y=1.765
+ $X2=6.005 $Y2=2.4
r239 21 85 25.4309 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.315 $Y=1.82
+ $X2=3.315 $Y2=1.58
r240 21 23 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.315 $Y=1.82
+ $X2=3.315 $Y2=2.315
r241 18 83 25.4309 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.865 $Y=1.82
+ $X2=2.865 $Y2=1.58
r242 18 20 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.865 $Y=1.82
+ $X2=2.865 $Y2=2.315
r243 15 83 17.7837 $w=3.93e-07 $l=3.03974e-07 $layer=POLY_cond $X=2.72 $Y=1.34
+ $X2=2.865 $Y2=1.58
r244 15 17 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.72 $Y=1.34
+ $X2=2.72 $Y2=0.945
r245 13 15 28.4128 $w=3.93e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.645 $Y=1.415
+ $X2=2.72 $Y2=1.34
r246 13 14 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.645 $Y=1.415
+ $X2=2.325 $Y2=1.415
r247 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.25 $Y=1.34
+ $X2=2.325 $Y2=1.415
r248 10 12 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.25 $Y=1.34
+ $X2=2.25 $Y2=0.945
r249 3 66 600 $w=1.7e-07 $l=2.55441e-07 $layer=licon1_PDIFF $count=1 $X=4.895
+ $Y=2.05 $X2=5.12 $Y2=1.985
r250 2 80 600 $w=1.7e-07 $l=2.32379e-07 $layer=licon1_PDIFF $count=1 $X=3.84
+ $Y=1.895 $X2=4.065 $Y2=1.91
r251 1 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.975
+ $Y=0.595 $X2=4.115 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__HA_4%B 3 5 7 10 12 14 15 16 18 19 20 21 22 23 26 29
+ 31 33 37 39 41 43 44 46 47
c135 47 0 1.898e-19 $X=2.16 $Y=1.665
c136 23 0 1.26877e-19 $X=3.765 $Y=1.82
c137 12 0 7.21125e-20 $X=1.845 $Y=1.885
c138 3 0 1.44963e-19 $X=1.36 $Y=0.945
r139 55 56 6.32697 $w=4.19e-07 $l=5.5e-08 $layer=POLY_cond $X=1.79 $Y=1.67
+ $X2=1.845 $Y2=1.67
r140 53 55 6.90215 $w=4.19e-07 $l=6e-08 $layer=POLY_cond $X=1.73 $Y=1.67
+ $X2=1.79 $Y2=1.67
r141 51 53 38.537 $w=4.19e-07 $l=3.35e-07 $layer=POLY_cond $X=1.395 $Y=1.67
+ $X2=1.73 $Y2=1.67
r142 50 51 4.02625 $w=4.19e-07 $l=3.5e-08 $layer=POLY_cond $X=1.36 $Y=1.67
+ $X2=1.395 $Y2=1.67
r143 46 47 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.62
+ $X2=2.16 $Y2=1.62
r144 46 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.62 $X2=1.73 $Y2=1.62
r145 39 44 74.0611 $w=1.8e-07 $l=1.85e-07 $layer=POLY_cond $X=4.37 $Y=2.965
+ $X2=4.37 $Y2=3.15
r146 39 41 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.37 $Y=2.965
+ $X2=4.37 $Y2=2.47
r147 35 37 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=4.33 $Y=1.53
+ $X2=4.33 $Y2=0.915
r148 34 42 13.9682 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.975 $Y=1.605
+ $X2=3.825 $Y2=1.605
r149 33 35 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.255 $Y=1.605
+ $X2=4.33 $Y2=1.53
r150 33 34 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.255 $Y=1.605
+ $X2=3.975 $Y2=1.605
r151 32 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.855 $Y=3.15
+ $X2=3.765 $Y2=3.15
r152 31 44 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.28 $Y=3.15 $X2=4.37
+ $Y2=3.15
r153 31 32 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.28 $Y=3.15
+ $X2=3.855 $Y2=3.15
r154 27 42 21.8618 $w=2.42e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.9 $Y=1.53
+ $X2=3.825 $Y2=1.605
r155 27 29 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.9 $Y=1.53
+ $X2=3.9 $Y2=0.915
r156 24 26 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.765 $Y=2.81
+ $X2=3.765 $Y2=2.315
r157 23 42 49.7461 $w=2.42e-07 $l=2.43156e-07 $layer=POLY_cond $X=3.765 $Y=1.82
+ $X2=3.825 $Y2=1.605
r158 23 26 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.765 $Y=1.82
+ $X2=3.765 $Y2=2.315
r159 22 43 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=3.075
+ $X2=3.765 $Y2=3.15
r160 21 24 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.765 $Y=2.9
+ $X2=3.765 $Y2=2.81
r161 21 22 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.765 $Y=2.9
+ $X2=3.765 $Y2=3.075
r162 19 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.675 $Y=3.15
+ $X2=3.765 $Y2=3.15
r163 19 20 638.394 $w=1.5e-07 $l=1.245e-06 $layer=POLY_cond $X=3.675 $Y=3.15
+ $X2=2.43 $Y2=3.15
r164 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.355 $Y=3.075
+ $X2=2.43 $Y2=3.15
r165 17 18 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=2.355 $Y=1.88
+ $X2=2.355 $Y2=3.075
r166 16 56 31.3489 $w=4.19e-07 $l=1.74284e-07 $layer=POLY_cond $X=1.935 $Y=1.805
+ $X2=1.845 $Y2=1.67
r167 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.28 $Y=1.805
+ $X2=2.355 $Y2=1.88
r168 15 16 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.28 $Y=1.805
+ $X2=1.935 $Y2=1.805
r169 12 56 27.0004 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.845 $Y=1.885
+ $X2=1.845 $Y2=1.67
r170 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.845 $Y=1.885
+ $X2=1.845 $Y2=2.46
r171 8 55 27.0004 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.79 $Y=1.455
+ $X2=1.79 $Y2=1.67
r172 8 10 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.79 $Y=1.455
+ $X2=1.79 $Y2=0.945
r173 5 51 27.0004 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.395 $Y=1.885
+ $X2=1.395 $Y2=1.67
r174 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.395 $Y=1.885
+ $X2=1.395 $Y2=2.46
r175 1 50 27.0004 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.36 $Y=1.455
+ $X2=1.36 $Y2=1.67
r176 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.36 $Y=1.455
+ $X2=1.36 $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_LS__HA_4%A 3 5 7 11 12 14 15 16 18 19 21 25 26 28 30 31
+ 33 34 35 36 37 38 46
c118 46 0 1.898e-19 $X=0.93 $Y=1.67
c119 28 0 1.39181e-20 $X=5.33 $Y=1.31
c120 12 0 5.25684e-20 $X=0.945 $Y=1.885
c121 5 0 2.13006e-19 $X=0.495 $Y=1.885
r122 46 47 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=0.93 $Y=1.67
+ $X2=0.945 $Y2=1.67
r123 44 46 26.1402 $w=3.78e-07 $l=2.05e-07 $layer=POLY_cond $X=0.725 $Y=1.67
+ $X2=0.93 $Y2=1.67
r124 42 44 29.328 $w=3.78e-07 $l=2.3e-07 $layer=POLY_cond $X=0.495 $Y=1.67
+ $X2=0.725 $Y2=1.67
r125 37 38 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.62
+ $X2=1.2 $Y2=1.62
r126 37 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.725
+ $Y=1.62 $X2=0.725 $Y2=1.62
r127 36 37 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.62
+ $X2=0.72 $Y2=1.62
r128 31 35 36.308 $w=1.5e-07 $l=4.97971e-07 $layer=POLY_cond $X=5.345 $Y=1.765
+ $X2=5.255 $Y2=1.31
r129 31 33 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.345 $Y=1.765
+ $X2=5.345 $Y2=2.26
r130 28 35 36.308 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.33 $Y=1.31
+ $X2=5.255 $Y2=1.31
r131 28 30 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.33 $Y=1.31
+ $X2=5.33 $Y2=0.915
r132 27 34 3.5291 $w=3.2e-07 $l=1.84932e-07 $layer=POLY_cond $X=4.91 $Y=1.47
+ $X2=4.73 $Y2=1.46
r133 26 35 4.67038 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=5.255 $Y=1.47
+ $X2=5.255 $Y2=1.31
r134 26 27 62.2124 $w=3.2e-07 $l=3.45e-07 $layer=POLY_cond $X=5.255 $Y=1.47
+ $X2=4.91 $Y2=1.47
r135 23 34 33.9972 $w=1.65e-07 $l=1.93649e-07 $layer=POLY_cond $X=4.83 $Y=1.31
+ $X2=4.73 $Y2=1.46
r136 23 25 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.83 $Y=1.31
+ $X2=4.83 $Y2=0.915
r137 22 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.83 $Y=0.255
+ $X2=4.83 $Y2=0.915
r138 19 21 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.82 $Y=1.975
+ $X2=4.82 $Y2=2.47
r139 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.82 $Y=1.885
+ $X2=4.82 $Y2=1.975
r140 17 34 33.9972 $w=1.65e-07 $l=2.10238e-07 $layer=POLY_cond $X=4.82 $Y=1.63
+ $X2=4.73 $Y2=1.46
r141 17 18 99.121 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=4.82 $Y=1.63
+ $X2=4.82 $Y2=1.885
r142 15 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.755 $Y=0.18
+ $X2=4.83 $Y2=0.255
r143 15 16 1922.87 $w=1.5e-07 $l=3.75e-06 $layer=POLY_cond $X=4.755 $Y=0.18
+ $X2=1.005 $Y2=0.18
r144 12 47 24.4846 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.945 $Y=1.885
+ $X2=0.945 $Y2=1.67
r145 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.945 $Y=1.885
+ $X2=0.945 $Y2=2.46
r146 9 46 24.4846 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.93 $Y=1.455
+ $X2=0.93 $Y2=1.67
r147 9 11 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.93 $Y=1.455
+ $X2=0.93 $Y2=0.945
r148 8 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.93 $Y=0.255
+ $X2=1.005 $Y2=0.18
r149 8 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.93 $Y=0.255
+ $X2=0.93 $Y2=0.945
r150 5 42 24.4846 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.495 $Y=1.885
+ $X2=0.495 $Y2=1.67
r151 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.885
+ $X2=0.495 $Y2=2.46
r152 1 42 24.4846 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.495 $Y=1.455
+ $X2=0.495 $Y2=1.67
r153 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.495 $Y=1.455
+ $X2=0.495 $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_LS__HA_4%A_294_392# 1 2 3 10 12 15 17 19 22 24 26 29 31
+ 32 35 37 39 42 46 49 50 52 54 57 58 63 64 67 68 69 72 74
c205 67 0 5.25684e-20 $X=1.62 $Y=2.12
c206 57 0 5.29972e-20 $X=7.81 $Y=2.32
c207 52 0 1.26877e-19 $X=3.9 $Y=2.25
c208 49 0 1.0136e-19 $X=2.585 $Y=1.905
c209 32 0 9.44376e-20 $X=9.025 $Y=1.485
c210 10 0 2.24074e-19 $X=7.965 $Y=1.765
r211 83 84 10.6693 $w=3.84e-07 $l=8.5e-08 $layer=POLY_cond $X=8.865 $Y=1.542
+ $X2=8.95 $Y2=1.542
r212 82 83 52.0911 $w=3.84e-07 $l=4.15e-07 $layer=POLY_cond $X=8.45 $Y=1.542
+ $X2=8.865 $Y2=1.542
r213 81 82 4.39323 $w=3.84e-07 $l=3.5e-08 $layer=POLY_cond $X=8.415 $Y=1.542
+ $X2=8.45 $Y2=1.542
r214 78 79 6.90365 $w=3.84e-07 $l=5.5e-08 $layer=POLY_cond $X=7.965 $Y=1.542
+ $X2=8.02 $Y2=1.542
r215 74 76 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.985 $Y=2.25
+ $X2=3.985 $Y2=2.405
r216 72 73 7.52055 $w=2.92e-07 $l=1.8e-07 $layer=LI1_cond $X=3.09 $Y=2.07
+ $X2=3.09 $Y2=2.25
r217 70 72 2.29795 $w=2.92e-07 $l=5.5e-08 $layer=LI1_cond $X=3.09 $Y=2.015
+ $X2=3.09 $Y2=2.07
r218 64 87 1.8075 $w=4e-07 $l=1.5e-08 $layer=POLY_cond $X=9.56 $Y=1.542
+ $X2=9.575 $Y2=1.542
r219 64 85 6.6275 $w=4e-07 $l=5.5e-08 $layer=POLY_cond $X=9.56 $Y=1.542
+ $X2=9.505 $Y2=1.542
r220 63 64 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=9.56
+ $Y=1.485 $X2=9.56 $Y2=1.485
r221 61 81 47.0703 $w=3.84e-07 $l=3.75e-07 $layer=POLY_cond $X=8.04 $Y=1.542
+ $X2=8.415 $Y2=1.542
r222 61 79 2.51042 $w=3.84e-07 $l=2e-08 $layer=POLY_cond $X=8.04 $Y=1.542
+ $X2=8.02 $Y2=1.542
r223 60 63 53.0822 $w=3.28e-07 $l=1.52e-06 $layer=LI1_cond $X=8.04 $Y=1.485
+ $X2=9.56 $Y2=1.485
r224 60 61 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=8.04
+ $Y=1.485 $X2=8.04 $Y2=1.485
r225 58 60 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=7.895 $Y=1.485
+ $X2=8.04 $Y2=1.485
r226 56 58 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.81 $Y=1.65
+ $X2=7.895 $Y2=1.485
r227 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.81 $Y=1.65
+ $X2=7.81 $Y2=2.32
r228 55 76 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=2.405
+ $X2=3.985 $Y2=2.405
r229 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.725 $Y=2.405
+ $X2=7.81 $Y2=2.32
r230 54 55 238.455 $w=1.68e-07 $l=3.655e-06 $layer=LI1_cond $X=7.725 $Y=2.405
+ $X2=4.07 $Y2=2.405
r231 53 73 3.90229 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=2.25
+ $X2=3.09 $Y2=2.25
r232 52 74 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.9 $Y=2.25
+ $X2=3.985 $Y2=2.25
r233 52 53 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.9 $Y=2.25
+ $X2=3.255 $Y2=2.25
r234 51 69 4.60183 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=2.015
+ $X2=2.585 $Y2=2.015
r235 50 70 2.3974 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=2.015
+ $X2=3.09 $Y2=2.015
r236 50 51 13.3579 $w=2.18e-07 $l=2.55e-07 $layer=LI1_cond $X=2.925 $Y=2.015
+ $X2=2.67 $Y2=2.015
r237 49 69 1.84097 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.585 $Y=1.905
+ $X2=2.585 $Y2=2.015
r238 49 68 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.585 $Y=1.905
+ $X2=2.585 $Y2=1.285
r239 44 68 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=1.12
+ $X2=2.505 $Y2=1.285
r240 44 46 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=2.505 $Y=1.12
+ $X2=2.505 $Y2=0.77
r241 43 67 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.735 $Y=2.04
+ $X2=1.595 $Y2=2.04
r242 42 69 4.60183 $w=1.95e-07 $l=9.66954e-08 $layer=LI1_cond $X=2.5 $Y=2.04
+ $X2=2.585 $Y2=2.015
r243 42 43 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.5 $Y=2.04
+ $X2=1.735 $Y2=2.04
r244 37 87 25.8619 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=9.575 $Y=1.765
+ $X2=9.575 $Y2=1.542
r245 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.575 $Y=1.765
+ $X2=9.575 $Y2=2.4
r246 33 85 25.8619 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=9.505 $Y=1.32
+ $X2=9.505 $Y2=1.542
r247 33 35 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.505 $Y=1.32
+ $X2=9.505 $Y2=0.74
r248 32 84 10.5016 $w=3.84e-07 $l=9.94987e-08 $layer=POLY_cond $X=9.025 $Y=1.485
+ $X2=8.95 $Y2=1.542
r249 31 85 10.6563 $w=4e-07 $l=9.94987e-08 $layer=POLY_cond $X=9.43 $Y=1.485
+ $X2=9.505 $Y2=1.542
r250 31 32 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=9.43 $Y=1.485
+ $X2=9.025 $Y2=1.485
r251 27 84 24.8669 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=8.95 $Y=1.32
+ $X2=8.95 $Y2=1.542
r252 27 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.95 $Y=1.32
+ $X2=8.95 $Y2=0.74
r253 24 83 24.8669 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=8.865 $Y=1.765
+ $X2=8.865 $Y2=1.542
r254 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.865 $Y=1.765
+ $X2=8.865 $Y2=2.4
r255 20 82 24.8669 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=8.45 $Y=1.32
+ $X2=8.45 $Y2=1.542
r256 20 22 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.45 $Y=1.32
+ $X2=8.45 $Y2=0.74
r257 17 81 24.8669 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=8.415 $Y=1.765
+ $X2=8.415 $Y2=1.542
r258 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.415 $Y=1.765
+ $X2=8.415 $Y2=2.4
r259 13 79 24.8669 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=8.02 $Y=1.32
+ $X2=8.02 $Y2=1.542
r260 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.02 $Y=1.32
+ $X2=8.02 $Y2=0.74
r261 10 78 24.8669 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.965 $Y=1.765
+ $X2=7.965 $Y2=1.542
r262 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.965 $Y=1.765
+ $X2=7.965 $Y2=2.4
r263 3 72 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.895 $X2=3.09 $Y2=2.07
r264 2 67 300 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=2 $X=1.47
+ $Y=1.96 $X2=1.62 $Y2=2.12
r265 1 46 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=2.325
+ $Y=0.625 $X2=2.505 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LS__HA_4%A_27_392# 1 2 3 10 12 14 16 19 20 21 24
c44 21 0 1.02086e-19 $X=1.255 $Y=2.99
c45 12 0 1.10921e-19 $X=0.27 $Y=2.8
r46 22 24 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=2.07 $Y=2.905
+ $X2=2.07 $Y2=2.38
r47 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.905 $Y=2.99
+ $X2=2.07 $Y2=2.905
r48 20 21 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.905 $Y=2.99
+ $X2=1.255 $Y2=2.99
r49 17 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.13 $Y=2.905
+ $X2=1.255 $Y2=2.99
r50 17 19 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.13 $Y=2.905 $X2=1.13
+ $Y2=2.815
r51 16 29 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=2.125
+ $X2=1.13 $Y2=2.04
r52 16 19 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=1.13 $Y=2.125
+ $X2=1.13 $Y2=2.815
r53 15 27 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.385 $Y=2.04
+ $X2=0.245 $Y2=2.04
r54 14 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.005 $Y=2.04
+ $X2=1.13 $Y2=2.04
r55 14 15 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.005 $Y=2.04
+ $X2=0.385 $Y2=2.04
r56 10 27 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=2.125
+ $X2=0.245 $Y2=2.04
r57 10 12 27.7821 $w=2.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.245 $Y=2.125
+ $X2=0.245 $Y2=2.8
r58 3 24 300 $w=1.7e-07 $l=4.89285e-07 $layer=licon1_PDIFF $count=2 $X=1.92
+ $Y=1.96 $X2=2.07 $Y2=2.38
r59 2 29 400 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.96 $X2=1.17 $Y2=2.12
r60 2 19 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.96 $X2=1.17 $Y2=2.815
r61 1 27 400 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.27 $Y2=2.12
r62 1 12 400 $w=1.7e-07 $l=9.04986e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.27 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_LS__HA_4%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 44 48 52 56
+ 60 62 64 67 68 70 71 73 74 75 77 82 90 95 110 115 118 121 124 127 131
c157 34 0 7.21125e-20 $X=2.64 $Y=2.57
c158 2 0 1.0136e-19 $X=2.505 $Y=1.895
r159 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r160 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r161 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r162 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r163 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r164 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r165 113 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r166 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r167 110 130 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=9.635 $Y=3.33
+ $X2=9.857 $Y2=3.33
r168 110 112 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.635 $Y=3.33
+ $X2=9.36 $Y2=3.33
r169 109 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r170 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r171 106 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r172 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r173 103 106 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r174 103 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=5.52 $Y2=3.33
r175 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r176 100 127 10.6558 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=5.945 $Y=3.33
+ $X2=5.717 $Y2=3.33
r177 100 102 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=5.945 $Y=3.33
+ $X2=6.48 $Y2=3.33
r178 99 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r179 99 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r180 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r181 96 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.54 $Y2=3.33
r182 96 98 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r183 95 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.595 $Y2=3.33
r184 95 98 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.08 $Y2=3.33
r185 94 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r186 94 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r187 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r188 91 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.64 $Y2=3.33
r189 91 93 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=3.12 $Y2=3.33
r190 90 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.54 $Y2=3.33
r191 90 93 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.12 $Y2=3.33
r192 89 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r193 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r194 86 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r195 86 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r196 85 88 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r197 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r198 83 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.68 $Y2=3.33
r199 83 85 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.2 $Y2=3.33
r200 82 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=3.33
+ $X2=2.64 $Y2=3.33
r201 82 88 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.475 $Y=3.33
+ $X2=2.16 $Y2=3.33
r202 80 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r203 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r204 77 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.68 $Y2=3.33
r205 77 79 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r206 75 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r207 75 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r208 73 108 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=8.475 $Y=3.33
+ $X2=8.4 $Y2=3.33
r209 73 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.475 $Y=3.33
+ $X2=8.64 $Y2=3.33
r210 72 112 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=8.805 $Y=3.33
+ $X2=9.36 $Y2=3.33
r211 72 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.805 $Y=3.33
+ $X2=8.64 $Y2=3.33
r212 70 105 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.575 $Y=3.33
+ $X2=7.44 $Y2=3.33
r213 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.575 $Y=3.33
+ $X2=7.74 $Y2=3.33
r214 69 108 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.905 $Y=3.33
+ $X2=8.4 $Y2=3.33
r215 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.905 $Y=3.33
+ $X2=7.74 $Y2=3.33
r216 67 102 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.675 $Y=3.33
+ $X2=6.48 $Y2=3.33
r217 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=3.33
+ $X2=6.84 $Y2=3.33
r218 66 105 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.005 $Y=3.33
+ $X2=7.44 $Y2=3.33
r219 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.005 $Y=3.33
+ $X2=6.84 $Y2=3.33
r220 62 130 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.8 $Y=3.245
+ $X2=9.857 $Y2=3.33
r221 62 64 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=9.8 $Y=3.245
+ $X2=9.8 $Y2=2.415
r222 58 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.64 $Y=3.245
+ $X2=8.64 $Y2=3.33
r223 58 60 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=8.64 $Y=3.245
+ $X2=8.64 $Y2=2.405
r224 54 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.74 $Y=3.245
+ $X2=7.74 $Y2=3.33
r225 54 56 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.74 $Y=3.245
+ $X2=7.74 $Y2=2.78
r226 50 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=3.245
+ $X2=6.84 $Y2=3.33
r227 50 52 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.84 $Y=3.245
+ $X2=6.84 $Y2=2.78
r228 46 127 1.82608 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=5.717 $Y=3.245
+ $X2=5.717 $Y2=3.33
r229 46 48 13.1437 $w=4.53e-07 $l=5e-07 $layer=LI1_cond $X=5.717 $Y=3.245
+ $X2=5.717 $Y2=2.745
r230 45 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.76 $Y=3.33
+ $X2=4.595 $Y2=3.33
r231 44 127 10.6558 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=5.49 $Y=3.33
+ $X2=5.717 $Y2=3.33
r232 44 45 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.49 $Y=3.33
+ $X2=4.76 $Y2=3.33
r233 40 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.595 $Y=3.245
+ $X2=4.595 $Y2=3.33
r234 40 42 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.595 $Y=3.245
+ $X2=4.595 $Y2=2.745
r235 36 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=3.245
+ $X2=3.54 $Y2=3.33
r236 36 38 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=3.54 $Y=3.245
+ $X2=3.54 $Y2=2.59
r237 32 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=3.245
+ $X2=2.64 $Y2=3.33
r238 32 34 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.64 $Y=3.245
+ $X2=2.64 $Y2=2.57
r239 28 115 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=3.245
+ $X2=0.68 $Y2=3.33
r240 28 30 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=0.68 $Y=3.245
+ $X2=0.68 $Y2=2.46
r241 9 64 300 $w=1.7e-07 $l=6.45659e-07 $layer=licon1_PDIFF $count=2 $X=9.65
+ $Y=1.84 $X2=9.8 $Y2=2.415
r242 8 60 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=8.49
+ $Y=1.84 $X2=8.64 $Y2=2.405
r243 7 56 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=7.59
+ $Y=1.84 $X2=7.74 $Y2=2.78
r244 6 52 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=6.69
+ $Y=1.84 $X2=6.84 $Y2=2.78
r245 5 48 600 $w=1.7e-07 $l=1.04211e-06 $layer=licon1_PDIFF $count=1 $X=5.42
+ $Y=1.84 $X2=5.715 $Y2=2.745
r246 4 42 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=4.445
+ $Y=2.05 $X2=4.595 $Y2=2.745
r247 3 38 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=3.39
+ $Y=1.895 $X2=3.54 $Y2=2.59
r248 2 34 600 $w=1.7e-07 $l=7.39425e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=1.895 $X2=2.64 $Y2=2.57
r249 1 30 300 $w=1.7e-07 $l=5.70088e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.96 $X2=0.72 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__HA_4%COUT 1 2 3 4 13 17 19 21 25 28 29 30 34
c51 28 0 1.49079e-19 $X=7.44 $Y=1.295
r52 30 34 3.3396 $w=3.45e-07 $l=1.65e-07 $layer=LI1_cond $X=7.382 $Y=1.985
+ $X2=7.382 $Y2=1.82
r53 29 34 5.17764 $w=3.43e-07 $l=1.55e-07 $layer=LI1_cond $X=7.382 $Y=1.665
+ $X2=7.382 $Y2=1.82
r54 28 29 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=7.382 $Y=1.295
+ $X2=7.382 $Y2=1.665
r55 25 28 5.51168 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=7.382 $Y=1.13
+ $X2=7.382 $Y2=1.295
r56 25 27 2.96505 $w=3.45e-07 $l=1.25e-07 $layer=LI1_cond $X=7.382 $Y=1.13
+ $X2=7.382 $Y2=1.005
r57 22 24 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.6 $Y=1.005
+ $X2=6.475 $Y2=1.005
r58 21 27 4.07991 $w=2.5e-07 $l=1.72e-07 $layer=LI1_cond $X=7.21 $Y=1.005
+ $X2=7.382 $Y2=1.005
r59 21 22 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=7.21 $Y=1.005
+ $X2=6.6 $Y2=1.005
r60 17 24 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.475 $Y=0.88
+ $X2=6.475 $Y2=1.005
r61 17 19 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=6.475 $Y=0.88
+ $X2=6.475 $Y2=0.515
r62 13 30 3.48128 $w=3.3e-07 $l=1.72e-07 $layer=LI1_cond $X=7.21 $Y=1.985
+ $X2=7.382 $Y2=1.985
r63 13 15 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=7.21 $Y=1.985
+ $X2=6.385 $Y2=1.985
r64 4 30 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.14
+ $Y=1.84 $X2=7.29 $Y2=1.985
r65 3 15 600 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=1 $X=6.08
+ $Y=1.84 $X2=6.385 $Y2=1.985
r66 2 27 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.235
+ $Y=0.37 $X2=7.375 $Y2=0.965
r67 1 24 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=6.375
+ $Y=0.37 $X2=6.515 $Y2=0.965
r68 1 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.375
+ $Y=0.37 $X2=6.515 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__HA_4%SUM 1 2 3 4 13 15 19 21 22 25 29 31 33 36 40 41
+ 43 44 45 50
c89 13 0 1.74057e-19 $X=8.19 $Y=2.15
r90 50 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=2.035
+ $X2=9.84 $Y2=2.035
r91 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=2.035
+ $X2=8.88 $Y2=2.035
r92 45 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.025 $Y=2.035
+ $X2=8.88 $Y2=2.035
r93 44 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.695 $Y=2.035
+ $X2=9.84 $Y2=2.035
r94 44 45 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=9.695 $Y=2.035
+ $X2=9.025 $Y2=2.035
r95 41 48 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=9.075 $Y=1.985
+ $X2=8.88 $Y2=1.985
r96 41 43 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.075 $Y=1.985
+ $X2=9.24 $Y2=1.985
r97 37 48 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=8.305 $Y=1.985
+ $X2=8.88 $Y2=1.985
r98 37 39 2.91733 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=8.305 $Y=1.985
+ $X2=8.19 $Y2=1.985
r99 36 54 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.91 $Y=1.82
+ $X2=9.91 $Y2=1.985
r100 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.91 $Y=1.15
+ $X2=9.91 $Y2=1.82
r101 34 43 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.405 $Y=1.985
+ $X2=9.24 $Y2=1.985
r102 33 54 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.825 $Y=1.985
+ $X2=9.91 $Y2=1.985
r103 33 34 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=9.825 $Y=1.985
+ $X2=9.405 $Y2=1.985
r104 32 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.4 $Y=1.065
+ $X2=9.235 $Y2=1.065
r105 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.825 $Y=1.065
+ $X2=9.91 $Y2=1.15
r106 31 32 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.825 $Y=1.065
+ $X2=9.4 $Y2=1.065
r107 27 43 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.24 $Y=2.15
+ $X2=9.24 $Y2=1.985
r108 27 29 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=9.24 $Y=2.15
+ $X2=9.24 $Y2=2.43
r109 23 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.235 $Y=0.98
+ $X2=9.235 $Y2=1.065
r110 23 25 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=9.235 $Y=0.98
+ $X2=9.235 $Y2=0.515
r111 21 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.07 $Y=1.065
+ $X2=9.235 $Y2=1.065
r112 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.07 $Y=1.065
+ $X2=8.4 $Y2=1.065
r113 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.275 $Y=0.98
+ $X2=8.4 $Y2=1.065
r114 17 19 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=8.275 $Y=0.98
+ $X2=8.275 $Y2=0.515
r115 13 39 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.19 $Y=2.15
+ $X2=8.19 $Y2=1.985
r116 13 15 14.0297 $w=2.28e-07 $l=2.8e-07 $layer=LI1_cond $X=8.19 $Y=2.15
+ $X2=8.19 $Y2=2.43
r117 4 43 600 $w=1.7e-07 $l=3.65377e-07 $layer=licon1_PDIFF $count=1 $X=8.94
+ $Y=1.84 $X2=9.24 $Y2=1.985
r118 4 29 300 $w=1.7e-07 $l=7.24638e-07 $layer=licon1_PDIFF $count=2 $X=8.94
+ $Y=1.84 $X2=9.24 $Y2=2.43
r119 3 39 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.04
+ $Y=1.84 $X2=8.19 $Y2=1.985
r120 3 15 300 $w=1.7e-07 $l=6.60757e-07 $layer=licon1_PDIFF $count=2 $X=8.04
+ $Y=1.84 $X2=8.19 $Y2=2.43
r121 2 25 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=9.025
+ $Y=0.37 $X2=9.235 $Y2=0.515
r122 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.095
+ $Y=0.37 $X2=8.235 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__HA_4%A_27_125# 1 2 3 4 15 17 18 21 23 28 29 30 33 35
c66 23 0 1.8401e-19 $X=1.84 $Y=1.2
c67 21 0 1.44963e-19 $X=1.145 $Y=0.77
r68 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.005 $Y=0.435
+ $X2=3.005 $Y2=0.77
r69 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.84 $Y=0.35
+ $X2=3.005 $Y2=0.435
r70 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.84 $Y=0.35
+ $X2=2.17 $Y2=0.35
r71 26 28 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.005 $Y=1.115
+ $X2=2.005 $Y2=0.77
r72 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.005 $Y=0.435
+ $X2=2.17 $Y2=0.35
r73 25 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.005 $Y=0.435
+ $X2=2.005 $Y2=0.77
r74 24 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.23 $Y=1.2
+ $X2=1.105 $Y2=1.2
r75 23 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.84 $Y=1.2
+ $X2=2.005 $Y2=1.115
r76 23 24 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.84 $Y=1.2 $X2=1.23
+ $Y2=1.2
r77 19 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.105 $Y=1.115
+ $X2=1.105 $Y2=1.2
r78 19 21 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=1.105 $Y=1.115
+ $X2=1.105 $Y2=0.77
r79 17 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.98 $Y=1.2
+ $X2=1.105 $Y2=1.2
r80 17 18 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.98 $Y=1.2
+ $X2=0.365 $Y2=1.2
r81 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.115
+ $X2=0.365 $Y2=1.2
r82 13 15 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.115
+ $X2=0.24 $Y2=0.77
r83 4 33 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.795
+ $Y=0.625 $X2=3.005 $Y2=0.77
r84 3 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.865
+ $Y=0.625 $X2=2.005 $Y2=0.77
r85 2 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.005
+ $Y=0.625 $X2=1.145 $Y2=0.77
r86 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.625 $X2=0.28 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LS__HA_4%VGND 1 2 3 4 5 6 7 8 27 31 35 37 41 45 49 53 55
+ 57 60 61 63 64 66 67 69 70 71 80 87 99 104 107 110 114
c126 49 0 9.44376e-20 $X=7.805 $Y=0.53
r127 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r128 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r129 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r130 102 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r131 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r132 99 113 4.36388 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=9.58 $Y=0 $X2=9.83
+ $Y2=0
r133 99 101 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=9.58 $Y=0 $X2=9.36
+ $Y2=0
r134 98 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r135 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r136 95 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r137 95 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r138 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r139 92 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.11 $Y=0
+ $X2=6.945 $Y2=0
r140 92 94 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.11 $Y=0 $X2=7.44
+ $Y2=0
r141 91 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r142 91 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r143 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r144 88 107 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.17 $Y=0
+ $X2=6.045 $Y2=0
r145 88 90 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.17 $Y=0 $X2=6.48
+ $Y2=0
r146 87 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.78 $Y=0
+ $X2=6.945 $Y2=0
r147 87 90 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.78 $Y=0 $X2=6.48
+ $Y2=0
r148 85 86 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r149 83 86 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=4.56 $Y2=0
r150 82 85 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=4.56
+ $Y2=0
r151 82 83 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r152 80 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.95 $Y=0
+ $X2=5.115 $Y2=0
r153 80 85 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.95 $Y=0 $X2=4.56
+ $Y2=0
r154 79 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r155 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r156 75 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r157 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r158 71 108 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r159 71 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r160 71 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r161 69 97 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.57 $Y=0 $X2=8.4
+ $Y2=0
r162 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.57 $Y=0 $X2=8.735
+ $Y2=0
r163 68 101 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=8.9 $Y=0 $X2=9.36
+ $Y2=0
r164 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.9 $Y=0 $X2=8.735
+ $Y2=0
r165 66 94 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.64 $Y=0 $X2=7.44
+ $Y2=0
r166 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.64 $Y=0 $X2=7.805
+ $Y2=0
r167 65 97 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.97 $Y=0 $X2=8.4
+ $Y2=0
r168 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.97 $Y=0 $X2=7.805
+ $Y2=0
r169 63 78 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.2
+ $Y2=0
r170 63 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.535
+ $Y2=0
r171 62 82 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.66 $Y=0 $X2=1.68
+ $Y2=0
r172 62 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.66 $Y=0 $X2=1.535
+ $Y2=0
r173 60 74 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r174 60 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.67
+ $Y2=0
r175 59 78 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.2
+ $Y2=0
r176 59 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.67
+ $Y2=0
r177 55 113 3.19436 $w=3.05e-07 $l=1.33918e-07 $layer=LI1_cond $X=9.732 $Y=0.085
+ $X2=9.83 $Y2=0
r178 55 57 21.1596 $w=3.03e-07 $l=5.6e-07 $layer=LI1_cond $X=9.732 $Y=0.085
+ $X2=9.732 $Y2=0.645
r179 51 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.735 $Y=0.085
+ $X2=8.735 $Y2=0
r180 51 53 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=8.735 $Y=0.085
+ $X2=8.735 $Y2=0.58
r181 47 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.805 $Y=0.085
+ $X2=7.805 $Y2=0
r182 47 49 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=7.805 $Y=0.085
+ $X2=7.805 $Y2=0.53
r183 43 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.945 $Y=0.085
+ $X2=6.945 $Y2=0
r184 43 45 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6.945 $Y=0.085
+ $X2=6.945 $Y2=0.53
r185 39 107 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.045 $Y=0.085
+ $X2=6.045 $Y2=0
r186 39 41 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.045 $Y=0.085
+ $X2=6.045 $Y2=0.515
r187 38 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.28 $Y=0
+ $X2=5.115 $Y2=0
r188 37 107 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.92 $Y=0
+ $X2=6.045 $Y2=0
r189 37 38 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.92 $Y=0 $X2=5.28
+ $Y2=0
r190 33 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.115 $Y=0.085
+ $X2=5.115 $Y2=0
r191 33 35 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=5.115 $Y=0.085
+ $X2=5.115 $Y2=0.74
r192 29 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=0.085
+ $X2=1.535 $Y2=0
r193 29 31 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=1.535 $Y=0.085
+ $X2=1.535 $Y2=0.775
r194 25 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r195 25 27 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.775
r196 8 57 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=9.58
+ $Y=0.37 $X2=9.72 $Y2=0.645
r197 7 53 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=8.525
+ $Y=0.37 $X2=8.735 $Y2=0.58
r198 6 49 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=7.665
+ $Y=0.37 $X2=7.805 $Y2=0.53
r199 5 45 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=6.805
+ $Y=0.37 $X2=6.945 $Y2=0.53
r200 4 41 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.95
+ $Y=0.37 $X2=6.085 $Y2=0.515
r201 3 35 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=4.905
+ $Y=0.595 $X2=5.115 $Y2=0.74
r202 2 31 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.625 $X2=1.575 $Y2=0.775
r203 1 27 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.625 $X2=0.71 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LS__HA_4%A_707_119# 1 2 3 12 14 15 19 20 21 24
c52 14 0 1.39181e-20 $X=4.45 $Y=0.4
r53 22 24 31.5769 $w=2.48e-07 $l=6.85e-07 $layer=LI1_cond $X=5.585 $Y=1.425
+ $X2=5.585 $Y2=0.74
r54 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.46 $Y=1.51
+ $X2=5.585 $Y2=1.425
r55 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.46 $Y=1.51
+ $X2=4.78 $Y2=1.51
r56 17 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.615 $Y=1.425
+ $X2=4.78 $Y2=1.51
r57 17 19 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=4.615 $Y=1.425
+ $X2=4.615 $Y2=0.74
r58 16 19 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.615 $Y=0.485
+ $X2=4.615 $Y2=0.74
r59 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.45 $Y=0.4
+ $X2=4.615 $Y2=0.485
r60 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.45 $Y=0.4 $X2=3.78
+ $Y2=0.4
r61 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.65 $Y=0.485
+ $X2=3.78 $Y2=0.4
r62 10 12 10.8596 $w=2.58e-07 $l=2.45e-07 $layer=LI1_cond $X=3.65 $Y=0.485
+ $X2=3.65 $Y2=0.73
r63 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.405
+ $Y=0.595 $X2=5.545 $Y2=0.74
r64 2 19 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=4.405
+ $Y=0.595 $X2=4.615 $Y2=0.74
r65 1 12 91 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=2 $X=3.535
+ $Y=0.595 $X2=3.685 $Y2=0.73
.ends

