# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__or4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__or4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.232500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 3.835000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.232500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.965000 1.350000 3.295000 2.890000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.455000 1.780000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.050000 1.315000 1.720000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.240000 1.820000 4.715000 2.980000 ;
        RECT 4.345000 0.350000 4.715000 1.130000 ;
        RECT 4.545000 1.130000 4.715000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  2.100000 0.795000 2.310000 ;
      RECT 0.115000  2.310000 1.285000 2.480000 ;
      RECT 0.115000  2.480000 0.445000 2.980000 ;
      RECT 0.140000  0.350000 0.470000 0.960000 ;
      RECT 0.140000  0.960000 0.795000 1.130000 ;
      RECT 0.615000  2.650000 0.945000 3.245000 ;
      RECT 0.625000  1.130000 0.795000 2.100000 ;
      RECT 0.640000  0.085000 0.970000 0.790000 ;
      RECT 1.115000  2.480000 1.285000 2.905000 ;
      RECT 1.115000  2.905000 2.755000 3.075000 ;
      RECT 1.140000  0.350000 1.655000 0.880000 ;
      RECT 1.150000  1.890000 1.655000 2.140000 ;
      RECT 1.485000  0.880000 1.655000 1.030000 ;
      RECT 1.485000  1.030000 1.905000 1.700000 ;
      RECT 1.485000  1.700000 1.655000 1.890000 ;
      RECT 1.825000  0.085000 2.075000 0.680000 ;
      RECT 1.845000  1.870000 2.245000 2.735000 ;
      RECT 2.075000  0.850000 3.640000 1.010000 ;
      RECT 2.075000  1.010000 4.175000 1.020000 ;
      RECT 2.075000  1.020000 2.245000 1.870000 ;
      RECT 2.245000  0.350000 2.575000 0.850000 ;
      RECT 2.425000  1.190000 2.755000 2.905000 ;
      RECT 2.745000  0.085000 3.140000 0.680000 ;
      RECT 3.310000  0.350000 3.640000 0.850000 ;
      RECT 3.310000  1.020000 4.175000 1.180000 ;
      RECT 3.740000  1.950000 4.070000 3.245000 ;
      RECT 3.810000  0.085000 4.140000 0.840000 ;
      RECT 4.005000  1.180000 4.175000 1.300000 ;
      RECT 4.005000  1.300000 4.375000 1.630000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_ls__or4bb_1
END LIBRARY
