* File: sky130_fd_sc_ls__o2111a_1.pxi.spice
* Created: Fri Aug 28 13:41:35 2020
* 
x_PM_SKY130_FD_SC_LS__O2111A_1%A_82_48# N_A_82_48#_M1009_s N_A_82_48#_M1003_d
+ N_A_82_48#_M1008_d N_A_82_48#_c_69_n N_A_82_48#_M1004_g N_A_82_48#_c_70_n
+ N_A_82_48#_M1006_g N_A_82_48#_c_71_n N_A_82_48#_c_72_n N_A_82_48#_c_82_p
+ N_A_82_48#_c_118_p N_A_82_48#_c_73_n N_A_82_48#_c_95_p N_A_82_48#_c_74_n
+ N_A_82_48#_c_77_n N_A_82_48#_c_78_n PM_SKY130_FD_SC_LS__O2111A_1%A_82_48#
x_PM_SKY130_FD_SC_LS__O2111A_1%D1 N_D1_c_143_n N_D1_M1003_g N_D1_c_144_n
+ N_D1_c_145_n N_D1_M1009_g N_D1_c_146_n D1 PM_SKY130_FD_SC_LS__O2111A_1%D1
x_PM_SKY130_FD_SC_LS__O2111A_1%C1 N_C1_c_183_n N_C1_M1007_g N_C1_M1010_g C1 C1
+ C1 C1 PM_SKY130_FD_SC_LS__O2111A_1%C1
x_PM_SKY130_FD_SC_LS__O2111A_1%B1 N_B1_M1011_g N_B1_c_224_n N_B1_c_225_n
+ N_B1_M1008_g B1 N_B1_c_222_n N_B1_c_223_n PM_SKY130_FD_SC_LS__O2111A_1%B1
x_PM_SKY130_FD_SC_LS__O2111A_1%A2 N_A2_M1002_g N_A2_c_258_n N_A2_M1001_g A2
+ PM_SKY130_FD_SC_LS__O2111A_1%A2
x_PM_SKY130_FD_SC_LS__O2111A_1%A1 N_A1_M1005_g N_A1_c_289_n N_A1_M1000_g A1
+ N_A1_c_290_n PM_SKY130_FD_SC_LS__O2111A_1%A1
x_PM_SKY130_FD_SC_LS__O2111A_1%X N_X_M1004_s N_X_M1006_s N_X_c_311_n N_X_c_312_n
+ X X X X N_X_c_313_n PM_SKY130_FD_SC_LS__O2111A_1%X
x_PM_SKY130_FD_SC_LS__O2111A_1%VPWR N_VPWR_M1006_d N_VPWR_M1007_d N_VPWR_M1000_d
+ N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_336_n N_VPWR_c_337_n VPWR
+ N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n
+ N_VPWR_c_333_n PM_SKY130_FD_SC_LS__O2111A_1%VPWR
x_PM_SKY130_FD_SC_LS__O2111A_1%VGND N_VGND_M1004_d N_VGND_M1002_d N_VGND_c_381_n
+ N_VGND_c_382_n VGND N_VGND_c_383_n N_VGND_c_384_n N_VGND_c_385_n
+ N_VGND_c_386_n N_VGND_c_387_n N_VGND_c_388_n PM_SKY130_FD_SC_LS__O2111A_1%VGND
x_PM_SKY130_FD_SC_LS__O2111A_1%A_471_74# N_A_471_74#_M1011_d N_A_471_74#_M1005_d
+ N_A_471_74#_c_425_n N_A_471_74#_c_426_n N_A_471_74#_c_427_n
+ N_A_471_74#_c_428_n PM_SKY130_FD_SC_LS__O2111A_1%A_471_74#
cc_1 VNB N_A_82_48#_c_69_n 0.0234345f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.22
cc_2 VNB N_A_82_48#_c_70_n 0.0442905f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_A_82_48#_c_71_n 0.00153124f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.07
cc_4 VNB N_A_82_48#_c_72_n 0.0174507f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.295
cc_5 VNB N_A_82_48#_c_73_n 0.0112873f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=0.515
cc_6 VNB N_A_82_48#_c_74_n 0.00538141f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.295
cc_7 VNB N_D1_c_143_n 0.0135911f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=0.37
cc_8 VNB N_D1_c_144_n 0.0135632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_D1_c_145_n 0.0165545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_D1_c_146_n 0.0324276f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_11 VNB D1 0.00165832f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_12 VNB N_C1_c_183_n 0.0136816f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=0.37
cc_13 VNB N_C1_M1010_g 0.0335784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB C1 0.0022543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_M1011_g 0.0291183f $X=-0.19 $Y=-0.245 $X2=2.465 $Y2=2.065
cc_16 VNB N_B1_c_222_n 0.0199249f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_17 VNB N_B1_c_223_n 0.00796532f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_18 VNB N_A2_M1002_g 0.0311844f $X=-0.19 $Y=-0.245 $X2=2.465 $Y2=2.065
cc_19 VNB N_A2_c_258_n 0.0185444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB A2 0.00520679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_M1005_g 0.0314484f $X=-0.19 $Y=-0.245 $X2=2.465 $Y2=2.065
cc_22 VNB N_A1_c_289_n 0.0604737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_c_290_n 0.00488709f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_24 VNB N_X_c_311_n 0.0235276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_312_n 0.00489291f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_26 VNB N_X_c_313_n 0.0284135f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.295
cc_27 VNB N_VPWR_c_333_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_381_n 0.0135318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_382_n 0.00975957f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_30 VNB N_VGND_c_383_n 0.0169946f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.07
cc_31 VNB N_VGND_c_384_n 0.0574108f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.21
cc_32 VNB N_VGND_c_385_n 0.0196288f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.295
cc_33 VNB N_VGND_c_386_n 0.249202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_387_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.385
cc_35 VNB N_VGND_c_388_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.24
cc_36 VNB N_A_471_74#_c_425_n 0.00335011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_471_74#_c_426_n 0.0131391f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_38 VNB N_A_471_74#_c_427_n 0.0095993f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_39 VNB N_A_471_74#_c_428_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_40 VPB N_A_82_48#_c_70_n 0.0285475f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_41 VPB N_A_82_48#_c_71_n 0.00314192f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.07
cc_42 VPB N_A_82_48#_c_77_n 0.00317243f $X=-0.19 $Y=1.66 $X2=1.36 $Y2=2.24
cc_43 VPB N_A_82_48#_c_78_n 0.00419846f $X=-0.19 $Y=1.66 $X2=2.7 $Y2=2.21
cc_44 VPB N_D1_c_143_n 0.0454261f $X=-0.19 $Y=1.66 $X2=1.105 $Y2=0.37
cc_45 VPB D1 0.00142441f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_46 VPB N_C1_c_183_n 0.0505577f $X=-0.19 $Y=1.66 $X2=1.105 $Y2=0.37
cc_47 VPB C1 0.00139918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_B1_c_224_n 0.0091881f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_B1_c_225_n 0.0247582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_B1_c_222_n 0.00899022f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_51 VPB N_B1_c_223_n 0.00470511f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_52 VPB N_A2_c_258_n 0.0303586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB A2 0.01111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A1_c_289_n 0.0314313f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A1_c_290_n 0.0072578f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=0.74
cc_56 VPB X 0.0130351f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_57 VPB X 0.0413071f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=0.515
cc_58 VPB N_X_c_313_n 0.0075834f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.295
cc_59 VPB N_VPWR_c_334_n 0.0112396f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=0.74
cc_60 VPB N_VPWR_c_335_n 0.0174875f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.55
cc_61 VPB N_VPWR_c_336_n 0.0118719f $X=-0.19 $Y=1.66 $X2=1.08 $Y2=1.295
cc_62 VPB N_VPWR_c_337_n 0.0513616f $X=-0.19 $Y=1.66 $X2=1.195 $Y2=2.155
cc_63 VPB N_VPWR_c_338_n 0.0189953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_339_n 0.0229347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_340_n 0.0331177f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.385
cc_66 VPB N_VPWR_c_341_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.587 $Y2=1.385
cc_67 VPB N_VPWR_c_342_n 0.0105532f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_333_n 0.0886544f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 N_A_82_48#_c_70_n N_D1_c_143_n 0.026643f $X=0.505 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_70 N_A_82_48#_c_71_n N_D1_c_143_n 0.00632537f $X=0.7 $Y=2.07 $X2=-0.19
+ $Y2=-0.245
cc_71 N_A_82_48#_c_72_n N_D1_c_143_n 0.0013382f $X=1.08 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_72 N_A_82_48#_c_82_p N_D1_c_143_n 0.0126958f $X=1.195 $Y=2.155 $X2=-0.19
+ $Y2=-0.245
cc_73 N_A_82_48#_c_77_n N_D1_c_143_n 0.0126005f $X=1.36 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_74 N_A_82_48#_c_72_n N_D1_c_144_n 0.00357242f $X=1.08 $Y=1.295 $X2=0 $Y2=0
cc_75 N_A_82_48#_c_74_n N_D1_c_144_n 0.00325742f $X=0.61 $Y=1.295 $X2=0 $Y2=0
cc_76 N_A_82_48#_c_73_n N_D1_c_145_n 0.0190115f $X=1.245 $Y=0.515 $X2=0 $Y2=0
cc_77 N_A_82_48#_c_69_n N_D1_c_146_n 4.52431e-19 $X=0.485 $Y=1.22 $X2=0 $Y2=0
cc_78 N_A_82_48#_c_70_n N_D1_c_146_n 0.00826486f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_79 N_A_82_48#_c_72_n N_D1_c_146_n 0.005455f $X=1.08 $Y=1.295 $X2=0 $Y2=0
cc_80 N_A_82_48#_c_73_n N_D1_c_146_n 0.00458903f $X=1.245 $Y=0.515 $X2=0 $Y2=0
cc_81 N_A_82_48#_c_71_n D1 0.0203563f $X=0.7 $Y=2.07 $X2=0 $Y2=0
cc_82 N_A_82_48#_c_72_n D1 0.0260844f $X=1.08 $Y=1.295 $X2=0 $Y2=0
cc_83 N_A_82_48#_c_82_p D1 0.0106923f $X=1.195 $Y=2.155 $X2=0 $Y2=0
cc_84 N_A_82_48#_c_77_n D1 0.00813566f $X=1.36 $Y=2.24 $X2=0 $Y2=0
cc_85 N_A_82_48#_c_95_p N_C1_c_183_n 0.0216559f $X=2.535 $Y=2.157 $X2=-0.19
+ $Y2=-0.245
cc_86 N_A_82_48#_c_77_n N_C1_c_183_n 0.00369784f $X=1.36 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_87 N_A_82_48#_c_72_n C1 0.0111966f $X=1.08 $Y=1.295 $X2=0 $Y2=0
cc_88 N_A_82_48#_c_73_n C1 0.0488331f $X=1.245 $Y=0.515 $X2=0 $Y2=0
cc_89 N_A_82_48#_c_95_p C1 0.0228671f $X=2.535 $Y=2.157 $X2=0 $Y2=0
cc_90 N_A_82_48#_c_95_p N_B1_c_225_n 0.0177773f $X=2.535 $Y=2.157 $X2=0 $Y2=0
cc_91 N_A_82_48#_c_78_n N_B1_c_225_n 0.0111095f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_92 N_A_82_48#_c_95_p N_B1_c_222_n 6.16889e-19 $X=2.535 $Y=2.157 $X2=0 $Y2=0
cc_93 N_A_82_48#_c_95_p N_B1_c_223_n 0.0212242f $X=2.535 $Y=2.157 $X2=0 $Y2=0
cc_94 N_A_82_48#_c_78_n N_A2_c_258_n 0.0182576f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_95 N_A_82_48#_c_78_n A2 0.00747271f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_96 N_A_82_48#_c_78_n N_A1_c_289_n 0.0025366f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_97 N_A_82_48#_c_69_n N_X_c_311_n 4.44442e-19 $X=0.485 $Y=1.22 $X2=0 $Y2=0
cc_98 N_A_82_48#_c_70_n X 0.00358528f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_82_48#_c_71_n X 0.0101424f $X=0.7 $Y=2.07 $X2=0 $Y2=0
cc_100 N_A_82_48#_c_74_n X 4.42944e-19 $X=0.61 $Y=1.295 $X2=0 $Y2=0
cc_101 N_A_82_48#_c_70_n X 0.0129519f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_82_48#_c_69_n N_X_c_313_n 0.013355f $X=0.485 $Y=1.22 $X2=0 $Y2=0
cc_103 N_A_82_48#_c_70_n N_X_c_313_n 0.00595318f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_104 N_A_82_48#_c_71_n N_X_c_313_n 0.012249f $X=0.7 $Y=2.07 $X2=0 $Y2=0
cc_105 N_A_82_48#_c_74_n N_X_c_313_n 0.02563f $X=0.61 $Y=1.295 $X2=0 $Y2=0
cc_106 N_A_82_48#_c_71_n N_VPWR_M1006_d 0.00455057f $X=0.7 $Y=2.07 $X2=-0.19
+ $Y2=-0.245
cc_107 N_A_82_48#_c_82_p N_VPWR_M1006_d 0.0130846f $X=1.195 $Y=2.155 $X2=-0.19
+ $Y2=-0.245
cc_108 N_A_82_48#_c_118_p N_VPWR_M1006_d 0.00301935f $X=0.785 $Y=2.155 $X2=-0.19
+ $Y2=-0.245
cc_109 N_A_82_48#_c_95_p N_VPWR_M1007_d 0.0156961f $X=2.535 $Y=2.157 $X2=0 $Y2=0
cc_110 N_A_82_48#_c_70_n N_VPWR_c_334_n 0.00799654f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_111 N_A_82_48#_c_82_p N_VPWR_c_334_n 0.0128995f $X=1.195 $Y=2.155 $X2=0 $Y2=0
cc_112 N_A_82_48#_c_118_p N_VPWR_c_334_n 0.0132989f $X=0.785 $Y=2.155 $X2=0
+ $Y2=0
cc_113 N_A_82_48#_c_77_n N_VPWR_c_334_n 0.0297396f $X=1.36 $Y=2.24 $X2=0 $Y2=0
cc_114 N_A_82_48#_c_95_p N_VPWR_c_335_n 0.034201f $X=2.535 $Y=2.157 $X2=0 $Y2=0
cc_115 N_A_82_48#_c_77_n N_VPWR_c_335_n 0.00139437f $X=1.36 $Y=2.24 $X2=0 $Y2=0
cc_116 N_A_82_48#_c_78_n N_VPWR_c_335_n 0.0150858f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_117 N_A_82_48#_c_78_n N_VPWR_c_337_n 0.0258853f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_118 N_A_82_48#_c_70_n N_VPWR_c_338_n 0.00445602f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_119 N_A_82_48#_c_77_n N_VPWR_c_339_n 0.0119397f $X=1.36 $Y=2.24 $X2=0 $Y2=0
cc_120 N_A_82_48#_c_78_n N_VPWR_c_340_n 0.0119397f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_121 N_A_82_48#_c_70_n N_VPWR_c_333_n 0.00865213f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_122 N_A_82_48#_c_77_n N_VPWR_c_333_n 0.0116912f $X=1.36 $Y=2.24 $X2=0 $Y2=0
cc_123 N_A_82_48#_c_78_n N_VPWR_c_333_n 0.0116912f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_124 N_A_82_48#_c_69_n N_VGND_c_381_n 0.0156276f $X=0.485 $Y=1.22 $X2=0 $Y2=0
cc_125 N_A_82_48#_c_70_n N_VGND_c_381_n 0.00140504f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_126 N_A_82_48#_c_72_n N_VGND_c_381_n 0.00658384f $X=1.08 $Y=1.295 $X2=0 $Y2=0
cc_127 N_A_82_48#_c_73_n N_VGND_c_381_n 0.0477412f $X=1.245 $Y=0.515 $X2=0 $Y2=0
cc_128 N_A_82_48#_c_74_n N_VGND_c_381_n 0.019655f $X=0.61 $Y=1.295 $X2=0 $Y2=0
cc_129 N_A_82_48#_c_69_n N_VGND_c_383_n 0.00383152f $X=0.485 $Y=1.22 $X2=0 $Y2=0
cc_130 N_A_82_48#_c_73_n N_VGND_c_384_n 0.011066f $X=1.245 $Y=0.515 $X2=0 $Y2=0
cc_131 N_A_82_48#_c_69_n N_VGND_c_386_n 0.00761163f $X=0.485 $Y=1.22 $X2=0 $Y2=0
cc_132 N_A_82_48#_c_73_n N_VGND_c_386_n 0.00915947f $X=1.245 $Y=0.515 $X2=0
+ $Y2=0
cc_133 N_D1_c_143_n N_C1_c_183_n 0.0450198f $X=1.135 $Y=1.99 $X2=-0.19
+ $Y2=-0.245
cc_134 N_D1_c_146_n N_C1_c_183_n 0.00342787f $X=1.53 $Y=1.26 $X2=-0.19
+ $Y2=-0.245
cc_135 D1 N_C1_c_183_n 0.00112962f $X=1.115 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_136 N_D1_c_144_n N_C1_M1010_g 0.0043485f $X=1.26 $Y=1.55 $X2=0 $Y2=0
cc_137 N_D1_c_145_n N_C1_M1010_g 0.0705403f $X=1.53 $Y=1.185 $X2=0 $Y2=0
cc_138 N_D1_c_143_n C1 0.00120371f $X=1.135 $Y=1.99 $X2=0 $Y2=0
cc_139 N_D1_c_144_n C1 0.00464587f $X=1.26 $Y=1.55 $X2=0 $Y2=0
cc_140 N_D1_c_145_n C1 0.0181159f $X=1.53 $Y=1.185 $X2=0 $Y2=0
cc_141 N_D1_c_146_n C1 0.00518893f $X=1.53 $Y=1.26 $X2=0 $Y2=0
cc_142 D1 C1 0.0209972f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_143 N_D1_c_143_n X 9.40448e-19 $X=1.135 $Y=1.99 $X2=0 $Y2=0
cc_144 N_D1_c_143_n N_VPWR_c_334_n 0.00813312f $X=1.135 $Y=1.99 $X2=0 $Y2=0
cc_145 N_D1_c_143_n N_VPWR_c_339_n 0.00523995f $X=1.135 $Y=1.99 $X2=0 $Y2=0
cc_146 N_D1_c_143_n N_VPWR_c_333_n 0.00528353f $X=1.135 $Y=1.99 $X2=0 $Y2=0
cc_147 N_D1_c_145_n N_VGND_c_381_n 0.00361162f $X=1.53 $Y=1.185 $X2=0 $Y2=0
cc_148 N_D1_c_145_n N_VGND_c_384_n 0.0039925f $X=1.53 $Y=1.185 $X2=0 $Y2=0
cc_149 N_D1_c_145_n N_VGND_c_386_n 0.00702246f $X=1.53 $Y=1.185 $X2=0 $Y2=0
cc_150 N_C1_M1010_g N_B1_M1011_g 0.0599213f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_151 C1 N_B1_M1011_g 0.00363173f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_152 N_C1_c_183_n N_B1_c_224_n 0.00615951f $X=1.635 $Y=1.99 $X2=0 $Y2=0
cc_153 C1 N_B1_c_224_n 6.48925e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_154 N_C1_c_183_n N_B1_c_225_n 0.0180292f $X=1.635 $Y=1.99 $X2=0 $Y2=0
cc_155 N_C1_M1010_g N_B1_c_222_n 0.0200714f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_156 C1 N_B1_c_222_n 2.77362e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_157 N_C1_M1010_g N_B1_c_223_n 0.0025595f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_158 C1 N_B1_c_223_n 0.0296056f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_159 N_C1_c_183_n N_VPWR_c_335_n 0.00784051f $X=1.635 $Y=1.99 $X2=0 $Y2=0
cc_160 N_C1_c_183_n N_VPWR_c_339_n 0.00537957f $X=1.635 $Y=1.99 $X2=0 $Y2=0
cc_161 N_C1_c_183_n N_VPWR_c_333_n 0.00528353f $X=1.635 $Y=1.99 $X2=0 $Y2=0
cc_162 N_C1_M1010_g N_VGND_c_384_n 0.0039925f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_163 C1 N_VGND_c_384_n 0.00851294f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_164 N_C1_M1010_g N_VGND_c_386_n 0.00696958f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_165 C1 N_VGND_c_386_n 0.0108483f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_166 C1 A_321_74# 0.00133334f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_167 C1 N_A_471_74#_c_427_n 0.0030385f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_168 N_B1_M1011_g N_A2_M1002_g 0.0179083f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_169 N_B1_c_224_n N_A2_c_258_n 0.00961814f $X=2.39 $Y=1.9 $X2=0 $Y2=0
cc_170 N_B1_c_225_n N_A2_c_258_n 0.0180664f $X=2.39 $Y=1.99 $X2=0 $Y2=0
cc_171 N_B1_c_222_n N_A2_c_258_n 0.0214219f $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_172 N_B1_c_223_n N_A2_c_258_n 5.21437e-19 $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_173 N_B1_c_222_n A2 4.13845e-19 $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_174 N_B1_c_223_n A2 0.0249368f $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_175 N_B1_c_225_n N_VPWR_c_335_n 0.00791639f $X=2.39 $Y=1.99 $X2=0 $Y2=0
cc_176 N_B1_c_225_n N_VPWR_c_340_n 0.00537957f $X=2.39 $Y=1.99 $X2=0 $Y2=0
cc_177 N_B1_c_225_n N_VPWR_c_333_n 0.00528353f $X=2.39 $Y=1.99 $X2=0 $Y2=0
cc_178 N_B1_M1011_g N_VGND_c_384_n 0.00461464f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_179 N_B1_M1011_g N_VGND_c_386_n 0.00909821f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B1_M1011_g N_A_471_74#_c_425_n 8.94767e-19 $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_181 N_B1_M1011_g N_A_471_74#_c_427_n 3.11521e-19 $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B1_c_222_n N_A_471_74#_c_427_n 0.00306064f $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_183 N_B1_c_223_n N_A_471_74#_c_427_n 0.00722443f $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_184 N_A2_M1002_g N_A1_M1005_g 0.0277451f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A2_c_258_n N_A1_c_289_n 0.078453f $X=2.925 $Y=1.83 $X2=0 $Y2=0
cc_186 A2 N_A1_c_289_n 0.00294298f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_187 N_A2_M1002_g N_A1_c_290_n 5.08722e-19 $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A2_c_258_n N_A1_c_290_n 2.55968e-19 $X=2.925 $Y=1.83 $X2=0 $Y2=0
cc_189 A2 N_A1_c_290_n 0.0299389f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_190 N_A2_c_258_n N_VPWR_c_337_n 0.00352411f $X=2.925 $Y=1.83 $X2=0 $Y2=0
cc_191 N_A2_c_258_n N_VPWR_c_340_n 0.00523995f $X=2.925 $Y=1.83 $X2=0 $Y2=0
cc_192 N_A2_c_258_n N_VPWR_c_333_n 0.00528353f $X=2.925 $Y=1.83 $X2=0 $Y2=0
cc_193 N_A2_M1002_g N_VGND_c_382_n 0.0036453f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A2_M1002_g N_VGND_c_384_n 0.00461464f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A2_M1002_g N_VGND_c_386_n 0.00909258f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A2_M1002_g N_A_471_74#_c_425_n 5.32432e-19 $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A2_M1002_g N_A_471_74#_c_426_n 0.0144173f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A2_c_258_n N_A_471_74#_c_426_n 0.00421088f $X=2.925 $Y=1.83 $X2=0 $Y2=0
cc_199 A2 N_A_471_74#_c_426_n 0.0270243f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_200 N_A2_M1002_g N_A_471_74#_c_428_n 6.2684e-19 $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A1_c_289_n N_VPWR_c_337_n 0.0230907f $X=3.345 $Y=1.83 $X2=0 $Y2=0
cc_202 N_A1_c_290_n N_VPWR_c_337_n 0.0266442f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_203 N_A1_c_289_n N_VPWR_c_340_n 0.0048289f $X=3.345 $Y=1.83 $X2=0 $Y2=0
cc_204 N_A1_c_289_n N_VPWR_c_333_n 0.0047904f $X=3.345 $Y=1.83 $X2=0 $Y2=0
cc_205 N_A1_M1005_g N_VGND_c_382_n 0.00572341f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A1_M1005_g N_VGND_c_385_n 0.00434272f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A1_M1005_g N_VGND_c_386_n 0.00824797f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A1_M1005_g N_A_471_74#_c_426_n 0.017525f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A1_c_289_n N_A_471_74#_c_426_n 0.00240389f $X=3.345 $Y=1.83 $X2=0 $Y2=0
cc_210 N_A1_c_290_n N_A_471_74#_c_426_n 0.0264387f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_211 N_A1_M1005_g N_A_471_74#_c_428_n 0.00977408f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_212 X N_VPWR_c_334_n 0.0223718f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_213 X N_VPWR_c_338_n 0.0154862f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_214 X N_VPWR_c_333_n 0.0127853f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_215 N_X_c_311_n N_VGND_c_381_n 0.0254628f $X=0.27 $Y=0.515 $X2=0 $Y2=0
cc_216 N_X_c_311_n N_VGND_c_383_n 0.0115164f $X=0.27 $Y=0.515 $X2=0 $Y2=0
cc_217 N_X_c_311_n N_VGND_c_386_n 0.00953044f $X=0.27 $Y=0.515 $X2=0 $Y2=0
cc_218 N_VGND_c_382_n N_A_471_74#_c_425_n 0.00158095f $X=3.045 $Y=0.57 $X2=0
+ $Y2=0
cc_219 N_VGND_c_384_n N_A_471_74#_c_425_n 0.0146357f $X=2.88 $Y=0 $X2=0 $Y2=0
cc_220 N_VGND_c_386_n N_A_471_74#_c_425_n 0.0121141f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_221 N_VGND_M1002_d N_A_471_74#_c_426_n 0.00318135f $X=2.865 $Y=0.37 $X2=0
+ $Y2=0
cc_222 N_VGND_c_382_n N_A_471_74#_c_426_n 0.022455f $X=3.045 $Y=0.57 $X2=0 $Y2=0
cc_223 N_VGND_c_382_n N_A_471_74#_c_428_n 0.0173003f $X=3.045 $Y=0.57 $X2=0
+ $Y2=0
cc_224 N_VGND_c_385_n N_A_471_74#_c_428_n 0.0145639f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_225 N_VGND_c_386_n N_A_471_74#_c_428_n 0.0119984f $X=3.6 $Y=0 $X2=0 $Y2=0
