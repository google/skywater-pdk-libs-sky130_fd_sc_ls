* NGSPICE file created from sky130_fd_sc_ls__or4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
M1000 a_182_270# B VGND VNB nshort w=640000u l=150000u
+  ad=5.192e+11p pd=4.27e+06u as=1.16472e+12p ps=9.37e+06u
M1001 a_548_110# C_N VPWR VPB phighvt w=840000u l=150000u
+  ad=2.436e+11p pd=2.26e+06u as=1.0664e+12p ps=8.54e+06u
M1002 X a_182_270# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1003 VGND a_182_270# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND D_N a_27_424# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1005 a_587_392# a_548_110# a_503_392# VPB phighvt w=1e+06u l=150000u
+  ad=3.6e+11p pd=2.72e+06u as=2.7e+11p ps=2.54e+06u
M1006 a_689_392# B a_587_392# VPB phighvt w=1e+06u l=150000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1007 a_548_110# C_N VGND VNB nshort w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1008 X a_182_270# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1009 a_503_392# a_27_424# a_182_270# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1010 VPWR D_N a_27_424# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.25e+06u
M1011 a_182_270# a_27_424# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A a_182_270# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_182_270# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_548_110# a_182_270# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A a_689_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

