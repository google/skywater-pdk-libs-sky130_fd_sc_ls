* NGSPICE file created from sky130_fd_sc_ls__and3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__and3b_4 A_N B C VGND VNB VPB VPWR X
M1000 a_239_98# a_27_74# a_298_368# VNB nshort w=640000u l=150000u
+  ad=5.44e+11p pd=5.54e+06u as=1.792e+11p ps=1.84e+06u
M1001 a_298_368# B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=9e+11p pd=7.8e+06u as=2.5708e+12p ps=1.76e+07u
M1002 a_498_98# C VGND VNB nshort w=640000u l=150000u
+  ad=4.032e+11p pd=3.82e+06u as=1.063e+12p ps=1.005e+07u
M1003 VGND a_298_368# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.662e+11p ps=4.22e+06u
M1004 a_298_368# C VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_298_368# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.72e+11p ps=5.68e+06u
M1006 X a_298_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_298_368# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B a_298_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR C a_298_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_298_368# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_298_368# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND C a_498_98# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A_N a_27_74# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1014 a_239_98# B a_498_98# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_498_98# B a_239_98# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_298_368# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_298_368# a_27_74# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_298_368# a_27_74# a_239_98# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A_N a_27_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1020 VPWR a_27_74# a_298_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_298_368# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

