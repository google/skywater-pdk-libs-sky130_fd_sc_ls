* File: sky130_fd_sc_ls__a222o_2.pxi.spice
* Created: Fri Aug 28 12:54:12 2020
* 
x_PM_SKY130_FD_SC_LS__A222O_2%C1 N_C1_M1001_g N_C1_M1013_g N_C1_c_91_n
+ N_C1_c_95_n C1 N_C1_c_92_n N_C1_c_93_n PM_SKY130_FD_SC_LS__A222O_2%C1
x_PM_SKY130_FD_SC_LS__A222O_2%C2 N_C2_M1011_g N_C2_c_124_n N_C2_c_128_n
+ N_C2_M1012_g C2 N_C2_c_125_n N_C2_c_126_n PM_SKY130_FD_SC_LS__A222O_2%C2
x_PM_SKY130_FD_SC_LS__A222O_2%A_27_82# N_A_27_82#_M1001_s N_A_27_82#_M1003_d
+ N_A_27_82#_M1013_s N_A_27_82#_M1012_d N_A_27_82#_c_161_n N_A_27_82#_M1002_g
+ N_A_27_82#_c_162_n N_A_27_82#_c_163_n N_A_27_82#_c_175_n N_A_27_82#_M1000_g
+ N_A_27_82#_c_164_n N_A_27_82#_M1006_g N_A_27_82#_c_176_n N_A_27_82#_M1004_g
+ N_A_27_82#_c_165_n N_A_27_82#_c_177_n N_A_27_82#_c_178_n N_A_27_82#_c_166_n
+ N_A_27_82#_c_167_n N_A_27_82#_c_179_n N_A_27_82#_c_202_n N_A_27_82#_c_168_n
+ N_A_27_82#_c_169_n N_A_27_82#_c_263_p N_A_27_82#_c_248_p N_A_27_82#_c_170_n
+ N_A_27_82#_c_171_n N_A_27_82#_c_172_n N_A_27_82#_c_264_p N_A_27_82#_c_173_n
+ N_A_27_82#_c_174_n PM_SKY130_FD_SC_LS__A222O_2%A_27_82#
x_PM_SKY130_FD_SC_LS__A222O_2%A1 N_A1_c_293_n N_A1_M1008_g N_A1_M1003_g A1 A1
+ N_A1_c_295_n PM_SKY130_FD_SC_LS__A222O_2%A1
x_PM_SKY130_FD_SC_LS__A222O_2%B1 N_B1_c_332_n N_B1_M1005_g N_B1_M1009_g B1
+ N_B1_c_334_n PM_SKY130_FD_SC_LS__A222O_2%B1
x_PM_SKY130_FD_SC_LS__A222O_2%B2 N_B2_M1007_g N_B2_c_362_n N_B2_M1010_g B2
+ N_B2_c_363_n PM_SKY130_FD_SC_LS__A222O_2%B2
x_PM_SKY130_FD_SC_LS__A222O_2%A2 N_A2_M1015_g N_A2_c_395_n N_A2_M1014_g A2
+ PM_SKY130_FD_SC_LS__A222O_2%A2
x_PM_SKY130_FD_SC_LS__A222O_2%A_116_392# N_A_116_392#_M1013_d
+ N_A_116_392#_M1005_d N_A_116_392#_c_417_n N_A_116_392#_c_431_n
+ N_A_116_392#_c_418_n PM_SKY130_FD_SC_LS__A222O_2%A_116_392#
x_PM_SKY130_FD_SC_LS__A222O_2%VPWR N_VPWR_M1000_s N_VPWR_M1004_s N_VPWR_M1014_d
+ N_VPWR_c_452_n N_VPWR_c_453_n N_VPWR_c_454_n N_VPWR_c_455_n N_VPWR_c_456_n
+ N_VPWR_c_457_n VPWR N_VPWR_c_458_n N_VPWR_c_459_n N_VPWR_c_460_n
+ N_VPWR_c_451_n PM_SKY130_FD_SC_LS__A222O_2%VPWR
x_PM_SKY130_FD_SC_LS__A222O_2%X N_X_M1002_d N_X_M1000_d N_X_c_501_n X
+ N_X_c_503_n PM_SKY130_FD_SC_LS__A222O_2%X
x_PM_SKY130_FD_SC_LS__A222O_2%A_639_368# N_A_639_368#_M1008_d
+ N_A_639_368#_M1010_d N_A_639_368#_c_530_n N_A_639_368#_c_531_n
+ N_A_639_368#_c_532_n PM_SKY130_FD_SC_LS__A222O_2%A_639_368#
x_PM_SKY130_FD_SC_LS__A222O_2%VGND N_VGND_M1011_d N_VGND_M1006_s N_VGND_M1007_d
+ N_VGND_c_553_n N_VGND_c_554_n N_VGND_c_555_n N_VGND_c_556_n N_VGND_c_557_n
+ N_VGND_c_558_n N_VGND_c_559_n N_VGND_c_560_n VGND N_VGND_c_561_n
+ N_VGND_c_562_n PM_SKY130_FD_SC_LS__A222O_2%VGND
x_PM_SKY130_FD_SC_LS__A222O_2%A_557_74# N_A_557_74#_M1003_s N_A_557_74#_M1015_d
+ N_A_557_74#_c_616_n N_A_557_74#_c_653_p N_A_557_74#_c_617_n
+ N_A_557_74#_c_618_n N_A_557_74#_c_619_n N_A_557_74#_c_620_n
+ PM_SKY130_FD_SC_LS__A222O_2%A_557_74#
cc_1 VNB N_C1_M1001_g 0.0329894f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_2 VNB N_C1_c_91_n 0.00186909f $X=-0.19 $Y=-0.245 $X2=0.497 $Y2=1.83
cc_3 VNB N_C1_c_92_n 0.00453376f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_C1_c_93_n 0.057529f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_5 VNB N_C2_M1011_g 0.0237179f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_6 VNB N_C2_c_124_n 0.00425652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_C2_c_125_n 0.0320644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_C2_c_126_n 0.00834647f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_9 VNB N_A_27_82#_c_161_n 0.0182542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_82#_c_162_n 0.013455f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_11 VNB N_A_27_82#_c_163_n 0.013716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_82#_c_164_n 0.0165924f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_13 VNB N_A_27_82#_c_165_n 0.0220451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_82#_c_166_n 0.0109097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_82#_c_167_n 0.00886217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_82#_c_168_n 0.0102068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_82#_c_169_n 0.0021754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_82#_c_170_n 0.00351331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_82#_c_171_n 0.0629583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_82#_c_172_n 0.0255526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_82#_c_173_n 0.00378718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_82#_c_174_n 0.0103491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_c_293_n 0.0280525f $X=-0.19 $Y=-0.245 $X2=0.492 $Y2=1.63
cc_24 VNB N_A1_M1003_g 0.0367638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_c_295_n 0.0016809f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_26 VNB N_B1_c_332_n 0.0315869f $X=-0.19 $Y=-0.245 $X2=0.492 $Y2=1.63
cc_27 VNB N_B1_M1009_g 0.0313709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B1_c_334_n 0.00240839f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_29 VNB N_B2_M1007_g 0.0290869f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_30 VNB N_B2_c_362_n 0.0224538f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_31 VNB N_B2_c_363_n 0.0054107f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_32 VNB N_A2_M1015_g 0.0411723f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_33 VNB N_A2_c_395_n 0.0276611f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_34 VNB A2 0.0159538f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_35 VNB N_VPWR_c_451_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_501_n 0.00209829f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_37 VNB N_VGND_c_553_n 0.00881119f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_38 VNB N_VGND_c_554_n 0.00671846f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_39 VNB N_VGND_c_555_n 0.0301057f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_40 VNB N_VGND_c_556_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_557_n 0.0168493f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_42 VNB N_VGND_c_558_n 0.0282128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_559_n 0.0443678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_560_n 0.00617641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_561_n 0.0215382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_562_n 0.330142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_557_74#_c_616_n 0.00610588f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_48 VNB N_A_557_74#_c_617_n 0.0269419f $X=-0.19 $Y=-0.245 $X2=0.497 $Y2=1.885
cc_49 VNB N_A_557_74#_c_618_n 0.00403445f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_50 VNB N_A_557_74#_c_619_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_51 VNB N_A_557_74#_c_620_n 0.00917671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VPB N_C1_c_91_n 0.0118236f $X=-0.19 $Y=1.66 $X2=0.497 $Y2=1.83
cc_53 VPB N_C1_c_95_n 0.0265759f $X=-0.19 $Y=1.66 $X2=0.497 $Y2=1.885
cc_54 VPB N_C1_c_92_n 0.00761937f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_55 VPB N_C2_c_124_n 0.00829991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_C2_c_128_n 0.0242543f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_57 VPB N_C2_c_126_n 0.00530202f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_58 VPB N_A_27_82#_c_175_n 0.0168457f $X=-0.19 $Y=1.66 $X2=0.492 $Y2=1.465
cc_59 VPB N_A_27_82#_c_176_n 0.0166737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_27_82#_c_177_n 0.0120621f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_27_82#_c_178_n 0.0310277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_27_82#_c_179_n 0.0175842f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_27_82#_c_168_n 0.00646682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_27_82#_c_171_n 0.0147183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A1_c_293_n 0.028304f $X=-0.19 $Y=1.66 $X2=0.492 $Y2=1.63
cc_66 VPB N_A1_c_295_n 0.00342331f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_67 VPB N_B1_c_332_n 0.0298433f $X=-0.19 $Y=1.66 $X2=0.492 $Y2=1.63
cc_68 VPB N_B1_c_334_n 0.00443927f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_69 VPB N_B2_c_362_n 0.0258518f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.73
cc_70 VPB N_B2_c_363_n 0.00567312f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_71 VPB N_A2_c_395_n 0.0311017f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.73
cc_72 VPB A2 0.00894665f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_73 VPB N_A_116_392#_c_417_n 0.015467f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_74 VPB N_A_116_392#_c_418_n 0.00256835f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_75 VPB N_VPWR_c_452_n 0.0150746f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_76 VPB N_VPWR_c_453_n 0.010686f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_77 VPB N_VPWR_c_454_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0.492 $Y2=1.465
cc_78 VPB N_VPWR_c_455_n 0.0515024f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_456_n 0.0234846f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_80 VPB N_VPWR_c_457_n 0.00632279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_458_n 0.0477633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_459_n 0.0459735f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_460_n 0.00632279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_451_n 0.0843705f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_X_c_501_n 0.00253211f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_86 VPB N_X_c_503_n 0.00644552f $X=-0.19 $Y=1.66 $X2=0.492 $Y2=1.465
cc_87 VPB N_A_639_368#_c_530_n 0.0151211f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_88 VPB N_A_639_368#_c_531_n 0.00140203f $X=-0.19 $Y=1.66 $X2=0.497 $Y2=1.885
cc_89 VPB N_A_639_368#_c_532_n 0.00624697f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_90 N_C1_M1001_g N_C2_M1011_g 0.0346947f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_91 N_C1_c_93_n N_C2_c_124_n 0.00480053f $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_92 N_C1_c_91_n N_C2_c_128_n 0.00480053f $X=0.497 $Y=1.83 $X2=0 $Y2=0
cc_93 N_C1_c_95_n N_C2_c_128_n 0.0248473f $X=0.497 $Y=1.885 $X2=0 $Y2=0
cc_94 N_C1_c_92_n N_C2_c_125_n 2.1027e-19 $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_95 N_C1_c_93_n N_C2_c_125_n 0.0346947f $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_96 N_C1_M1001_g N_C2_c_126_n 0.00533482f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_97 N_C1_c_92_n N_C2_c_126_n 0.0395606f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_98 N_C1_M1001_g N_A_27_82#_c_165_n 5.45389e-19 $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_99 N_C1_c_92_n N_A_27_82#_c_177_n 0.0228254f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_100 N_C1_c_93_n N_A_27_82#_c_177_n 0.00137994f $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_101 N_C1_c_95_n N_A_27_82#_c_178_n 0.00607013f $X=0.497 $Y=1.885 $X2=0 $Y2=0
cc_102 N_C1_M1001_g N_A_27_82#_c_166_n 0.0174317f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_103 N_C1_c_92_n N_A_27_82#_c_166_n 0.00448606f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_104 N_C1_c_93_n N_A_27_82#_c_166_n 3.67898e-19 $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_105 N_C1_c_92_n N_A_27_82#_c_167_n 0.0185799f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_106 N_C1_c_93_n N_A_27_82#_c_167_n 0.00192177f $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_107 N_C1_c_95_n N_A_27_82#_c_179_n 0.0202448f $X=0.497 $Y=1.885 $X2=0 $Y2=0
cc_108 N_C1_c_92_n N_A_27_82#_c_179_n 0.00568215f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_109 N_C1_c_93_n N_A_27_82#_c_179_n 2.49658e-19 $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_110 N_C1_c_95_n N_A_116_392#_c_418_n 0.007054f $X=0.497 $Y=1.885 $X2=0 $Y2=0
cc_111 N_C1_c_95_n N_VPWR_c_458_n 0.00445602f $X=0.497 $Y=1.885 $X2=0 $Y2=0
cc_112 N_C1_c_95_n N_VPWR_c_451_n 0.00861929f $X=0.497 $Y=1.885 $X2=0 $Y2=0
cc_113 N_C1_M1001_g N_VGND_c_553_n 0.00160827f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_114 N_C1_M1001_g N_VGND_c_555_n 0.00548708f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_115 N_C1_M1001_g N_VGND_c_562_n 0.00533081f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_116 N_C2_M1011_g N_A_27_82#_c_161_n 0.009666f $X=0.885 $Y=0.73 $X2=0 $Y2=0
cc_117 N_C2_c_125_n N_A_27_82#_c_163_n 0.00361438f $X=0.975 $Y=1.425 $X2=0 $Y2=0
cc_118 N_C2_M1011_g N_A_27_82#_c_166_n 0.0150237f $X=0.885 $Y=0.73 $X2=0 $Y2=0
cc_119 N_C2_c_125_n N_A_27_82#_c_166_n 0.00435908f $X=0.975 $Y=1.425 $X2=0 $Y2=0
cc_120 N_C2_c_126_n N_A_27_82#_c_166_n 0.0419923f $X=0.975 $Y=1.425 $X2=0 $Y2=0
cc_121 N_C2_c_128_n N_A_27_82#_c_179_n 0.0117748f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_122 N_C2_c_125_n N_A_27_82#_c_179_n 6.93298e-19 $X=0.975 $Y=1.425 $X2=0 $Y2=0
cc_123 N_C2_c_126_n N_A_27_82#_c_179_n 0.0438342f $X=0.975 $Y=1.425 $X2=0 $Y2=0
cc_124 N_C2_M1011_g N_A_27_82#_c_202_n 0.00296638f $X=0.885 $Y=0.73 $X2=0 $Y2=0
cc_125 N_C2_M1011_g N_A_27_82#_c_168_n 0.00304065f $X=0.885 $Y=0.73 $X2=0 $Y2=0
cc_126 N_C2_c_124_n N_A_27_82#_c_168_n 0.00420027f $X=0.955 $Y=1.795 $X2=0 $Y2=0
cc_127 N_C2_c_128_n N_A_27_82#_c_168_n 0.00185743f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_128 N_C2_c_125_n N_A_27_82#_c_168_n 0.001751f $X=0.975 $Y=1.425 $X2=0 $Y2=0
cc_129 N_C2_c_126_n N_A_27_82#_c_168_n 0.0348642f $X=0.975 $Y=1.425 $X2=0 $Y2=0
cc_130 N_C2_c_128_n N_A_116_392#_c_417_n 0.0109425f $X=0.955 $Y=1.885 $X2=0
+ $Y2=0
cc_131 N_C2_c_128_n N_A_116_392#_c_418_n 0.019456f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_132 N_C2_c_128_n N_VPWR_c_452_n 0.00947784f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_133 N_C2_c_128_n N_VPWR_c_458_n 0.00445602f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_134 N_C2_c_128_n N_VPWR_c_451_n 0.00447124f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_135 N_C2_c_128_n N_X_c_503_n 4.19771e-19 $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_136 N_C2_M1011_g N_VGND_c_553_n 0.0110632f $X=0.885 $Y=0.73 $X2=0 $Y2=0
cc_137 N_C2_M1011_g N_VGND_c_555_n 0.00455951f $X=0.885 $Y=0.73 $X2=0 $Y2=0
cc_138 N_C2_M1011_g N_VGND_c_562_n 0.00447788f $X=0.885 $Y=0.73 $X2=0 $Y2=0
cc_139 N_A_27_82#_c_176_n N_A1_c_293_n 0.0276252f $X=2.5 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_140 N_A_27_82#_c_170_n N_A1_c_293_n 9.97553e-19 $X=2.395 $Y=1.425 $X2=-0.19
+ $Y2=-0.245
cc_141 N_A_27_82#_c_171_n N_A1_c_293_n 0.0133229f $X=2.395 $Y=1.425 $X2=-0.19
+ $Y2=-0.245
cc_142 N_A_27_82#_c_172_n N_A1_c_293_n 0.00125579f $X=3.265 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A_27_82#_c_170_n N_A1_M1003_g 0.00245637f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_144 N_A_27_82#_c_171_n N_A1_M1003_g 0.00233427f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_145 N_A_27_82#_c_172_n N_A1_M1003_g 0.0132844f $X=3.265 $Y=1.095 $X2=0 $Y2=0
cc_146 N_A_27_82#_c_174_n N_A1_M1003_g 0.00113123f $X=3.505 $Y=0.865 $X2=0 $Y2=0
cc_147 N_A_27_82#_c_176_n N_A1_c_295_n 0.0039021f $X=2.5 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A_27_82#_c_170_n N_A1_c_295_n 0.00975019f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_149 N_A_27_82#_c_171_n N_A1_c_295_n 0.00344746f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_150 N_A_27_82#_c_172_n N_A1_c_295_n 0.0256551f $X=3.265 $Y=1.095 $X2=0 $Y2=0
cc_151 N_A_27_82#_c_174_n N_B1_c_332_n 0.00197779f $X=3.505 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A_27_82#_c_174_n N_B1_M1009_g 0.0132613f $X=3.505 $Y=0.865 $X2=0 $Y2=0
cc_153 N_A_27_82#_c_174_n N_B1_c_334_n 0.0236445f $X=3.505 $Y=0.865 $X2=0 $Y2=0
cc_154 N_A_27_82#_c_174_n N_B2_M1007_g 2.25597e-19 $X=3.505 $Y=0.865 $X2=0 $Y2=0
cc_155 N_A_27_82#_c_179_n N_A_116_392#_M1013_d 0.00200085f $X=1.355 $Y=2.075
+ $X2=-0.19 $Y2=-0.245
cc_156 N_A_27_82#_M1012_d N_A_116_392#_c_417_n 0.00818441f $X=1.03 $Y=1.96 $X2=0
+ $Y2=0
cc_157 N_A_27_82#_c_175_n N_A_116_392#_c_417_n 0.0138924f $X=2.05 $Y=1.765 $X2=0
+ $Y2=0
cc_158 N_A_27_82#_c_176_n N_A_116_392#_c_417_n 0.016816f $X=2.5 $Y=1.765 $X2=0
+ $Y2=0
cc_159 N_A_27_82#_c_179_n N_A_116_392#_c_417_n 0.0437127f $X=1.355 $Y=2.075
+ $X2=0 $Y2=0
cc_160 N_A_27_82#_c_178_n N_A_116_392#_c_418_n 0.0416015f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_27_82#_c_179_n N_A_116_392#_c_418_n 0.0176481f $X=1.355 $Y=2.075
+ $X2=0 $Y2=0
cc_162 N_A_27_82#_c_175_n N_VPWR_c_452_n 0.0156805f $X=2.05 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_27_82#_c_176_n N_VPWR_c_453_n 0.0124283f $X=2.5 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A_27_82#_c_175_n N_VPWR_c_456_n 0.00461464f $X=2.05 $Y=1.765 $X2=0
+ $Y2=0
cc_165 N_A_27_82#_c_176_n N_VPWR_c_456_n 0.00461464f $X=2.5 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A_27_82#_c_178_n N_VPWR_c_458_n 0.011066f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A_27_82#_c_175_n N_VPWR_c_451_n 0.00456645f $X=2.05 $Y=1.765 $X2=0
+ $Y2=0
cc_168 N_A_27_82#_c_176_n N_VPWR_c_451_n 0.00456645f $X=2.5 $Y=1.765 $X2=0 $Y2=0
cc_169 N_A_27_82#_c_178_n N_VPWR_c_451_n 0.00915947f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_27_82#_c_169_n N_X_M1002_d 0.00435233f $X=2.23 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_171 N_A_27_82#_c_161_n N_X_c_501_n 0.0052405f $X=1.645 $Y=1.26 $X2=0 $Y2=0
cc_172 N_A_27_82#_c_162_n N_X_c_501_n 0.0105762f $X=1.96 $Y=1.335 $X2=0 $Y2=0
cc_173 N_A_27_82#_c_163_n N_X_c_501_n 0.00207346f $X=1.72 $Y=1.335 $X2=0 $Y2=0
cc_174 N_A_27_82#_c_175_n N_X_c_501_n 0.0023312f $X=2.05 $Y=1.765 $X2=0 $Y2=0
cc_175 N_A_27_82#_c_164_n N_X_c_501_n 0.00554882f $X=2.075 $Y=1.26 $X2=0 $Y2=0
cc_176 N_A_27_82#_c_176_n N_X_c_501_n 2.7342e-19 $X=2.5 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A_27_82#_c_168_n N_X_c_501_n 0.0542206f $X=1.44 $Y=1.95 $X2=0 $Y2=0
cc_178 N_A_27_82#_c_169_n N_X_c_501_n 0.0170777f $X=2.23 $Y=0.665 $X2=0 $Y2=0
cc_179 N_A_27_82#_c_248_p N_X_c_501_n 0.00572056f $X=2.315 $Y=1.01 $X2=0 $Y2=0
cc_180 N_A_27_82#_c_170_n N_X_c_501_n 0.0267529f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_181 N_A_27_82#_c_171_n N_X_c_501_n 0.0189862f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_182 N_A_27_82#_c_173_n N_X_c_501_n 0.012203f $X=2.395 $Y=1.095 $X2=0 $Y2=0
cc_183 N_A_27_82#_c_163_n N_X_c_503_n 7.04168e-19 $X=1.72 $Y=1.335 $X2=0 $Y2=0
cc_184 N_A_27_82#_c_175_n N_X_c_503_n 0.0201899f $X=2.05 $Y=1.765 $X2=0 $Y2=0
cc_185 N_A_27_82#_c_176_n N_X_c_503_n 0.00728842f $X=2.5 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A_27_82#_c_179_n N_X_c_503_n 0.0233303f $X=1.355 $Y=2.075 $X2=0 $Y2=0
cc_187 N_A_27_82#_c_168_n N_X_c_503_n 0.0108574f $X=1.44 $Y=1.95 $X2=0 $Y2=0
cc_188 N_A_27_82#_c_170_n N_X_c_503_n 0.0140238f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_189 N_A_27_82#_c_171_n N_X_c_503_n 0.00615917f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_190 N_A_27_82#_c_166_n A_114_82# 0.0048076f $X=1.355 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_191 N_A_27_82#_c_166_n N_VGND_M1011_d 0.0111604f $X=1.355 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_192 N_A_27_82#_c_202_n N_VGND_M1011_d 0.00267073f $X=1.44 $Y=0.92 $X2=-0.19
+ $Y2=-0.245
cc_193 N_A_27_82#_c_168_n N_VGND_M1011_d 0.00133961f $X=1.44 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_194 N_A_27_82#_c_263_p N_VGND_M1011_d 0.00463907f $X=1.525 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_195 N_A_27_82#_c_264_p N_VGND_M1011_d 0.00142544f $X=1.44 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_196 N_A_27_82#_c_169_n N_VGND_M1006_s 0.00562426f $X=2.23 $Y=0.665 $X2=0
+ $Y2=0
cc_197 N_A_27_82#_c_248_p N_VGND_M1006_s 0.011885f $X=2.315 $Y=1.01 $X2=0 $Y2=0
cc_198 N_A_27_82#_c_173_n N_VGND_M1006_s 0.00193901f $X=2.395 $Y=1.095 $X2=0
+ $Y2=0
cc_199 N_A_27_82#_c_161_n N_VGND_c_553_n 0.0062784f $X=1.645 $Y=1.26 $X2=0 $Y2=0
cc_200 N_A_27_82#_c_165_n N_VGND_c_553_n 0.00509935f $X=0.28 $Y=0.555 $X2=0
+ $Y2=0
cc_201 N_A_27_82#_c_166_n N_VGND_c_553_n 0.015373f $X=1.355 $Y=1.005 $X2=0 $Y2=0
cc_202 N_A_27_82#_c_263_p N_VGND_c_553_n 0.0141996f $X=1.525 $Y=0.665 $X2=0
+ $Y2=0
cc_203 N_A_27_82#_c_165_n N_VGND_c_555_n 0.00955085f $X=0.28 $Y=0.555 $X2=0
+ $Y2=0
cc_204 N_A_27_82#_c_164_n N_VGND_c_557_n 0.00546687f $X=2.075 $Y=1.26 $X2=0
+ $Y2=0
cc_205 N_A_27_82#_c_169_n N_VGND_c_557_n 0.0157799f $X=2.23 $Y=0.665 $X2=0 $Y2=0
cc_206 N_A_27_82#_c_173_n N_VGND_c_557_n 0.00480154f $X=2.395 $Y=1.095 $X2=0
+ $Y2=0
cc_207 N_A_27_82#_c_161_n N_VGND_c_558_n 0.00414982f $X=1.645 $Y=1.26 $X2=0
+ $Y2=0
cc_208 N_A_27_82#_c_164_n N_VGND_c_558_n 0.00414982f $X=2.075 $Y=1.26 $X2=0
+ $Y2=0
cc_209 N_A_27_82#_c_169_n N_VGND_c_558_n 0.0113015f $X=2.23 $Y=0.665 $X2=0 $Y2=0
cc_210 N_A_27_82#_c_263_p N_VGND_c_558_n 0.00358211f $X=1.525 $Y=0.665 $X2=0
+ $Y2=0
cc_211 N_A_27_82#_c_161_n N_VGND_c_562_n 0.00533081f $X=1.645 $Y=1.26 $X2=0
+ $Y2=0
cc_212 N_A_27_82#_c_164_n N_VGND_c_562_n 0.00533081f $X=2.075 $Y=1.26 $X2=0
+ $Y2=0
cc_213 N_A_27_82#_c_165_n N_VGND_c_562_n 0.00894475f $X=0.28 $Y=0.555 $X2=0
+ $Y2=0
cc_214 N_A_27_82#_c_169_n N_VGND_c_562_n 0.0210788f $X=2.23 $Y=0.665 $X2=0 $Y2=0
cc_215 N_A_27_82#_c_263_p N_VGND_c_562_n 0.00537088f $X=1.525 $Y=0.665 $X2=0
+ $Y2=0
cc_216 N_A_27_82#_M1003_d N_A_557_74#_c_616_n 0.00478343f $X=3.255 $Y=0.37 $X2=0
+ $Y2=0
cc_217 N_A_27_82#_c_172_n N_A_557_74#_c_616_n 0.00462336f $X=3.265 $Y=1.095
+ $X2=0 $Y2=0
cc_218 N_A_27_82#_c_174_n N_A_557_74#_c_616_n 0.0272186f $X=3.505 $Y=0.865 $X2=0
+ $Y2=0
cc_219 N_A_27_82#_c_174_n N_A_557_74#_c_618_n 0.0146766f $X=3.505 $Y=0.865 $X2=0
+ $Y2=0
cc_220 N_A_27_82#_c_164_n N_A_557_74#_c_620_n 0.00501373f $X=2.075 $Y=1.26 $X2=0
+ $Y2=0
cc_221 N_A_27_82#_c_169_n N_A_557_74#_c_620_n 0.00852177f $X=2.23 $Y=0.665 $X2=0
+ $Y2=0
cc_222 N_A_27_82#_c_248_p N_A_557_74#_c_620_n 0.00405254f $X=2.315 $Y=1.01 $X2=0
+ $Y2=0
cc_223 N_A_27_82#_c_172_n N_A_557_74#_c_620_n 0.0244887f $X=3.265 $Y=1.095 $X2=0
+ $Y2=0
cc_224 N_A1_c_293_n N_B1_c_332_n 0.0461053f $X=3.12 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_225 N_A1_c_295_n N_B1_c_332_n 0.00619734f $X=3.09 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_226 N_A1_M1003_g N_B1_M1009_g 0.0259476f $X=3.18 $Y=0.69 $X2=0 $Y2=0
cc_227 N_A1_c_293_n N_B1_c_334_n 0.00152252f $X=3.12 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A1_c_295_n N_B1_c_334_n 0.0280926f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_229 N_A1_c_293_n N_A_116_392#_c_417_n 0.0147342f $X=3.12 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A1_c_295_n N_A_116_392#_c_417_n 0.0134522f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_231 N_A1_c_293_n N_A_116_392#_c_431_n 0.0011267f $X=3.12 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A1_c_295_n N_A_116_392#_c_431_n 0.00593546f $X=3.09 $Y=1.515 $X2=0
+ $Y2=0
cc_233 N_A1_c_295_n N_VPWR_M1004_s 0.00522949f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_234 N_A1_c_293_n N_VPWR_c_453_n 0.00296264f $X=3.12 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A1_c_293_n N_VPWR_c_459_n 0.0049405f $X=3.12 $Y=1.765 $X2=0 $Y2=0
cc_236 N_A1_c_293_n N_VPWR_c_451_n 0.00508379f $X=3.12 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A1_c_293_n N_X_c_503_n 5.05129e-19 $X=3.12 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A1_c_295_n N_X_c_503_n 0.011999f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_239 N_A1_c_295_n N_A_639_368#_M1008_d 0.00500256f $X=3.09 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_240 N_A1_c_293_n N_A_639_368#_c_532_n 0.00309115f $X=3.12 $Y=1.765 $X2=0
+ $Y2=0
cc_241 N_A1_M1003_g N_VGND_c_557_n 0.00265086f $X=3.18 $Y=0.69 $X2=0 $Y2=0
cc_242 N_A1_M1003_g N_VGND_c_559_n 0.00291649f $X=3.18 $Y=0.69 $X2=0 $Y2=0
cc_243 N_A1_M1003_g N_VGND_c_562_n 0.00365718f $X=3.18 $Y=0.69 $X2=0 $Y2=0
cc_244 N_A1_M1003_g N_A_557_74#_c_616_n 0.0115929f $X=3.18 $Y=0.69 $X2=0 $Y2=0
cc_245 N_A1_M1003_g N_A_557_74#_c_620_n 0.00168345f $X=3.18 $Y=0.69 $X2=0 $Y2=0
cc_246 N_B1_M1009_g N_B2_M1007_g 0.0355648f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_247 N_B1_c_332_n N_B2_c_362_n 0.057175f $X=3.775 $Y=1.765 $X2=0 $Y2=0
cc_248 N_B1_c_334_n N_B2_c_362_n 3.64648e-19 $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_249 N_B1_c_332_n N_B2_c_363_n 0.00318816f $X=3.775 $Y=1.765 $X2=0 $Y2=0
cc_250 N_B1_c_334_n N_B2_c_363_n 0.0350349f $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_251 N_B1_c_332_n N_A_116_392#_c_417_n 0.0173193f $X=3.775 $Y=1.765 $X2=0
+ $Y2=0
cc_252 N_B1_c_334_n N_A_116_392#_c_417_n 0.00928034f $X=3.63 $Y=1.515 $X2=0
+ $Y2=0
cc_253 N_B1_c_332_n N_A_116_392#_c_431_n 0.00971005f $X=3.775 $Y=1.765 $X2=0
+ $Y2=0
cc_254 N_B1_c_332_n N_VPWR_c_459_n 7.26245e-19 $X=3.775 $Y=1.765 $X2=0 $Y2=0
cc_255 N_B1_c_332_n N_A_639_368#_c_530_n 0.00776105f $X=3.775 $Y=1.765 $X2=0
+ $Y2=0
cc_256 N_B1_c_332_n N_A_639_368#_c_532_n 0.00553388f $X=3.775 $Y=1.765 $X2=0
+ $Y2=0
cc_257 N_B1_M1009_g N_VGND_c_554_n 7.59698e-19 $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_258 N_B1_M1009_g N_VGND_c_559_n 0.00291649f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_259 N_B1_M1009_g N_VGND_c_562_n 0.00360429f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_260 N_B1_M1009_g N_A_557_74#_c_616_n 0.0139417f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_261 N_B1_M1009_g N_A_557_74#_c_618_n 0.00130469f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_262 N_B2_M1007_g N_A2_M1015_g 0.0231299f $X=4.19 $Y=0.69 $X2=0 $Y2=0
cc_263 N_B2_c_362_n N_A2_c_395_n 0.048535f $X=4.225 $Y=1.765 $X2=0 $Y2=0
cc_264 N_B2_c_363_n N_A2_c_395_n 8.4048e-19 $X=4.28 $Y=1.515 $X2=0 $Y2=0
cc_265 N_B2_c_362_n A2 5.53912e-19 $X=4.225 $Y=1.765 $X2=0 $Y2=0
cc_266 N_B2_c_363_n A2 0.026473f $X=4.28 $Y=1.515 $X2=0 $Y2=0
cc_267 N_B2_c_362_n N_A_116_392#_c_417_n 0.00378309f $X=4.225 $Y=1.765 $X2=0
+ $Y2=0
cc_268 N_B2_c_362_n N_A_116_392#_c_431_n 0.00494592f $X=4.225 $Y=1.765 $X2=0
+ $Y2=0
cc_269 N_B2_c_363_n N_A_116_392#_c_431_n 0.0148925f $X=4.28 $Y=1.515 $X2=0 $Y2=0
cc_270 N_B2_c_362_n N_VPWR_c_455_n 2.39035e-19 $X=4.225 $Y=1.765 $X2=0 $Y2=0
cc_271 N_B2_c_362_n N_VPWR_c_459_n 7.26245e-19 $X=4.225 $Y=1.765 $X2=0 $Y2=0
cc_272 N_B2_c_362_n N_A_639_368#_c_530_n 0.0112073f $X=4.225 $Y=1.765 $X2=0
+ $Y2=0
cc_273 N_B2_c_362_n N_A_639_368#_c_531_n 0.00777893f $X=4.225 $Y=1.765 $X2=0
+ $Y2=0
cc_274 N_B2_c_363_n N_A_639_368#_c_531_n 0.00869275f $X=4.28 $Y=1.515 $X2=0
+ $Y2=0
cc_275 N_B2_M1007_g N_VGND_c_554_n 0.00890008f $X=4.19 $Y=0.69 $X2=0 $Y2=0
cc_276 N_B2_M1007_g N_VGND_c_559_n 0.00444681f $X=4.19 $Y=0.69 $X2=0 $Y2=0
cc_277 N_B2_M1007_g N_VGND_c_562_n 0.00877228f $X=4.19 $Y=0.69 $X2=0 $Y2=0
cc_278 N_B2_M1007_g N_A_557_74#_c_616_n 7.44093e-19 $X=4.19 $Y=0.69 $X2=0 $Y2=0
cc_279 N_B2_M1007_g N_A_557_74#_c_617_n 0.0147396f $X=4.19 $Y=0.69 $X2=0 $Y2=0
cc_280 N_B2_c_362_n N_A_557_74#_c_617_n 0.00418988f $X=4.225 $Y=1.765 $X2=0
+ $Y2=0
cc_281 N_B2_c_363_n N_A_557_74#_c_617_n 0.0267388f $X=4.28 $Y=1.515 $X2=0 $Y2=0
cc_282 N_B2_c_363_n N_A_557_74#_c_618_n 0.011271f $X=4.28 $Y=1.515 $X2=0 $Y2=0
cc_283 N_B2_M1007_g N_A_557_74#_c_619_n 9.43881e-19 $X=4.19 $Y=0.69 $X2=0 $Y2=0
cc_284 N_A2_c_395_n N_VPWR_c_455_n 0.0176177f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_285 A2 N_VPWR_c_455_n 0.0255179f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_286 N_A2_c_395_n N_VPWR_c_459_n 0.00443511f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_287 N_A2_c_395_n N_VPWR_c_451_n 0.00460931f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_288 N_A2_c_395_n N_A_639_368#_c_530_n 6.49559e-19 $X=4.775 $Y=1.765 $X2=0
+ $Y2=0
cc_289 N_A2_c_395_n N_A_639_368#_c_531_n 0.00589778f $X=4.775 $Y=1.765 $X2=0
+ $Y2=0
cc_290 N_A2_M1015_g N_VGND_c_554_n 0.00752319f $X=4.76 $Y=0.69 $X2=0 $Y2=0
cc_291 N_A2_M1015_g N_VGND_c_561_n 0.00434272f $X=4.76 $Y=0.69 $X2=0 $Y2=0
cc_292 N_A2_M1015_g N_VGND_c_562_n 0.00826173f $X=4.76 $Y=0.69 $X2=0 $Y2=0
cc_293 N_A2_M1015_g N_A_557_74#_c_617_n 0.0159753f $X=4.76 $Y=0.69 $X2=0 $Y2=0
cc_294 N_A2_c_395_n N_A_557_74#_c_617_n 0.00426868f $X=4.775 $Y=1.765 $X2=0
+ $Y2=0
cc_295 A2 N_A_557_74#_c_617_n 0.0378526f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_296 N_A2_M1015_g N_A_557_74#_c_619_n 0.00970393f $X=4.76 $Y=0.69 $X2=0 $Y2=0
cc_297 N_A_116_392#_c_417_n N_VPWR_M1000_s 0.00530189f $X=3.835 $Y=2.455
+ $X2=-0.19 $Y2=1.66
cc_298 N_A_116_392#_c_417_n N_VPWR_M1004_s 0.0168889f $X=3.835 $Y=2.455 $X2=0
+ $Y2=0
cc_299 N_A_116_392#_c_417_n N_VPWR_c_452_n 0.0264652f $X=3.835 $Y=2.455 $X2=0
+ $Y2=0
cc_300 N_A_116_392#_c_417_n N_VPWR_c_453_n 0.0260584f $X=3.835 $Y=2.455 $X2=0
+ $Y2=0
cc_301 N_A_116_392#_c_418_n N_VPWR_c_458_n 0.0144379f $X=0.73 $Y=2.455 $X2=0
+ $Y2=0
cc_302 N_A_116_392#_c_417_n N_VPWR_c_451_n 0.0616189f $X=3.835 $Y=2.455 $X2=0
+ $Y2=0
cc_303 N_A_116_392#_c_418_n N_VPWR_c_451_n 0.0119346f $X=0.73 $Y=2.455 $X2=0
+ $Y2=0
cc_304 N_A_116_392#_c_417_n N_X_M1000_d 0.00556049f $X=3.835 $Y=2.455 $X2=0
+ $Y2=0
cc_305 N_A_116_392#_c_417_n N_X_c_503_n 0.043448f $X=3.835 $Y=2.455 $X2=0 $Y2=0
cc_306 N_A_116_392#_c_417_n N_A_639_368#_M1008_d 0.0167516f $X=3.835 $Y=2.455
+ $X2=-0.19 $Y2=1.66
cc_307 N_A_116_392#_c_417_n N_A_639_368#_c_530_n 0.026807f $X=3.835 $Y=2.455
+ $X2=0 $Y2=0
cc_308 N_A_116_392#_c_417_n N_A_639_368#_c_532_n 0.0290159f $X=3.835 $Y=2.455
+ $X2=0 $Y2=0
cc_309 N_VPWR_M1000_s N_X_c_503_n 0.00387385f $X=1.595 $Y=2.73 $X2=0 $Y2=0
cc_310 N_VPWR_c_455_n N_A_639_368#_c_530_n 0.0147692f $X=5 $Y=2.115 $X2=0 $Y2=0
cc_311 N_VPWR_c_459_n N_A_639_368#_c_530_n 0.0690424f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_451_n N_A_639_368#_c_530_n 0.0393321f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_455_n N_A_639_368#_c_531_n 0.038455f $X=5 $Y=2.115 $X2=0 $Y2=0
cc_314 N_VPWR_c_453_n N_A_639_368#_c_532_n 0.0206835f $X=2.81 $Y=2.875 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_459_n N_A_639_368#_c_532_n 0.0248486f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_451_n N_A_639_368#_c_532_n 0.0138941f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_317 N_VGND_c_554_n N_A_557_74#_c_616_n 0.00729485f $X=4.425 $Y=0.635 $X2=0
+ $Y2=0
cc_318 N_VGND_c_559_n N_A_557_74#_c_616_n 0.0401161f $X=4.26 $Y=0 $X2=0 $Y2=0
cc_319 N_VGND_c_562_n N_A_557_74#_c_616_n 0.0340164f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_320 N_VGND_c_554_n N_A_557_74#_c_617_n 0.0245379f $X=4.425 $Y=0.635 $X2=0
+ $Y2=0
cc_321 N_VGND_c_554_n N_A_557_74#_c_619_n 0.0312316f $X=4.425 $Y=0.635 $X2=0
+ $Y2=0
cc_322 N_VGND_c_561_n N_A_557_74#_c_619_n 0.0145639f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_323 N_VGND_c_562_n N_A_557_74#_c_619_n 0.0119984f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_324 N_VGND_c_557_n N_A_557_74#_c_620_n 0.00404517f $X=2.37 $Y=0 $X2=0 $Y2=0
cc_325 N_VGND_c_559_n N_A_557_74#_c_620_n 0.0142934f $X=4.26 $Y=0 $X2=0 $Y2=0
cc_326 N_VGND_c_562_n N_A_557_74#_c_620_n 0.0119825f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_327 N_A_557_74#_c_653_p A_775_74# 9.797e-19 $X=4.005 $Y=1.01 $X2=-0.19
+ $Y2=-0.245
