* File: sky130_fd_sc_ls__a22o_4.spice
* Created: Wed Sep  2 10:50:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a22o_4.pex.spice"
.subckt sky130_fd_sc_ls__a22o_4  VNB VPB B2 B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1002 N_X_M1002_d N_A_95_306#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75004.8 A=0.111 P=1.78 MULT=1
MM1004 N_X_M1002_d N_A_95_306#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75004.4 A=0.111 P=1.78 MULT=1
MM1017 N_X_M1017_d N_A_95_306#_M1017_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75003.9 A=0.111 P=1.78 MULT=1
MM1020 N_X_M1017_d N_A_95_306#_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.136042 PD=1.02 PS=1.17435 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1020_s N_B2_M1021_g N_A_645_120#_M1021_s VNB NSHORT L=0.15 W=0.64
+ AD=0.117658 AS=0.0896 PD=1.01565 PS=0.92 NRD=14.052 NRS=0 M=1 R=4.26667
+ SA=75002 SB=75003.5 A=0.096 P=1.58 MULT=1
MM1000 N_A_95_306#_M1000_d N_B1_M1000_g N_A_645_120#_M1021_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.4 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1018 N_A_95_306#_M1000_d N_B1_M1018_g N_A_645_120#_M1018_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.105312 PD=0.92 PS=0.98 NRD=0 NRS=3.744 M=1 R=4.26667
+ SA=75002.8 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1023 N_VGND_M1023_d N_B2_M1023_g N_A_645_120#_M1018_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1952 AS=0.105312 PD=1.25 PS=0.98 NRD=0 NRS=4.68 M=1 R=4.26667 SA=75003.2
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1001 N_A_1064_123#_M1001_d N_A2_M1001_g N_VGND_M1023_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1952 PD=0.92 PS=1.25 NRD=0 NRS=61.872 M=1 R=4.26667
+ SA=75004 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1003 N_A_95_306#_M1003_d N_A1_M1003_g N_A_1064_123#_M1001_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.4 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1016 N_A_95_306#_M1003_d N_A1_M1016_g N_A_1064_123#_M1016_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.9 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1022 N_A_1064_123#_M1016_s N_A2_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75005.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_X_M1007_d N_A_95_306#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1008 N_X_M1007_d N_A_95_306#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1013 N_X_M1013_d N_A_95_306#_M1013_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1019 N_X_M1013_d N_A_95_306#_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1009 N_A_95_306#_M1009_d N_B2_M1009_g N_A_555_392#_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75003.6 A=0.15 P=2.3 MULT=1
MM1010 N_A_95_306#_M1009_d N_B1_M1010_g N_A_555_392#_M1010_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.6 SB=75003.1 A=0.15 P=2.3 MULT=1
MM1014 N_A_95_306#_M1014_d N_B1_M1014_g N_A_555_392#_M1010_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1015 N_A_95_306#_M1014_d N_B2_M1015_g N_A_555_392#_M1015_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.165 PD=1.3 PS=1.33 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.5 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A2_M1006_g N_A_555_392#_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2575 AS=0.165 PD=1.515 PS=1.33 NRD=19.7 NRS=7.8603 M=1 R=6.66667 SA=75002
+ SB=75001.8 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1006_d N_A1_M1005_g N_A_555_392#_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2575 AS=0.15 PD=1.515 PS=1.3 NRD=26.5753 NRS=1.9503 M=1 R=6.66667
+ SA=75002.7 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_A1_M1011_g N_A_555_392#_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75003.1
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1011_d N_A2_M1012_g N_A_555_392#_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75003.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=14.0988 P=18.88
*
.include "sky130_fd_sc_ls__a22o_4.pxi.spice"
*
.ends
*
*
