* File: sky130_fd_sc_ls__or2_2.pex.spice
* Created: Fri Aug 28 13:57:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__OR2_2%B 1 3 4 6 7
c23 7 0 1.41453e-19 $X=0.24 $Y=1.295
c24 1 0 1.44963e-19 $X=0.49 $Y=1.22
r25 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r26 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r27 4 10 67.6304 $w=3.61e-07 $l=4.48776e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.345 $Y2=1.385
r28 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.34
r29 1 10 38.924 $w=3.61e-07 $l=2.26164e-07 $layer=POLY_cond $X=0.49 $Y=1.22
+ $X2=0.345 $Y2=1.385
r30 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.49 $Y=1.22 $X2=0.49
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_2%A 1 3 6 8 9 14
c41 1 0 1.41453e-19 $X=0.885 $Y=1.765
r42 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=1.515 $X2=0.96 $Y2=1.515
r43 8 9 9.691 $w=4.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.825 $Y=1.665 $X2=0.825
+ $Y2=2.035
r44 8 14 3.92878 $w=4.38e-07 $l=1.5e-07 $layer=LI1_cond $X=0.825 $Y=1.665
+ $X2=0.825 $Y2=1.515
r45 4 13 38.5562 $w=2.99e-07 $l=1.83916e-07 $layer=POLY_cond $X=0.92 $Y=1.35
+ $X2=0.96 $Y2=1.515
r46 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.92 $Y=1.35 $X2=0.92
+ $Y2=0.79
r47 1 13 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.885 $Y=1.765
+ $X2=0.96 $Y2=1.515
r48 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.885 $Y=1.765
+ $X2=0.885 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_2%A_27_368# 1 2 9 11 13 16 18 20 23 27 29 33 35
+ 36 38 39 42 43 44 46 52
c97 33 0 1.44963e-19 $X=0.705 $Y=0.615
r98 51 52 5.07368 $w=3.8e-07 $l=4e-08 $layer=POLY_cond $X=1.855 $Y=1.532
+ $X2=1.895 $Y2=1.532
r99 50 51 54.5421 $w=3.8e-07 $l=4.3e-07 $layer=POLY_cond $X=1.425 $Y=1.532
+ $X2=1.855 $Y2=1.532
r100 47 52 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=2.13 $Y=1.532
+ $X2=1.895 $Y2=1.532
r101 46 49 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.13 $Y=1.465
+ $X2=2.13 $Y2=1.63
r102 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.465 $X2=2.13 $Y2=1.465
r103 42 49 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.21 $Y=2.32
+ $X2=2.21 $Y2=1.63
r104 40 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.385 $Y=2.405
+ $X2=1.3 $Y2=2.405
r105 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.125 $Y=2.405
+ $X2=2.21 $Y2=2.32
r106 39 40 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.125 $Y=2.405
+ $X2=1.385 $Y2=2.405
r107 38 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=2.32 $X2=1.3
+ $Y2=2.405
r108 37 38 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=1.3 $Y=1.18
+ $X2=1.3 $Y2=2.32
r109 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.215 $Y=1.095
+ $X2=1.3 $Y2=1.18
r110 35 36 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.215 $Y=1.095
+ $X2=0.87 $Y2=1.095
r111 31 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.745 $Y=1.01
+ $X2=0.87 $Y2=1.095
r112 31 33 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=0.745 $Y=1.01
+ $X2=0.745 $Y2=0.615
r113 30 43 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=2.405
+ $X2=0.27 $Y2=2.405
r114 29 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=2.405
+ $X2=1.3 $Y2=2.405
r115 29 30 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.215 $Y=2.405
+ $X2=0.435 $Y2=2.405
r116 25 43 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.49
+ $X2=0.27 $Y2=2.405
r117 25 27 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.27 $Y=2.49
+ $X2=0.27 $Y2=2.695
r118 21 43 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.32
+ $X2=0.27 $Y2=2.405
r119 21 23 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.27 $Y=2.32
+ $X2=0.27 $Y2=1.985
r120 18 52 24.6126 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.895 $Y=1.765
+ $X2=1.895 $Y2=1.532
r121 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.895 $Y=1.765
+ $X2=1.895 $Y2=2.4
r122 14 51 24.6126 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.855 $Y=1.3
+ $X2=1.855 $Y2=1.532
r123 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.855 $Y=1.3
+ $X2=1.855 $Y2=0.74
r124 11 50 24.6126 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.425 $Y=1.765
+ $X2=1.425 $Y2=1.532
r125 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.425 $Y=1.765
+ $X2=1.425 $Y2=2.4
r126 7 50 24.6126 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.425 $Y=1.3
+ $X2=1.425 $Y2=1.532
r127 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.425 $Y=1.3
+ $X2=1.425 $Y2=0.74
r128 2 27 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.695
r129 2 23 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=1.985
r130 1 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.47 $X2=0.705 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_2%VPWR 1 2 9 11 13 15 17 22 28 32
r36 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 23 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=3.33
+ $X2=1.2 $Y2=3.33
r40 23 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.365 $Y=3.33
+ $X2=1.68 $Y2=3.33
r41 22 31 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=2.177 $Y2=3.33
r42 22 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 17 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 17 19 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 15 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 11 31 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.177 $Y2=3.33
r50 11 13 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=2.78
r51 7 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=3.245 $X2=1.2
+ $Y2=3.33
r52 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.2 $Y=3.245 $X2=1.2
+ $Y2=2.78
r53 2 13 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=1.84 $X2=2.12 $Y2=2.78
r54 1 9 600 $w=1.7e-07 $l=1.05319e-06 $layer=licon1_PDIFF $count=1 $X=0.96
+ $Y=1.84 $X2=1.2 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_2%X 1 2 7 8 9 10 11
r21 11 30 7.05875 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.695 $Y=1.985
+ $X2=1.695 $Y2=1.82
r22 10 30 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=1.675 $Y=1.665
+ $X2=1.675 $Y2=1.82
r23 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.675 $Y=1.295
+ $X2=1.675 $Y2=1.665
r24 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.675 $Y=0.925
+ $X2=1.675 $Y2=1.295
r25 7 8 19.6876 $w=2.38e-07 $l=4.1e-07 $layer=LI1_cond $X=1.675 $Y=0.515
+ $X2=1.675 $Y2=0.925
r26 2 11 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.84 $X2=1.66 $Y2=1.985
r27 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.5 $Y=0.37
+ $X2=1.64 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_2%VGND 1 2 3 10 12 16 18 20 22 24 29 38 42
r37 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 33 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r40 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r41 30 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.21
+ $Y2=0
r42 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.68
+ $Y2=0
r43 29 41 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.97 $Y=0 $X2=2.185
+ $Y2=0
r44 29 32 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.97 $Y=0 $X2=1.68
+ $Y2=0
r45 28 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r46 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r47 25 35 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.22
+ $Y2=0
r48 25 27 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.72
+ $Y2=0
r49 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.21
+ $Y2=0
r50 24 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.72
+ $Y2=0
r51 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r52 22 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r53 22 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 18 41 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=2.135 $Y=0.085
+ $X2=2.185 $Y2=0
r55 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.135 $Y=0.085
+ $X2=2.135 $Y2=0.515
r56 14 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r57 14 16 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.65
r58 10 35 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.22 $Y2=0
r59 10 12 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.835
r60 3 20 91 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=2 $X=1.93
+ $Y=0.37 $X2=2.135 $Y2=0.515
r61 2 16 182 $w=1.7e-07 $l=2.91419e-07 $layer=licon1_NDIFF $count=1 $X=0.995
+ $Y=0.47 $X2=1.21 $Y2=0.65
r62 1 12 182 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.47 $X2=0.275 $Y2=0.835
.ends

