* File: sky130_fd_sc_ls__and4bb_1.spice
* Created: Fri Aug 28 13:06:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__and4bb_1.pex.spice"
.subckt sky130_fd_sc_ls__and4bb_1  VNB VPB A_N C D B_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B_N	B_N
* D	D
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_A_N_M1012_g N_A_27_74#_M1012_s VNB NSHORT L=0.15 W=0.55
+ AD=0.0964632 AS=0.15675 PD=0.90814 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1002 N_X_M1002_d N_A_179_48#_M1002_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.129787 PD=2.05 PS=1.22186 NRD=0 NRS=7.296 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 A_455_74# N_A_27_74#_M1004_g N_A_179_48#_M1004_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1005 A_533_74# N_A_503_48#_M1005_g A_455_74# VNB NSHORT L=0.15 W=0.64
+ AD=0.1344 AS=0.0768 PD=1.06 PS=0.88 NRD=29.052 NRS=12.18 M=1 R=4.26667
+ SA=75000.6 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1010 A_647_74# N_C_M1010_g A_533_74# VNB NSHORT L=0.15 W=0.64 AD=0.1152
+ AS=0.1344 PD=1 PS=1.06 NRD=23.436 NRS=29.052 M=1 R=4.26667 SA=75001.2
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1000_d N_D_M1000_g A_647_74# VNB NSHORT L=0.15 W=0.64 AD=0.163308
+ AS=0.1152 PD=1.21008 PS=1 NRD=11.244 NRS=23.436 M=1 R=4.26667 SA=75001.7
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1007 N_A_503_48#_M1007_d N_B_N_M1007_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.55
+ AD=0.15675 AS=0.140342 PD=1.67 PS=1.03992 NRD=0 NRS=32.724 M=1 R=3.66667
+ SA=75002.3 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1008 N_VPWR_M1008_d N_A_N_M1008_g N_A_27_74#_M1008_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.174 AS=0.2478 PD=1.29 PS=2.27 NRD=35.6767 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75000.9 A=0.126 P=1.98 MULT=1
MM1011 N_X_M1011_d N_A_179_48#_M1011_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.4816 AS=0.232 PD=3.1 PS=1.72 NRD=13.1793 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75000.4 A=0.168 P=2.54 MULT=1
MM1009 N_A_179_48#_M1009_d N_A_27_74#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.147 AS=0.2478 PD=1.19 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1013 N_VPWR_M1013_d N_A_503_48#_M1013_g N_A_179_48#_M1009_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.168 AS=0.147 PD=1.24 PS=1.19 NRD=14.0658 NRS=2.3443 M=1 R=5.6
+ SA=75000.7 SB=75001.8 A=0.126 P=1.98 MULT=1
MM1001 N_A_179_48#_M1001_d N_C_M1001_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.168 PD=1.14 PS=1.24 NRD=2.3443 NRS=14.0658 M=1 R=5.6 SA=75001.3
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1006 N_VPWR_M1006_d N_D_M1006_g N_A_179_48#_M1001_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1764 AS=0.126 PD=1.26 PS=1.14 NRD=18.7544 NRS=2.3443 M=1 R=5.6 SA=75001.7
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1003 N_A_503_48#_M1003_d N_B_N_M1003_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2478 AS=0.1764 PD=2.27 PS=1.26 NRD=2.3443 NRS=14.0658 M=1 R=5.6
+ SA=75002.3 SB=75000.2 A=0.126 P=1.98 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
c_96 VPB 0 1.20215e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__and4bb_1.pxi.spice"
*
.ends
*
*
