* File: sky130_fd_sc_ls__nor2_1.spice
* Created: Wed Sep  2 11:13:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nor2_1.pex.spice"
.subckt sky130_fd_sc_ls__nor2_1  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_A_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75000.6
+ A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_B_M1002_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.74 AD=0.2109
+ AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1001 A_116_368# N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.12 AD=0.1512
+ AS=0.3304 PD=1.39 PS=2.83 NRD=14.0658 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75000.6 A=0.168 P=2.54 MULT=1
MM1000 N_Y_M1000_d N_B_M1000_g A_116_368# VPB PHIGHVT L=0.15 W=1.12 AD=0.3304
+ AS=0.1512 PD=2.83 PS=1.39 NRD=1.7533 NRS=14.0658 M=1 R=7.46667 SA=75000.6
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.3852 P=7.36
*
.include "sky130_fd_sc_ls__nor2_1.pxi.spice"
*
.ends
*
*
