* File: sky130_fd_sc_ls__nor3_4.spice
* Created: Wed Sep  2 11:14:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nor3_4.pex.spice"
.subckt sky130_fd_sc_ls__nor3_4  VNB VPB A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.74 AD=0.2109
+ AS=0.1073 PD=2.05 PS=1.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75002.9
+ A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_A_M1014_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.74 AD=0.1517
+ AS=0.1073 PD=1.15 PS=1.03 NRD=9.72 NRS=1.62 M=1 R=4.93333 SA=75000.6
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1517 PD=1.02 PS=1.15 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.2 SB=75001.9
+ A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1003_d N_B_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.6 SB=75001.5
+ A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_C_M1001_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.2 SB=75000.9
+ A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1001_d N_C_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.40425 PD=1.02 PS=2.58 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.6 SB=75000.5
+ A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_27_368#_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3248 PD=1.42 PS=2.82 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75005.9 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1000_d N_A_M1004_g N_A_27_368#_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75005.5 A=0.168 P=2.54 MULT=1
MM1008 N_A_27_368#_M1004_s N_B_M1008_g N_A_295_368#_M1008_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.2713 PD=1.42 PS=1.695 NRD=1.7533 NRS=16.7056 M=1
+ R=7.46667 SA=75001.1 SB=75005 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1006_d N_C_M1006_g N_A_295_368#_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.26145 AS=0.2713 PD=1.64 PS=1.695 NRD=15.8191 NRS=15.8191 M=1 R=7.46667
+ SA=75001.7 SB=75004.4 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1006_d N_C_M1007_g N_A_295_368#_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.26145 AS=0.2744 PD=1.64 PS=1.7 NRD=15.8191 NRS=16.7056 M=1 R=7.46667
+ SA=75002.3 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1012 N_Y_M1012_d N_C_M1012_g N_A_295_368#_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.26145 AS=0.2744 PD=1.64 PS=1.7 NRD=15.8191 NRS=16.7056 M=1 R=7.46667
+ SA=75002.9 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1017 N_Y_M1012_d N_C_M1017_g N_A_295_368#_M1017_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.26145 AS=0.2744 PD=1.64 PS=1.7 NRD=15.8191 NRS=16.7056 M=1 R=7.46667
+ SA=75003.5 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1013 N_A_27_368#_M1013_d N_B_M1013_g N_A_295_368#_M1017_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.2744 PD=1.42 PS=1.7 NRD=1.7533 NRS=16.7056 M=1 R=7.46667
+ SA=75004.1 SB=75002 A=0.168 P=2.54 MULT=1
MM1015 N_A_27_368#_M1013_d N_B_M1015_g N_A_295_368#_M1015_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.6 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1016 N_A_27_368#_M1016_d N_B_M1016_g N_A_295_368#_M1015_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1010 N_VPWR_M1010_d N_A_M1010_g N_A_27_368#_M1016_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.5 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1010_d N_A_M1011_g N_A_27_368#_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.9 SB=75000.2 A=0.168 P=2.54 MULT=1
DX18_noxref VNB VPB NWDIODE A=13.3495 P=18.06
c_107 VPB 0 3.61225e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__nor3_4.pxi.spice"
*
.ends
*
*
