* File: sky130_fd_sc_ls__dfrtp_1.pxi.spice
* Created: Wed Sep  2 11:01:06 2020
* 
x_PM_SKY130_FD_SC_LS__DFRTP_1%D N_D_c_238_n N_D_c_243_n N_D_c_244_n N_D_M1018_g
+ N_D_M1020_g D D D N_D_c_240_n N_D_c_241_n N_D_c_246_n
+ PM_SKY130_FD_SC_LS__DFRTP_1%D
x_PM_SKY130_FD_SC_LS__DFRTP_1%CLK N_CLK_M1006_g N_CLK_M1030_g CLK N_CLK_c_274_n
+ N_CLK_c_275_n PM_SKY130_FD_SC_LS__DFRTP_1%CLK
x_PM_SKY130_FD_SC_LS__DFRTP_1%A_490_390# N_A_490_390#_M1025_d
+ N_A_490_390#_M1011_d N_A_490_390#_c_321_n N_A_490_390#_c_343_n
+ N_A_490_390#_M1009_g N_A_490_390#_c_322_n N_A_490_390#_c_323_n
+ N_A_490_390#_M1027_g N_A_490_390#_c_325_n N_A_490_390#_M1022_g
+ N_A_490_390#_c_326_n N_A_490_390#_c_327_n N_A_490_390#_c_346_n
+ N_A_490_390#_M1001_g N_A_490_390#_c_347_n N_A_490_390#_c_328_n
+ N_A_490_390#_c_329_n N_A_490_390#_c_330_n N_A_490_390#_c_353_p
+ N_A_490_390#_c_331_n N_A_490_390#_c_332_n N_A_490_390#_c_333_n
+ N_A_490_390#_c_334_n N_A_490_390#_c_335_n N_A_490_390#_c_336_n
+ N_A_490_390#_c_337_n N_A_490_390#_c_338_n N_A_490_390#_c_339_n
+ N_A_490_390#_c_340_n N_A_490_390#_c_341_n
+ PM_SKY130_FD_SC_LS__DFRTP_1%A_490_390#
x_PM_SKY130_FD_SC_LS__DFRTP_1%A_830_359# N_A_830_359#_M1026_d
+ N_A_830_359#_M1005_d N_A_830_359#_c_527_n N_A_830_359#_M1003_g
+ N_A_830_359#_M1012_g N_A_830_359#_c_524_n N_A_830_359#_c_542_n
+ N_A_830_359#_c_544_n N_A_830_359#_c_530_n N_A_830_359#_c_525_n
+ N_A_830_359#_c_526_n PM_SKY130_FD_SC_LS__DFRTP_1%A_830_359#
x_PM_SKY130_FD_SC_LS__DFRTP_1%RESET_B N_RESET_B_M1008_g N_RESET_B_c_607_n
+ N_RESET_B_c_617_n N_RESET_B_M1000_g N_RESET_B_c_608_n N_RESET_B_c_609_n
+ N_RESET_B_M1004_g N_RESET_B_c_618_n N_RESET_B_M1029_g N_RESET_B_c_611_n
+ N_RESET_B_M1028_g N_RESET_B_c_621_n N_RESET_B_M1010_g N_RESET_B_c_622_n
+ N_RESET_B_c_613_n N_RESET_B_c_623_n N_RESET_B_c_624_n N_RESET_B_c_625_n
+ N_RESET_B_c_626_n N_RESET_B_c_627_n N_RESET_B_c_628_n RESET_B
+ N_RESET_B_c_614_n N_RESET_B_c_615_n N_RESET_B_c_630_n N_RESET_B_c_631_n
+ N_RESET_B_c_632_n PM_SKY130_FD_SC_LS__DFRTP_1%RESET_B
x_PM_SKY130_FD_SC_LS__DFRTP_1%A_695_457# N_A_695_457#_M1031_d
+ N_A_695_457#_M1009_d N_A_695_457#_M1029_d N_A_695_457#_M1026_g
+ N_A_695_457#_c_833_n N_A_695_457#_M1005_g N_A_695_457#_c_827_n
+ N_A_695_457#_c_861_n N_A_695_457#_c_828_n N_A_695_457#_c_829_n
+ N_A_695_457#_c_830_n N_A_695_457#_c_831_n N_A_695_457#_c_837_n
+ N_A_695_457#_c_832_n N_A_695_457#_c_838_n N_A_695_457#_c_839_n
+ N_A_695_457#_c_875_n PM_SKY130_FD_SC_LS__DFRTP_1%A_695_457#
x_PM_SKY130_FD_SC_LS__DFRTP_1%A_306_96# N_A_306_96#_M1030_s N_A_306_96#_M1006_s
+ N_A_306_96#_M1011_g N_A_306_96#_c_952_n N_A_306_96#_M1025_g
+ N_A_306_96#_c_964_n N_A_306_96#_c_965_n N_A_306_96#_c_966_n
+ N_A_306_96#_c_953_n N_A_306_96#_c_954_n N_A_306_96#_c_955_n
+ N_A_306_96#_M1031_g N_A_306_96#_M1019_g N_A_306_96#_c_969_n
+ N_A_306_96#_M1015_g N_A_306_96#_c_956_n N_A_306_96#_c_957_n
+ N_A_306_96#_M1016_g N_A_306_96#_c_973_n N_A_306_96#_c_974_n
+ N_A_306_96#_c_959_n N_A_306_96#_c_960_n N_A_306_96#_c_989_n
+ N_A_306_96#_c_961_n N_A_306_96#_c_976_n N_A_306_96#_c_1035_n
+ N_A_306_96#_c_962_n PM_SKY130_FD_SC_LS__DFRTP_1%A_306_96#
x_PM_SKY130_FD_SC_LS__DFRTP_1%A_1518_203# N_A_1518_203#_M1017_d
+ N_A_1518_203#_M1010_d N_A_1518_203#_c_1149_n N_A_1518_203#_c_1150_n
+ N_A_1518_203#_c_1151_n N_A_1518_203#_M1024_g N_A_1518_203#_M1014_g
+ N_A_1518_203#_c_1142_n N_A_1518_203#_c_1143_n N_A_1518_203#_c_1144_n
+ N_A_1518_203#_c_1153_n N_A_1518_203#_c_1154_n N_A_1518_203#_c_1145_n
+ N_A_1518_203#_c_1146_n N_A_1518_203#_c_1147_n N_A_1518_203#_c_1156_n
+ N_A_1518_203#_c_1157_n N_A_1518_203#_c_1148_n
+ PM_SKY130_FD_SC_LS__DFRTP_1%A_1518_203#
x_PM_SKY130_FD_SC_LS__DFRTP_1%A_1266_74# N_A_1266_74#_M1022_d
+ N_A_1266_74#_M1015_d N_A_1266_74#_M1017_g N_A_1266_74#_c_1274_n
+ N_A_1266_74#_c_1275_n N_A_1266_74#_M1021_g N_A_1266_74#_c_1261_n
+ N_A_1266_74#_c_1262_n N_A_1266_74#_c_1263_n N_A_1266_74#_c_1278_n
+ N_A_1266_74#_c_1279_n N_A_1266_74#_M1013_g N_A_1266_74#_c_1264_n
+ N_A_1266_74#_c_1265_n N_A_1266_74#_c_1266_n N_A_1266_74#_M1023_g
+ N_A_1266_74#_c_1267_n N_A_1266_74#_c_1287_n N_A_1266_74#_c_1268_n
+ N_A_1266_74#_c_1281_n N_A_1266_74#_c_1269_n N_A_1266_74#_c_1303_n
+ N_A_1266_74#_c_1404_p N_A_1266_74#_c_1282_n N_A_1266_74#_c_1270_n
+ N_A_1266_74#_c_1271_n N_A_1266_74#_c_1272_n N_A_1266_74#_c_1273_n
+ PM_SKY130_FD_SC_LS__DFRTP_1%A_1266_74#
x_PM_SKY130_FD_SC_LS__DFRTP_1%A_1864_409# N_A_1864_409#_M1023_d
+ N_A_1864_409#_M1013_d N_A_1864_409#_c_1426_n N_A_1864_409#_M1007_g
+ N_A_1864_409#_M1002_g N_A_1864_409#_c_1422_n N_A_1864_409#_c_1423_n
+ N_A_1864_409#_c_1429_n N_A_1864_409#_c_1424_n N_A_1864_409#_c_1425_n
+ PM_SKY130_FD_SC_LS__DFRTP_1%A_1864_409#
x_PM_SKY130_FD_SC_LS__DFRTP_1%VPWR N_VPWR_M1018_s N_VPWR_M1000_d N_VPWR_M1006_d
+ N_VPWR_M1003_d N_VPWR_M1005_s N_VPWR_M1024_d N_VPWR_M1021_d N_VPWR_M1007_d
+ N_VPWR_c_1476_n N_VPWR_c_1477_n N_VPWR_c_1478_n N_VPWR_c_1479_n
+ N_VPWR_c_1480_n N_VPWR_c_1481_n N_VPWR_c_1482_n N_VPWR_c_1483_n
+ N_VPWR_c_1484_n N_VPWR_c_1485_n N_VPWR_c_1486_n N_VPWR_c_1487_n VPWR
+ N_VPWR_c_1488_n N_VPWR_c_1489_n N_VPWR_c_1490_n N_VPWR_c_1491_n
+ N_VPWR_c_1492_n N_VPWR_c_1493_n N_VPWR_c_1494_n N_VPWR_c_1495_n
+ N_VPWR_c_1496_n N_VPWR_c_1497_n N_VPWR_c_1498_n N_VPWR_c_1475_n
+ PM_SKY130_FD_SC_LS__DFRTP_1%VPWR
x_PM_SKY130_FD_SC_LS__DFRTP_1%A_30_78# N_A_30_78#_M1020_s N_A_30_78#_M1031_s
+ N_A_30_78#_M1018_d N_A_30_78#_M1009_s N_A_30_78#_c_1624_n N_A_30_78#_c_1631_n
+ N_A_30_78#_c_1625_n N_A_30_78#_c_1633_n N_A_30_78#_c_1634_n
+ N_A_30_78#_c_1635_n N_A_30_78#_c_1626_n N_A_30_78#_c_1636_n
+ N_A_30_78#_c_1627_n N_A_30_78#_c_1628_n N_A_30_78#_c_1638_n
+ N_A_30_78#_c_1639_n N_A_30_78#_c_1629_n N_A_30_78#_c_1630_n
+ PM_SKY130_FD_SC_LS__DFRTP_1%A_30_78#
x_PM_SKY130_FD_SC_LS__DFRTP_1%Q N_Q_M1002_s N_Q_M1007_s N_Q_c_1761_n
+ N_Q_c_1762_n Q Q Q N_Q_c_1763_n PM_SKY130_FD_SC_LS__DFRTP_1%Q
x_PM_SKY130_FD_SC_LS__DFRTP_1%VGND N_VGND_M1008_d N_VGND_M1030_d N_VGND_M1004_d
+ N_VGND_M1014_d N_VGND_M1023_s N_VGND_M1002_d N_VGND_c_1791_n N_VGND_c_1792_n
+ N_VGND_c_1793_n N_VGND_c_1794_n N_VGND_c_1795_n N_VGND_c_1796_n
+ N_VGND_c_1797_n N_VGND_c_1798_n VGND N_VGND_c_1799_n N_VGND_c_1800_n
+ N_VGND_c_1801_n N_VGND_c_1802_n N_VGND_c_1803_n N_VGND_c_1804_n
+ N_VGND_c_1805_n N_VGND_c_1806_n N_VGND_c_1807_n
+ PM_SKY130_FD_SC_LS__DFRTP_1%VGND
cc_1 VNB N_D_c_238_n 0.0406028f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.828
cc_2 VNB N_D_M1020_g 0.0286471f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_3 VNB N_D_c_240_n 0.0216279f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_4 VNB N_D_c_241_n 0.0281582f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_5 VNB CLK 0.00286388f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1
cc_6 VNB N_CLK_c_274_n 0.02183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_CLK_c_275_n 0.0156096f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_A_490_390#_c_321_n 0.00873028f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.75
cc_9 VNB N_A_490_390#_c_322_n 0.0107055f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_A_490_390#_c_323_n 0.022198f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_11 VNB N_A_490_390#_M1027_g 0.0243473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_490_390#_c_325_n 0.0192767f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.165
cc_13 VNB N_A_490_390#_c_326_n 0.0205614f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1
cc_14 VNB N_A_490_390#_c_327_n 0.0110312f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.845
cc_15 VNB N_A_490_390#_c_328_n 0.00232577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_490_390#_c_329_n 0.0343517f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.845
cc_17 VNB N_A_490_390#_c_330_n 0.00301641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_490_390#_c_331_n 0.0169659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_490_390#_c_332_n 9.76919e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_490_390#_c_333_n 0.00385029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_490_390#_c_334_n 0.0019226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_490_390#_c_335_n 0.00257231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_490_390#_c_336_n 0.0129351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_490_390#_c_337_n 0.00403594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_490_390#_c_338_n 0.00385106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_490_390#_c_339_n 0.00724203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_490_390#_c_340_n 0.0313598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_490_390#_c_341_n 0.00797767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_830_359#_M1012_g 0.0345594f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_30 VNB N_A_830_359#_c_524_n 0.00347288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_830_359#_c_525_n 0.00275035f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.295
cc_32 VNB N_A_830_359#_c_526_n 0.00947395f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.845
cc_33 VNB N_RESET_B_M1008_g 0.0204705f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.375
cc_34 VNB N_RESET_B_c_607_n 0.0251526f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.75
cc_35 VNB N_RESET_B_c_608_n 0.280422f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_36 VNB N_RESET_B_c_609_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_37 VNB N_RESET_B_M1004_g 0.0323607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_RESET_B_c_611_n 0.0197602f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.845
cc_39 VNB N_RESET_B_M1028_g 0.0510668f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=2.01
cc_40 VNB N_RESET_B_c_613_n 0.0134203f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.035
cc_41 VNB N_RESET_B_c_614_n 0.0348755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_RESET_B_c_615_n 0.00330649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_695_457#_M1026_g 0.0231233f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_44 VNB N_A_695_457#_c_827_n 0.00347163f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.845
cc_45 VNB N_A_695_457#_c_828_n 0.00148166f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.165
cc_46 VNB N_A_695_457#_c_829_n 0.00289685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_695_457#_c_830_n 0.00804496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_695_457#_c_831_n 0.0411633f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.665
cc_49 VNB N_A_695_457#_c_832_n 0.00235244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_306_96#_c_952_n 0.0152221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_306_96#_c_953_n 0.0279252f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.165
cc_52 VNB N_A_306_96#_c_954_n 0.0621263f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_53 VNB N_A_306_96#_c_955_n 0.0171286f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_54 VNB N_A_306_96#_c_956_n 0.0226279f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.035
cc_55 VNB N_A_306_96#_c_957_n 0.0014655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_306_96#_M1016_g 0.0517191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_306_96#_c_959_n 0.0125997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_306_96#_c_960_n 0.00793516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_306_96#_c_961_n 0.00308834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_306_96#_c_962_n 5.17386e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1518_203#_M1014_g 0.0207732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1518_203#_c_1142_n 0.0156636f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.165
cc_63 VNB N_A_1518_203#_c_1143_n 0.0155514f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_64 VNB N_A_1518_203#_c_1144_n 0.0105463f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=2.01
cc_65 VNB N_A_1518_203#_c_1145_n 0.0023345f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.665
cc_66 VNB N_A_1518_203#_c_1146_n 0.00392193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1518_203#_c_1147_n 0.0310153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1518_203#_c_1148_n 0.0124417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1266_74#_M1017_g 0.04091f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_70 VNB N_A_1266_74#_c_1261_n 0.0182931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1266_74#_c_1262_n 0.016718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1266_74#_c_1263_n 0.0126324f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_73 VNB N_A_1266_74#_c_1264_n 0.0232568f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=2.01
cc_74 VNB N_A_1266_74#_c_1265_n 0.0100399f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.165
cc_75 VNB N_A_1266_74#_c_1266_n 0.0210614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1266_74#_c_1267_n 0.0123873f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.665
cc_77 VNB N_A_1266_74#_c_1268_n 0.00445288f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.845
cc_78 VNB N_A_1266_74#_c_1269_n 0.00403288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1266_74#_c_1270_n 0.00637997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1266_74#_c_1271_n 0.00599516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1266_74#_c_1272_n 0.00266453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1266_74#_c_1273_n 0.00109446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1864_409#_M1002_g 0.0383367f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_84 VNB N_A_1864_409#_c_1422_n 0.0564146f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_85 VNB N_A_1864_409#_c_1423_n 0.0212559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1864_409#_c_1424_n 0.014962f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.845
cc_87 VNB N_A_1864_409#_c_1425_n 0.00445066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VPWR_c_1475_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_30_78#_c_1624_n 0.003401f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_90 VNB N_A_30_78#_c_1625_n 0.00542054f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_91 VNB N_A_30_78#_c_1626_n 9.45585e-19 $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.295
cc_92 VNB N_A_30_78#_c_1627_n 0.00327425f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.845
cc_93 VNB N_A_30_78#_c_1628_n 0.0223919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_30_78#_c_1629_n 0.00159616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_30_78#_c_1630_n 0.00594002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_Q_c_1761_n 0.00811762f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_97 VNB N_Q_c_1762_n 0.00208381f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_98 VNB N_Q_c_1763_n 0.00535471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1791_n 0.0119629f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1
cc_100 VNB N_VGND_c_1792_n 0.0116406f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=2.01
cc_101 VNB N_VGND_c_1793_n 0.0111809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1794_n 0.0145996f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.035
cc_103 VNB N_VGND_c_1795_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1796_n 0.0505973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1797_n 0.0297253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1798_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1799_n 0.019672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1800_n 0.0769928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1801_n 0.0580863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1802_n 0.0325483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1803_n 0.0345892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1804_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1805_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1806_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1807_n 0.588959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VPB N_D_c_238_n 0.0142152f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.828
cc_117 VPB N_D_c_243_n 0.0278711f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.375
cc_118 VPB N_D_c_244_n 0.0265124f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.465
cc_119 VPB N_D_c_241_n 0.0243342f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_120 VPB N_D_c_246_n 0.0207718f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_121 VPB N_CLK_M1006_g 0.0222472f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.01
cc_122 VPB CLK 0.00475607f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_123 VPB N_CLK_c_274_n 0.0119254f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_490_390#_c_321_n 0.0261847f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_125 VPB N_A_490_390#_c_343_n 0.00830698f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_126 VPB N_A_490_390#_c_322_n 0.00918328f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_127 VPB N_A_490_390#_c_323_n 0.00501058f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_128 VPB N_A_490_390#_c_346_n 0.0624804f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_129 VPB N_A_490_390#_c_347_n 0.0191437f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.165
cc_130 VPB N_A_490_390#_c_333_n 0.00559228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_490_390#_c_335_n 0.0078646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_830_359#_c_527_n 0.0637681f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_133 VPB N_A_830_359#_M1012_g 0.00734817f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_134 VPB N_A_830_359#_c_524_n 0.0022958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_830_359#_c_530_n 0.00215186f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=2.01
cc_136 VPB N_A_830_359#_c_526_n 0.00382281f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.845
cc_137 VPB N_RESET_B_c_607_n 0.0208628f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_138 VPB N_RESET_B_c_617_n 0.0166267f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_139 VPB N_RESET_B_c_618_n 0.0169713f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.165
cc_140 VPB N_RESET_B_c_611_n 0.00904598f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_141 VPB N_RESET_B_M1028_g 0.0151047f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=2.01
cc_142 VPB N_RESET_B_c_621_n 0.0572287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_RESET_B_c_622_n 0.0237358f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.665
cc_144 VPB N_RESET_B_c_623_n 0.0192441f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_RESET_B_c_624_n 0.00371129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_RESET_B_c_625_n 0.0198788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_RESET_B_c_626_n 0.00169127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_RESET_B_c_627_n 0.00495528f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_RESET_B_c_628_n 0.00335799f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_RESET_B_c_615_n 9.70225e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_RESET_B_c_630_n 0.0305069f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_RESET_B_c_631_n 0.0539371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_RESET_B_c_632_n 0.00620787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_695_457#_c_833_n 0.0172536f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_155 VPB N_A_695_457#_c_827_n 0.00892422f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_156 VPB N_A_695_457#_c_828_n 0.00538964f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.165
cc_157 VPB N_A_695_457#_c_831_n 0.0241647f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.665
cc_158 VPB N_A_695_457#_c_837_n 0.00256103f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_695_457#_c_838_n 0.00288386f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_695_457#_c_839_n 0.00198824f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_306_96#_M1011_g 0.019846f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_162 VPB N_A_306_96#_c_964_n 0.075647f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_306_96#_c_965_n 0.0561094f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_306_96#_c_966_n 0.0125211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_306_96#_c_954_n 0.0140691f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_166 VPB N_A_306_96#_M1019_g 0.0389765f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=2.01
cc_167 VPB N_A_306_96#_c_969_n 0.179344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_306_96#_M1015_g 0.0110598f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.845
cc_169 VPB N_A_306_96#_c_956_n 0.0299618f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=2.035
cc_170 VPB N_A_306_96#_c_957_n 0.012343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_306_96#_c_973_n 0.00749069f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_306_96#_c_974_n 0.0254973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_306_96#_c_960_n 0.00485186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_306_96#_c_976_n 0.00744406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_1518_203#_c_1149_n 0.0069195f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_176 VPB N_A_1518_203#_c_1150_n 0.0240163f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_177 VPB N_A_1518_203#_c_1151_n 0.0216466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_1518_203#_c_1142_n 0.0041544f $X=-0.19 $Y=1.66 $X2=0.402
+ $Y2=1.165
cc_179 VPB N_A_1518_203#_c_1153_n 0.00705277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_1518_203#_c_1154_n 0.00198797f $X=-0.19 $Y=1.66 $X2=0.32
+ $Y2=1.295
cc_181 VPB N_A_1518_203#_c_1145_n 0.00168296f $X=-0.19 $Y=1.66 $X2=0.32
+ $Y2=1.665
cc_182 VPB N_A_1518_203#_c_1156_n 0.00942442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_1518_203#_c_1157_n 0.00312494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1266_74#_c_1274_n 0.0330758f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_185 VPB N_A_1266_74#_c_1275_n 0.0210347f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_186 VPB N_A_1266_74#_c_1261_n 0.00533618f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_1266_74#_c_1262_n 0.003846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_1266_74#_c_1278_n 0.0108549f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1
cc_189 VPB N_A_1266_74#_c_1279_n 0.022831f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_190 VPB N_A_1266_74#_c_1267_n 9.60226e-19 $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.665
cc_191 VPB N_A_1266_74#_c_1281_n 0.00279628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_1266_74#_c_1282_n 0.00553847f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_1266_74#_c_1270_n 0.00921317f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1266_74#_c_1272_n 2.00274e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_1266_74#_c_1273_n 9.16426e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_1864_409#_c_1426_n 0.0221503f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_197 VPB N_A_1864_409#_c_1422_n 0.0304841f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_198 VPB N_A_1864_409#_c_1423_n 0.00967318f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1864_409#_c_1429_n 0.00988755f $X=-0.19 $Y=1.66 $X2=0.402
+ $Y2=1.165
cc_200 VPB N_A_1864_409#_c_1425_n 0.00279207f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1476_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=2.01
cc_202 VPB N_VPWR_c_1477_n 0.0314475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1478_n 0.00881664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1479_n 0.00367595f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1480_n 0.0150154f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1481_n 0.0203282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1482_n 0.0249158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1483_n 0.019026f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1484_n 0.0204007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1485_n 0.0144553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1486_n 0.0120152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1487_n 0.0660664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1488_n 0.0174851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1489_n 0.0191861f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1490_n 0.056798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1491_n 0.0543442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1492_n 0.0380491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1493_n 0.00613227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1494_n 0.00613824f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1495_n 0.00436844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1496_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1497_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1498_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1475_n 0.11399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_30_78#_c_1631_n 0.00218276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_30_78#_c_1625_n 0.00572962f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_227 VPB N_A_30_78#_c_1633_n 0.0117463f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1
cc_228 VPB N_A_30_78#_c_1634_n 2.77842e-19 $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_229 VPB N_A_30_78#_c_1635_n 0.00299175f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=2.01
cc_230 VPB N_A_30_78#_c_1636_n 0.00146209f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_30_78#_c_1627_n 0.00691983f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.845
cc_232 VPB N_A_30_78#_c_1638_n 0.00633757f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_30_78#_c_1639_n 0.00843421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB Q 0.0106664f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_235 VPB Q 0.0225117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_Q_c_1763_n 0.00313086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 N_D_M1020_g N_RESET_B_M1008_g 0.0245154f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_238 N_D_c_241_n N_RESET_B_M1008_g 9.92331e-19 $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_239 N_D_c_238_n N_RESET_B_c_607_n 0.0245154f $X=0.402 $Y=1.828 $X2=0 $Y2=0
cc_240 N_D_c_243_n N_RESET_B_c_617_n 0.00650355f $X=0.495 $Y=2.375 $X2=0 $Y2=0
cc_241 N_D_c_244_n N_RESET_B_c_622_n 0.016022f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_242 N_D_c_240_n N_RESET_B_c_614_n 0.0245154f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_243 N_D_c_246_n N_RESET_B_c_630_n 0.0245154f $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_244 N_D_c_244_n N_VPWR_c_1477_n 0.00596f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_245 N_D_c_241_n N_VPWR_c_1477_n 0.0129077f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_246 N_D_c_246_n N_VPWR_c_1477_n 7.18884e-19 $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_247 N_D_c_244_n N_VPWR_c_1478_n 4.24767e-19 $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_248 N_D_c_244_n N_VPWR_c_1488_n 0.00445602f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_249 N_D_c_244_n N_VPWR_c_1475_n 0.00898825f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_250 N_D_M1020_g N_A_30_78#_c_1624_n 0.0108589f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_251 N_D_c_241_n N_A_30_78#_c_1624_n 0.00411346f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_252 N_D_c_244_n N_A_30_78#_c_1631_n 0.00411415f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_253 N_D_M1020_g N_A_30_78#_c_1625_n 0.0145237f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_254 N_D_c_241_n N_A_30_78#_c_1625_n 0.0884076f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_255 N_D_M1020_g N_A_30_78#_c_1628_n 0.00806237f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_256 N_D_c_240_n N_A_30_78#_c_1628_n 0.00161806f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_257 N_D_c_241_n N_A_30_78#_c_1628_n 0.0286676f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_258 N_D_c_243_n N_A_30_78#_c_1638_n 0.00464415f $X=0.495 $Y=2.375 $X2=0 $Y2=0
cc_259 N_D_c_244_n N_A_30_78#_c_1638_n 0.00480701f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_260 N_D_M1020_g N_VGND_c_1791_n 0.00190636f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_261 N_D_M1020_g N_VGND_c_1797_n 0.00429844f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_262 N_D_M1020_g N_VGND_c_1807_n 0.00539454f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_263 N_CLK_M1006_g N_A_490_390#_c_335_n 0.00117088f $X=1.925 $Y=2.45 $X2=0
+ $Y2=0
cc_264 CLK N_A_490_390#_c_335_n 0.00246327f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_265 N_CLK_M1006_g N_RESET_B_c_607_n 0.00513392f $X=1.925 $Y=2.45 $X2=0 $Y2=0
cc_266 N_CLK_c_274_n N_RESET_B_c_607_n 0.00753785f $X=1.91 $Y=1.61 $X2=0 $Y2=0
cc_267 N_CLK_c_275_n N_RESET_B_c_608_n 0.0104164f $X=1.91 $Y=1.435 $X2=0 $Y2=0
cc_268 N_CLK_M1006_g N_RESET_B_c_623_n 0.00374052f $X=1.925 $Y=2.45 $X2=0 $Y2=0
cc_269 CLK N_RESET_B_c_623_n 0.0129811f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_270 N_CLK_c_275_n N_RESET_B_c_614_n 0.00429864f $X=1.91 $Y=1.435 $X2=0 $Y2=0
cc_271 N_CLK_M1006_g N_RESET_B_c_615_n 2.69506e-19 $X=1.925 $Y=2.45 $X2=0 $Y2=0
cc_272 CLK N_A_306_96#_M1030_s 4.93455e-19 $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_273 N_CLK_M1006_g N_A_306_96#_M1011_g 0.042279f $X=1.925 $Y=2.45 $X2=0 $Y2=0
cc_274 CLK N_A_306_96#_c_952_n 7.59256e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_275 N_CLK_c_275_n N_A_306_96#_c_952_n 0.0246727f $X=1.91 $Y=1.435 $X2=0 $Y2=0
cc_276 CLK N_A_306_96#_c_954_n 0.00402032f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_277 N_CLK_c_274_n N_A_306_96#_c_954_n 0.0202235f $X=1.91 $Y=1.61 $X2=0 $Y2=0
cc_278 N_CLK_c_275_n N_A_306_96#_c_954_n 0.00111896f $X=1.91 $Y=1.435 $X2=0
+ $Y2=0
cc_279 N_CLK_c_275_n N_A_306_96#_c_959_n 0.00654248f $X=1.91 $Y=1.435 $X2=0
+ $Y2=0
cc_280 N_CLK_M1006_g N_A_306_96#_c_960_n 0.00252075f $X=1.925 $Y=2.45 $X2=0
+ $Y2=0
cc_281 CLK N_A_306_96#_c_960_n 0.0368206f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_282 N_CLK_c_274_n N_A_306_96#_c_960_n 0.00297206f $X=1.91 $Y=1.61 $X2=0 $Y2=0
cc_283 N_CLK_c_275_n N_A_306_96#_c_960_n 0.00292393f $X=1.91 $Y=1.435 $X2=0
+ $Y2=0
cc_284 CLK N_A_306_96#_c_989_n 0.0262776f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_285 N_CLK_c_275_n N_A_306_96#_c_989_n 0.0131294f $X=1.91 $Y=1.435 $X2=0 $Y2=0
cc_286 CLK N_A_306_96#_c_961_n 0.00201688f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_287 N_CLK_c_274_n N_A_306_96#_c_961_n 0.00215961f $X=1.91 $Y=1.61 $X2=0 $Y2=0
cc_288 N_CLK_M1006_g N_A_306_96#_c_976_n 0.00437328f $X=1.925 $Y=2.45 $X2=0
+ $Y2=0
cc_289 CLK N_A_306_96#_c_976_n 0.00507476f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_290 N_CLK_c_274_n N_A_306_96#_c_976_n 0.00240115f $X=1.91 $Y=1.61 $X2=0 $Y2=0
cc_291 CLK N_A_306_96#_c_962_n 0.0311526f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_292 N_CLK_c_275_n N_A_306_96#_c_962_n 0.00104584f $X=1.91 $Y=1.435 $X2=0
+ $Y2=0
cc_293 N_CLK_M1006_g N_VPWR_c_1478_n 0.00566599f $X=1.925 $Y=2.45 $X2=0 $Y2=0
cc_294 N_CLK_M1006_g N_VPWR_c_1479_n 0.00947197f $X=1.925 $Y=2.45 $X2=0 $Y2=0
cc_295 N_CLK_M1006_g N_VPWR_c_1489_n 0.00403581f $X=1.925 $Y=2.45 $X2=0 $Y2=0
cc_296 N_CLK_M1006_g N_VPWR_c_1475_n 0.00492022f $X=1.925 $Y=2.45 $X2=0 $Y2=0
cc_297 N_CLK_M1006_g N_A_30_78#_c_1633_n 0.00265624f $X=1.925 $Y=2.45 $X2=0
+ $Y2=0
cc_298 N_CLK_M1006_g N_A_30_78#_c_1634_n 0.0107512f $X=1.925 $Y=2.45 $X2=0 $Y2=0
cc_299 CLK N_A_30_78#_c_1634_n 6.22319e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_300 N_CLK_M1006_g N_A_30_78#_c_1635_n 0.00727501f $X=1.925 $Y=2.45 $X2=0
+ $Y2=0
cc_301 CLK N_A_30_78#_c_1635_n 0.0038074f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_302 CLK N_VGND_M1030_d 0.00233115f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_303 N_CLK_c_275_n N_VGND_c_1792_n 0.00254438f $X=1.91 $Y=1.435 $X2=0 $Y2=0
cc_304 N_CLK_c_275_n N_VGND_c_1807_n 9.39239e-19 $X=1.91 $Y=1.435 $X2=0 $Y2=0
cc_305 N_A_490_390#_c_330_n N_A_830_359#_M1026_d 0.00330812f $X=5.48 $Y=0.65
+ $X2=-0.19 $Y2=-0.245
cc_306 N_A_490_390#_c_353_p N_A_830_359#_M1026_d 0.00218198f $X=5.565 $Y=0.565
+ $X2=-0.19 $Y2=-0.245
cc_307 N_A_490_390#_c_331_n N_A_830_359#_M1026_d 0.00764003f $X=7.25 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_308 N_A_490_390#_c_321_n N_A_830_359#_c_527_n 0.00467059f $X=3.412 $Y=1.985
+ $X2=0 $Y2=0
cc_309 N_A_490_390#_c_323_n N_A_830_359#_M1012_g 0.00466042f $X=4.005 $Y=1.405
+ $X2=0 $Y2=0
cc_310 N_A_490_390#_M1027_g N_A_830_359#_M1012_g 0.0529911f $X=4.005 $Y=0.9
+ $X2=0 $Y2=0
cc_311 N_A_490_390#_c_330_n N_A_830_359#_M1012_g 0.00341287f $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_312 N_A_490_390#_c_339_n N_A_830_359#_M1012_g 0.00599849f $X=4.355 $Y=0.415
+ $X2=0 $Y2=0
cc_313 N_A_490_390#_c_323_n N_A_830_359#_c_524_n 3.61909e-19 $X=4.005 $Y=1.405
+ $X2=0 $Y2=0
cc_314 N_A_490_390#_M1027_g N_A_830_359#_c_524_n 0.00131686f $X=4.005 $Y=0.9
+ $X2=0 $Y2=0
cc_315 N_A_490_390#_c_330_n N_A_830_359#_c_542_n 0.0658997f $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_316 N_A_490_390#_c_331_n N_A_830_359#_c_542_n 0.00571426f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_317 N_A_490_390#_c_330_n N_A_830_359#_c_544_n 3.80876e-19 $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_318 N_A_490_390#_c_339_n N_A_830_359#_c_544_n 0.00969153f $X=4.355 $Y=0.415
+ $X2=0 $Y2=0
cc_319 N_A_490_390#_c_327_n N_A_830_359#_c_530_n 0.00388841f $X=6.33 $Y=1.27
+ $X2=0 $Y2=0
cc_320 N_A_490_390#_c_325_n N_A_830_359#_c_525_n 0.00184952f $X=6.255 $Y=1.195
+ $X2=0 $Y2=0
cc_321 N_A_490_390#_c_330_n N_A_830_359#_c_525_n 0.00596144f $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_322 N_A_490_390#_c_331_n N_A_830_359#_c_525_n 0.0168368f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_323 N_A_490_390#_c_327_n N_A_830_359#_c_526_n 0.00184952f $X=6.33 $Y=1.27
+ $X2=0 $Y2=0
cc_324 N_A_490_390#_M1027_g N_RESET_B_c_608_n 0.00526413f $X=4.005 $Y=0.9 $X2=0
+ $Y2=0
cc_325 N_A_490_390#_c_329_n N_RESET_B_c_608_n 0.0234047f $X=4.27 $Y=0.415 $X2=0
+ $Y2=0
cc_326 N_A_490_390#_c_330_n N_RESET_B_c_608_n 0.0029296f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_327 N_A_490_390#_c_336_n N_RESET_B_c_608_n 0.0109521f $X=2.797 $Y=0.415 $X2=0
+ $Y2=0
cc_328 N_A_490_390#_c_339_n N_RESET_B_c_608_n 0.00219835f $X=4.355 $Y=0.415
+ $X2=0 $Y2=0
cc_329 N_A_490_390#_c_330_n N_RESET_B_M1004_g 0.0122094f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_330 N_A_490_390#_c_353_p N_RESET_B_M1004_g 6.19914e-19 $X=5.565 $Y=0.565
+ $X2=0 $Y2=0
cc_331 N_A_490_390#_c_339_n N_RESET_B_M1004_g 0.00649083f $X=4.355 $Y=0.415
+ $X2=0 $Y2=0
cc_332 N_A_490_390#_c_321_n N_RESET_B_c_623_n 0.00282958f $X=3.412 $Y=1.985
+ $X2=0 $Y2=0
cc_333 N_A_490_390#_c_343_n N_RESET_B_c_623_n 0.00383268f $X=3.412 $Y=2.123
+ $X2=0 $Y2=0
cc_334 N_A_490_390#_c_322_n N_RESET_B_c_623_n 0.00429293f $X=3.79 $Y=1.635 $X2=0
+ $Y2=0
cc_335 N_A_490_390#_c_335_n N_RESET_B_c_623_n 0.0452109f $X=3.03 $Y=1.882 $X2=0
+ $Y2=0
cc_336 N_A_490_390#_c_338_n N_RESET_B_c_623_n 5.22657e-19 $X=2.99 $Y=1.345 $X2=0
+ $Y2=0
cc_337 N_A_490_390#_c_346_n N_RESET_B_c_625_n 0.00268688f $X=7.265 $Y=2.39 $X2=0
+ $Y2=0
cc_338 N_A_490_390#_c_333_n N_RESET_B_c_625_n 0.0220527f $X=7.13 $Y=2.14 $X2=0
+ $Y2=0
cc_339 N_A_490_390#_c_325_n N_A_695_457#_M1026_g 0.00895705f $X=6.255 $Y=1.195
+ $X2=0 $Y2=0
cc_340 N_A_490_390#_c_330_n N_A_695_457#_M1026_g 0.0118282f $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_341 N_A_490_390#_c_353_p N_A_695_457#_M1026_g 0.0047339f $X=5.565 $Y=0.565
+ $X2=0 $Y2=0
cc_342 N_A_490_390#_c_332_n N_A_695_457#_M1026_g 0.00591041f $X=5.65 $Y=0.34
+ $X2=0 $Y2=0
cc_343 N_A_490_390#_c_323_n N_A_695_457#_c_827_n 0.0112879f $X=4.005 $Y=1.405
+ $X2=0 $Y2=0
cc_344 N_A_490_390#_M1027_g N_A_695_457#_c_827_n 0.00941138f $X=4.005 $Y=0.9
+ $X2=0 $Y2=0
cc_345 N_A_490_390#_c_347_n N_A_695_457#_c_827_n 5.3662e-19 $X=3.412 $Y=2.21
+ $X2=0 $Y2=0
cc_346 N_A_490_390#_c_327_n N_A_695_457#_c_831_n 0.00170129f $X=6.33 $Y=1.27
+ $X2=0 $Y2=0
cc_347 N_A_490_390#_c_322_n N_A_695_457#_c_832_n 7.94787e-19 $X=3.79 $Y=1.635
+ $X2=0 $Y2=0
cc_348 N_A_490_390#_c_323_n N_A_695_457#_c_832_n 0.00370718f $X=4.005 $Y=1.405
+ $X2=0 $Y2=0
cc_349 N_A_490_390#_M1027_g N_A_695_457#_c_832_n 0.00808934f $X=4.005 $Y=0.9
+ $X2=0 $Y2=0
cc_350 N_A_490_390#_c_329_n N_A_695_457#_c_832_n 0.0356492f $X=4.27 $Y=0.415
+ $X2=0 $Y2=0
cc_351 N_A_490_390#_c_339_n N_A_695_457#_c_832_n 0.00147569f $X=4.355 $Y=0.415
+ $X2=0 $Y2=0
cc_352 N_A_490_390#_c_347_n N_A_695_457#_c_838_n 0.00280663f $X=3.412 $Y=2.21
+ $X2=0 $Y2=0
cc_353 N_A_490_390#_c_335_n N_A_306_96#_M1011_g 0.00691852f $X=3.03 $Y=1.882
+ $X2=0 $Y2=0
cc_354 N_A_490_390#_c_336_n N_A_306_96#_c_952_n 0.00644381f $X=2.797 $Y=0.415
+ $X2=0 $Y2=0
cc_355 N_A_490_390#_c_337_n N_A_306_96#_c_952_n 0.00500076f $X=2.99 $Y=1.195
+ $X2=0 $Y2=0
cc_356 N_A_490_390#_c_343_n N_A_306_96#_c_964_n 0.0205243f $X=3.412 $Y=2.123
+ $X2=0 $Y2=0
cc_357 N_A_490_390#_c_335_n N_A_306_96#_c_964_n 0.0188445f $X=3.03 $Y=1.882
+ $X2=0 $Y2=0
cc_358 N_A_490_390#_c_347_n N_A_306_96#_c_965_n 0.00899647f $X=3.412 $Y=2.21
+ $X2=0 $Y2=0
cc_359 N_A_490_390#_c_321_n N_A_306_96#_c_953_n 0.0231012f $X=3.412 $Y=1.985
+ $X2=0 $Y2=0
cc_360 N_A_490_390#_c_328_n N_A_306_96#_c_953_n 4.22569e-19 $X=3.03 $Y=1.56
+ $X2=0 $Y2=0
cc_361 N_A_490_390#_c_335_n N_A_306_96#_c_953_n 0.00382077f $X=3.03 $Y=1.882
+ $X2=0 $Y2=0
cc_362 N_A_490_390#_c_338_n N_A_306_96#_c_953_n 0.00249449f $X=2.99 $Y=1.345
+ $X2=0 $Y2=0
cc_363 N_A_490_390#_c_321_n N_A_306_96#_c_954_n 0.0249553f $X=3.412 $Y=1.985
+ $X2=0 $Y2=0
cc_364 N_A_490_390#_c_323_n N_A_306_96#_c_954_n 7.47803e-19 $X=4.005 $Y=1.405
+ $X2=0 $Y2=0
cc_365 N_A_490_390#_c_328_n N_A_306_96#_c_954_n 0.0105491f $X=3.03 $Y=1.56 $X2=0
+ $Y2=0
cc_366 N_A_490_390#_c_335_n N_A_306_96#_c_954_n 0.0119493f $X=3.03 $Y=1.882
+ $X2=0 $Y2=0
cc_367 N_A_490_390#_c_336_n N_A_306_96#_c_954_n 0.00526481f $X=2.797 $Y=0.415
+ $X2=0 $Y2=0
cc_368 N_A_490_390#_c_338_n N_A_306_96#_c_954_n 0.00910693f $X=2.99 $Y=1.345
+ $X2=0 $Y2=0
cc_369 N_A_490_390#_M1027_g N_A_306_96#_c_955_n 0.0182908f $X=4.005 $Y=0.9 $X2=0
+ $Y2=0
cc_370 N_A_490_390#_c_329_n N_A_306_96#_c_955_n 0.00349197f $X=4.27 $Y=0.415
+ $X2=0 $Y2=0
cc_371 N_A_490_390#_c_336_n N_A_306_96#_c_955_n 0.00465637f $X=2.797 $Y=0.415
+ $X2=0 $Y2=0
cc_372 N_A_490_390#_c_322_n N_A_306_96#_M1019_g 0.00459329f $X=3.79 $Y=1.635
+ $X2=0 $Y2=0
cc_373 N_A_490_390#_c_347_n N_A_306_96#_M1019_g 0.0147557f $X=3.412 $Y=2.21
+ $X2=0 $Y2=0
cc_374 N_A_490_390#_c_346_n N_A_306_96#_M1015_g 0.00735807f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_375 N_A_490_390#_c_326_n N_A_306_96#_c_956_n 0.0196234f $X=6.69 $Y=1.27 $X2=0
+ $Y2=0
cc_376 N_A_490_390#_c_346_n N_A_306_96#_c_956_n 0.0220783f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_377 N_A_490_390#_c_333_n N_A_306_96#_c_956_n 0.0164562f $X=7.13 $Y=2.14 $X2=0
+ $Y2=0
cc_378 N_A_490_390#_c_341_n N_A_306_96#_c_956_n 0.00266664f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_379 N_A_490_390#_c_327_n N_A_306_96#_c_957_n 0.0196234f $X=6.33 $Y=1.27 $X2=0
+ $Y2=0
cc_380 N_A_490_390#_c_331_n N_A_306_96#_M1016_g 0.0088085f $X=7.25 $Y=0.34 $X2=0
+ $Y2=0
cc_381 N_A_490_390#_c_333_n N_A_306_96#_M1016_g 0.00923892f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_382 N_A_490_390#_c_334_n N_A_306_96#_M1016_g 0.0233298f $X=7.335 $Y=1.015
+ $X2=0 $Y2=0
cc_383 N_A_490_390#_c_340_n N_A_306_96#_M1016_g 0.0213806f $X=6.855 $Y=1.18
+ $X2=0 $Y2=0
cc_384 N_A_490_390#_c_341_n N_A_306_96#_M1016_g 0.011895f $X=7.335 $Y=1.18 $X2=0
+ $Y2=0
cc_385 N_A_490_390#_c_346_n N_A_306_96#_c_974_n 0.00118457f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_386 N_A_490_390#_M1025_d N_A_306_96#_c_989_n 0.00252881f $X=2.575 $Y=0.595
+ $X2=0 $Y2=0
cc_387 N_A_490_390#_c_336_n N_A_306_96#_c_989_n 0.00667592f $X=2.797 $Y=0.415
+ $X2=0 $Y2=0
cc_388 N_A_490_390#_c_337_n N_A_306_96#_c_989_n 0.0136439f $X=2.99 $Y=1.195
+ $X2=0 $Y2=0
cc_389 N_A_490_390#_c_335_n N_A_306_96#_c_976_n 0.00494199f $X=3.03 $Y=1.882
+ $X2=0 $Y2=0
cc_390 N_A_490_390#_c_328_n N_A_306_96#_c_1035_n 0.00496499f $X=3.03 $Y=1.56
+ $X2=0 $Y2=0
cc_391 N_A_490_390#_c_335_n N_A_306_96#_c_1035_n 0.0357325f $X=3.03 $Y=1.882
+ $X2=0 $Y2=0
cc_392 N_A_490_390#_M1025_d N_A_306_96#_c_962_n 0.00180532f $X=2.575 $Y=0.595
+ $X2=0 $Y2=0
cc_393 N_A_490_390#_c_328_n N_A_306_96#_c_962_n 0.00765569f $X=3.03 $Y=1.56
+ $X2=0 $Y2=0
cc_394 N_A_490_390#_c_337_n N_A_306_96#_c_962_n 0.0156102f $X=2.99 $Y=1.195
+ $X2=0 $Y2=0
cc_395 N_A_490_390#_c_346_n N_A_1518_203#_c_1150_n 0.0222944f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_396 N_A_490_390#_c_333_n N_A_1518_203#_c_1150_n 3.6309e-19 $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_397 N_A_490_390#_c_346_n N_A_1518_203#_c_1151_n 0.029186f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_398 N_A_490_390#_c_331_n N_A_1518_203#_M1014_g 0.00107872f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_399 N_A_490_390#_c_334_n N_A_1518_203#_M1014_g 0.0045389f $X=7.335 $Y=1.015
+ $X2=0 $Y2=0
cc_400 N_A_490_390#_c_333_n N_A_1518_203#_c_1142_n 0.00240511f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_401 N_A_490_390#_c_341_n N_A_1518_203#_c_1146_n 0.0276613f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_402 N_A_490_390#_c_341_n N_A_1518_203#_c_1147_n 0.00201148f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_403 N_A_490_390#_c_331_n N_A_1266_74#_M1022_d 0.00949775f $X=7.25 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_404 N_A_490_390#_c_325_n N_A_1266_74#_c_1287_n 0.0033591f $X=6.255 $Y=1.195
+ $X2=0 $Y2=0
cc_405 N_A_490_390#_c_330_n N_A_1266_74#_c_1287_n 0.00205017f $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_406 N_A_490_390#_c_331_n N_A_1266_74#_c_1287_n 0.00851496f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_407 N_A_490_390#_c_325_n N_A_1266_74#_c_1268_n 0.00750067f $X=6.255 $Y=1.195
+ $X2=0 $Y2=0
cc_408 N_A_490_390#_c_326_n N_A_1266_74#_c_1268_n 0.00921579f $X=6.69 $Y=1.27
+ $X2=0 $Y2=0
cc_409 N_A_490_390#_c_327_n N_A_1266_74#_c_1268_n 0.00149703f $X=6.33 $Y=1.27
+ $X2=0 $Y2=0
cc_410 N_A_490_390#_c_333_n N_A_1266_74#_c_1268_n 0.00662434f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_411 N_A_490_390#_c_340_n N_A_1266_74#_c_1268_n 6.18001e-19 $X=6.855 $Y=1.18
+ $X2=0 $Y2=0
cc_412 N_A_490_390#_c_341_n N_A_1266_74#_c_1268_n 0.0224751f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_413 N_A_490_390#_c_346_n N_A_1266_74#_c_1281_n 0.00556629f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_414 N_A_490_390#_c_333_n N_A_1266_74#_c_1281_n 0.0279379f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_415 N_A_490_390#_c_326_n N_A_1266_74#_c_1269_n 0.00430336f $X=6.69 $Y=1.27
+ $X2=0 $Y2=0
cc_416 N_A_490_390#_c_331_n N_A_1266_74#_c_1269_n 0.0414158f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_417 N_A_490_390#_c_334_n N_A_1266_74#_c_1269_n 0.0196081f $X=7.335 $Y=1.015
+ $X2=0 $Y2=0
cc_418 N_A_490_390#_c_340_n N_A_1266_74#_c_1269_n 0.00746605f $X=6.855 $Y=1.18
+ $X2=0 $Y2=0
cc_419 N_A_490_390#_c_341_n N_A_1266_74#_c_1269_n 0.030444f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_420 N_A_490_390#_c_346_n N_A_1266_74#_c_1303_n 0.0145082f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_421 N_A_490_390#_c_333_n N_A_1266_74#_c_1303_n 0.0232672f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_422 N_A_490_390#_c_346_n N_A_1266_74#_c_1282_n 0.00566122f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_423 N_A_490_390#_c_333_n N_A_1266_74#_c_1282_n 0.0462528f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_424 N_A_490_390#_c_333_n N_A_1266_74#_c_1271_n 0.0142973f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_425 N_A_490_390#_c_326_n N_A_1266_74#_c_1272_n 0.0016242f $X=6.69 $Y=1.27
+ $X2=0 $Y2=0
cc_426 N_A_490_390#_c_333_n N_A_1266_74#_c_1272_n 0.00830682f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_427 N_A_490_390#_c_346_n N_VPWR_c_1491_n 0.00391396f $X=7.265 $Y=2.39 $X2=0
+ $Y2=0
cc_428 N_A_490_390#_c_346_n N_VPWR_c_1475_n 0.0052212f $X=7.265 $Y=2.39 $X2=0
+ $Y2=0
cc_429 N_A_490_390#_c_347_n N_VPWR_c_1475_n 9.49986e-19 $X=3.412 $Y=2.21 $X2=0
+ $Y2=0
cc_430 N_A_490_390#_M1011_d N_A_30_78#_c_1635_n 0.00666319f $X=2.45 $Y=1.95
+ $X2=0 $Y2=0
cc_431 N_A_490_390#_c_335_n N_A_30_78#_c_1635_n 0.0265502f $X=3.03 $Y=1.882
+ $X2=0 $Y2=0
cc_432 N_A_490_390#_M1027_g N_A_30_78#_c_1626_n 4.91816e-19 $X=4.005 $Y=0.9
+ $X2=0 $Y2=0
cc_433 N_A_490_390#_c_337_n N_A_30_78#_c_1626_n 0.00848291f $X=2.99 $Y=1.195
+ $X2=0 $Y2=0
cc_434 N_A_490_390#_c_338_n N_A_30_78#_c_1626_n 0.00178482f $X=2.99 $Y=1.345
+ $X2=0 $Y2=0
cc_435 N_A_490_390#_c_322_n N_A_30_78#_c_1636_n 0.00228024f $X=3.79 $Y=1.635
+ $X2=0 $Y2=0
cc_436 N_A_490_390#_c_347_n N_A_30_78#_c_1636_n 0.0120307f $X=3.412 $Y=2.21
+ $X2=0 $Y2=0
cc_437 N_A_490_390#_c_335_n N_A_30_78#_c_1636_n 0.00502749f $X=3.03 $Y=1.882
+ $X2=0 $Y2=0
cc_438 N_A_490_390#_c_321_n N_A_30_78#_c_1627_n 0.00782591f $X=3.412 $Y=1.985
+ $X2=0 $Y2=0
cc_439 N_A_490_390#_c_322_n N_A_30_78#_c_1627_n 0.0132482f $X=3.79 $Y=1.635
+ $X2=0 $Y2=0
cc_440 N_A_490_390#_c_323_n N_A_30_78#_c_1627_n 0.00301777f $X=4.005 $Y=1.405
+ $X2=0 $Y2=0
cc_441 N_A_490_390#_M1027_g N_A_30_78#_c_1627_n 2.69467e-19 $X=4.005 $Y=0.9
+ $X2=0 $Y2=0
cc_442 N_A_490_390#_c_328_n N_A_30_78#_c_1627_n 0.00627045f $X=3.03 $Y=1.56
+ $X2=0 $Y2=0
cc_443 N_A_490_390#_c_335_n N_A_30_78#_c_1627_n 0.0335712f $X=3.03 $Y=1.882
+ $X2=0 $Y2=0
cc_444 N_A_490_390#_c_321_n N_A_30_78#_c_1639_n 0.0011758f $X=3.412 $Y=1.985
+ $X2=0 $Y2=0
cc_445 N_A_490_390#_c_347_n N_A_30_78#_c_1639_n 0.00336023f $X=3.412 $Y=2.21
+ $X2=0 $Y2=0
cc_446 N_A_490_390#_c_335_n N_A_30_78#_c_1639_n 0.0228903f $X=3.03 $Y=1.882
+ $X2=0 $Y2=0
cc_447 N_A_490_390#_c_329_n N_A_30_78#_c_1629_n 0.0192833f $X=4.27 $Y=0.415
+ $X2=0 $Y2=0
cc_448 N_A_490_390#_c_335_n N_A_30_78#_c_1629_n 0.00300061f $X=3.03 $Y=1.882
+ $X2=0 $Y2=0
cc_449 N_A_490_390#_c_336_n N_A_30_78#_c_1629_n 0.0293939f $X=2.797 $Y=0.415
+ $X2=0 $Y2=0
cc_450 N_A_490_390#_c_321_n N_A_30_78#_c_1630_n 0.00403943f $X=3.412 $Y=1.985
+ $X2=0 $Y2=0
cc_451 N_A_490_390#_c_322_n N_A_30_78#_c_1630_n 8.36337e-19 $X=3.79 $Y=1.635
+ $X2=0 $Y2=0
cc_452 N_A_490_390#_M1027_g N_A_30_78#_c_1630_n 0.0016508f $X=4.005 $Y=0.9 $X2=0
+ $Y2=0
cc_453 N_A_490_390#_c_335_n N_A_30_78#_c_1630_n 0.0101271f $X=3.03 $Y=1.882
+ $X2=0 $Y2=0
cc_454 N_A_490_390#_c_338_n N_A_30_78#_c_1630_n 0.0129594f $X=2.99 $Y=1.345
+ $X2=0 $Y2=0
cc_455 N_A_490_390#_c_330_n N_VGND_M1004_d 0.00922416f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_456 N_A_490_390#_c_336_n N_VGND_c_1792_n 0.0302166f $X=2.797 $Y=0.415 $X2=0
+ $Y2=0
cc_457 N_A_490_390#_c_331_n N_VGND_c_1793_n 0.00831292f $X=7.25 $Y=0.34 $X2=0
+ $Y2=0
cc_458 N_A_490_390#_c_334_n N_VGND_c_1793_n 0.00983536f $X=7.335 $Y=1.015 $X2=0
+ $Y2=0
cc_459 N_A_490_390#_c_329_n N_VGND_c_1800_n 0.0540738f $X=4.27 $Y=0.415 $X2=0
+ $Y2=0
cc_460 N_A_490_390#_c_330_n N_VGND_c_1800_n 0.0389968f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_461 N_A_490_390#_c_332_n N_VGND_c_1800_n 0.0107916f $X=5.65 $Y=0.34 $X2=0
+ $Y2=0
cc_462 N_A_490_390#_c_336_n N_VGND_c_1800_n 0.0225471f $X=2.797 $Y=0.415 $X2=0
+ $Y2=0
cc_463 N_A_490_390#_c_339_n N_VGND_c_1800_n 0.0103964f $X=4.355 $Y=0.415 $X2=0
+ $Y2=0
cc_464 N_A_490_390#_c_325_n N_VGND_c_1801_n 0.00278271f $X=6.255 $Y=1.195 $X2=0
+ $Y2=0
cc_465 N_A_490_390#_c_330_n N_VGND_c_1801_n 0.00286598f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_466 N_A_490_390#_c_331_n N_VGND_c_1801_n 0.114761f $X=7.25 $Y=0.34 $X2=0
+ $Y2=0
cc_467 N_A_490_390#_c_332_n N_VGND_c_1801_n 0.0117553f $X=5.65 $Y=0.34 $X2=0
+ $Y2=0
cc_468 N_A_490_390#_c_325_n N_VGND_c_1807_n 0.00361111f $X=6.255 $Y=1.195 $X2=0
+ $Y2=0
cc_469 N_A_490_390#_c_329_n N_VGND_c_1807_n 0.0393214f $X=4.27 $Y=0.415 $X2=0
+ $Y2=0
cc_470 N_A_490_390#_c_330_n N_VGND_c_1807_n 0.0191089f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_471 N_A_490_390#_c_331_n N_VGND_c_1807_n 0.0660751f $X=7.25 $Y=0.34 $X2=0
+ $Y2=0
cc_472 N_A_490_390#_c_332_n N_VGND_c_1807_n 0.00639038f $X=5.65 $Y=0.34 $X2=0
+ $Y2=0
cc_473 N_A_490_390#_c_336_n N_VGND_c_1807_n 0.0156523f $X=2.797 $Y=0.415 $X2=0
+ $Y2=0
cc_474 N_A_490_390#_c_339_n N_VGND_c_1807_n 0.0055037f $X=4.355 $Y=0.415 $X2=0
+ $Y2=0
cc_475 N_A_490_390#_c_330_n A_894_138# 0.00134267f $X=5.48 $Y=0.65 $X2=-0.19
+ $Y2=-0.245
cc_476 N_A_830_359#_M1012_g N_RESET_B_c_608_n 0.00555255f $X=4.395 $Y=0.9 $X2=0
+ $Y2=0
cc_477 N_A_830_359#_M1012_g N_RESET_B_M1004_g 0.0417175f $X=4.395 $Y=0.9 $X2=0
+ $Y2=0
cc_478 N_A_830_359#_c_524_n N_RESET_B_M1004_g 0.00105981f $X=4.355 $Y=1.96 $X2=0
+ $Y2=0
cc_479 N_A_830_359#_c_542_n N_RESET_B_M1004_g 0.0111445f $X=5.82 $Y=0.99 $X2=0
+ $Y2=0
cc_480 N_A_830_359#_c_527_n N_RESET_B_c_618_n 0.0131923f $X=4.24 $Y=2.21 $X2=0
+ $Y2=0
cc_481 N_A_830_359#_M1012_g N_RESET_B_c_611_n 0.0138167f $X=4.395 $Y=0.9 $X2=0
+ $Y2=0
cc_482 N_A_830_359#_c_524_n N_RESET_B_c_611_n 2.97938e-19 $X=4.355 $Y=1.96 $X2=0
+ $Y2=0
cc_483 N_A_830_359#_c_542_n N_RESET_B_c_613_n 0.00240316f $X=5.82 $Y=0.99 $X2=0
+ $Y2=0
cc_484 N_A_830_359#_c_527_n N_RESET_B_c_623_n 0.0115525f $X=4.24 $Y=2.21 $X2=0
+ $Y2=0
cc_485 N_A_830_359#_c_524_n N_RESET_B_c_623_n 0.0166498f $X=4.355 $Y=1.96 $X2=0
+ $Y2=0
cc_486 N_A_830_359#_M1005_d N_RESET_B_c_625_n 0.00144653f $X=5.955 $Y=1.735
+ $X2=0 $Y2=0
cc_487 N_A_830_359#_c_530_n N_RESET_B_c_625_n 0.0389295f $X=6.145 $Y=2.03 $X2=0
+ $Y2=0
cc_488 N_A_830_359#_c_527_n N_RESET_B_c_631_n 0.0191507f $X=4.24 $Y=2.21 $X2=0
+ $Y2=0
cc_489 N_A_830_359#_c_524_n N_RESET_B_c_631_n 3.38963e-19 $X=4.355 $Y=1.96 $X2=0
+ $Y2=0
cc_490 N_A_830_359#_c_542_n N_A_695_457#_M1026_g 0.0122404f $X=5.82 $Y=0.99
+ $X2=0 $Y2=0
cc_491 N_A_830_359#_c_525_n N_A_695_457#_M1026_g 0.00563857f $X=5.985 $Y=0.855
+ $X2=0 $Y2=0
cc_492 N_A_830_359#_c_526_n N_A_695_457#_M1026_g 0.0019205f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_493 N_A_830_359#_c_526_n N_A_695_457#_c_833_n 0.00373472f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_494 N_A_830_359#_c_527_n N_A_695_457#_c_827_n 0.00709856f $X=4.24 $Y=2.21
+ $X2=0 $Y2=0
cc_495 N_A_830_359#_M1012_g N_A_695_457#_c_827_n 0.00223534f $X=4.395 $Y=0.9
+ $X2=0 $Y2=0
cc_496 N_A_830_359#_c_524_n N_A_695_457#_c_827_n 0.074703f $X=4.355 $Y=1.96
+ $X2=0 $Y2=0
cc_497 N_A_830_359#_c_527_n N_A_695_457#_c_861_n 0.0113183f $X=4.24 $Y=2.21
+ $X2=0 $Y2=0
cc_498 N_A_830_359#_c_524_n N_A_695_457#_c_861_n 0.00697489f $X=4.355 $Y=1.96
+ $X2=0 $Y2=0
cc_499 N_A_830_359#_c_527_n N_A_695_457#_c_828_n 0.00375838f $X=4.24 $Y=2.21
+ $X2=0 $Y2=0
cc_500 N_A_830_359#_M1012_g N_A_695_457#_c_828_n 0.00139327f $X=4.395 $Y=0.9
+ $X2=0 $Y2=0
cc_501 N_A_830_359#_c_524_n N_A_695_457#_c_828_n 0.0386081f $X=4.355 $Y=1.96
+ $X2=0 $Y2=0
cc_502 N_A_830_359#_M1012_g N_A_695_457#_c_829_n 0.00230788f $X=4.395 $Y=0.9
+ $X2=0 $Y2=0
cc_503 N_A_830_359#_c_524_n N_A_695_457#_c_829_n 0.0266749f $X=4.355 $Y=1.96
+ $X2=0 $Y2=0
cc_504 N_A_830_359#_c_542_n N_A_695_457#_c_829_n 0.0115313f $X=5.82 $Y=0.99
+ $X2=0 $Y2=0
cc_505 N_A_830_359#_c_542_n N_A_695_457#_c_830_n 0.0585986f $X=5.82 $Y=0.99
+ $X2=0 $Y2=0
cc_506 N_A_830_359#_c_526_n N_A_695_457#_c_830_n 0.0159069f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_507 N_A_830_359#_c_542_n N_A_695_457#_c_831_n 0.00636706f $X=5.82 $Y=0.99
+ $X2=0 $Y2=0
cc_508 N_A_830_359#_c_525_n N_A_695_457#_c_831_n 0.00593666f $X=5.985 $Y=0.855
+ $X2=0 $Y2=0
cc_509 N_A_830_359#_c_526_n N_A_695_457#_c_831_n 0.00831051f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_510 N_A_830_359#_c_527_n N_A_695_457#_c_839_n 0.00932733f $X=4.24 $Y=2.21
+ $X2=0 $Y2=0
cc_511 N_A_830_359#_c_527_n N_A_695_457#_c_875_n 8.25025e-19 $X=4.24 $Y=2.21
+ $X2=0 $Y2=0
cc_512 N_A_830_359#_c_527_n N_A_306_96#_M1019_g 0.0341022f $X=4.24 $Y=2.21 $X2=0
+ $Y2=0
cc_513 N_A_830_359#_c_527_n N_A_306_96#_c_969_n 0.00845256f $X=4.24 $Y=2.21
+ $X2=0 $Y2=0
cc_514 N_A_830_359#_c_530_n N_A_306_96#_c_969_n 0.00611621f $X=6.145 $Y=2.03
+ $X2=0 $Y2=0
cc_515 N_A_830_359#_c_530_n N_A_306_96#_M1015_g 0.00116389f $X=6.145 $Y=2.03
+ $X2=0 $Y2=0
cc_516 N_A_830_359#_c_526_n N_A_306_96#_M1015_g 4.46008e-19 $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_517 N_A_830_359#_c_530_n N_A_306_96#_c_957_n 6.78448e-19 $X=6.145 $Y=2.03
+ $X2=0 $Y2=0
cc_518 N_A_830_359#_c_526_n N_A_306_96#_c_957_n 0.00196898f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_519 N_A_830_359#_c_525_n N_A_1266_74#_c_1268_n 0.03852f $X=5.985 $Y=0.855
+ $X2=0 $Y2=0
cc_520 N_A_830_359#_c_530_n N_A_1266_74#_c_1281_n 0.0206296f $X=6.145 $Y=2.03
+ $X2=0 $Y2=0
cc_521 N_A_830_359#_c_526_n N_A_1266_74#_c_1281_n 0.00813918f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_522 N_A_830_359#_c_526_n N_A_1266_74#_c_1272_n 0.0129729f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_523 N_A_830_359#_c_527_n N_VPWR_c_1480_n 0.00274139f $X=4.24 $Y=2.21 $X2=0
+ $Y2=0
cc_524 N_A_830_359#_c_542_n N_VPWR_c_1482_n 0.00363609f $X=5.82 $Y=0.99 $X2=0
+ $Y2=0
cc_525 N_A_830_359#_c_530_n N_VPWR_c_1482_n 0.0405057f $X=6.145 $Y=2.03 $X2=0
+ $Y2=0
cc_526 N_A_830_359#_c_530_n N_VPWR_c_1491_n 0.00670512f $X=6.145 $Y=2.03 $X2=0
+ $Y2=0
cc_527 N_A_830_359#_c_527_n N_VPWR_c_1475_n 9.49986e-19 $X=4.24 $Y=2.21 $X2=0
+ $Y2=0
cc_528 N_A_830_359#_c_530_n N_VPWR_c_1475_n 0.00907985f $X=6.145 $Y=2.03 $X2=0
+ $Y2=0
cc_529 N_A_830_359#_c_542_n N_VGND_M1004_d 0.00954133f $X=5.82 $Y=0.99 $X2=0
+ $Y2=0
cc_530 N_A_830_359#_c_542_n A_894_138# 0.00503032f $X=5.82 $Y=0.99 $X2=-0.19
+ $Y2=-0.245
cc_531 N_RESET_B_c_608_n N_A_695_457#_M1026_g 0.0212385f $X=4.71 $Y=0.18 $X2=0
+ $Y2=0
cc_532 N_RESET_B_c_613_n N_A_695_457#_M1026_g 0.00219471f $X=4.875 $Y=1.26 $X2=0
+ $Y2=0
cc_533 N_RESET_B_c_625_n N_A_695_457#_c_833_n 0.0113891f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_534 N_RESET_B_c_623_n N_A_695_457#_c_827_n 0.0128588f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_535 N_RESET_B_c_623_n N_A_695_457#_c_861_n 0.00774799f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_536 N_RESET_B_c_618_n N_A_695_457#_c_828_n 0.00234023f $X=4.86 $Y=2.21 $X2=0
+ $Y2=0
cc_537 N_RESET_B_c_611_n N_A_695_457#_c_828_n 0.0056545f $X=4.875 $Y=1.795 $X2=0
+ $Y2=0
cc_538 N_RESET_B_c_623_n N_A_695_457#_c_828_n 0.0207498f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_539 N_RESET_B_c_626_n N_A_695_457#_c_828_n 0.00237384f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_540 N_RESET_B_c_627_n N_A_695_457#_c_828_n 0.0234789f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_541 N_RESET_B_c_631_n N_A_695_457#_c_828_n 0.0103538f $X=4.875 $Y=2.002 $X2=0
+ $Y2=0
cc_542 N_RESET_B_c_613_n N_A_695_457#_c_829_n 0.00393752f $X=4.875 $Y=1.26 $X2=0
+ $Y2=0
cc_543 N_RESET_B_c_611_n N_A_695_457#_c_830_n 0.0121734f $X=4.875 $Y=1.795 $X2=0
+ $Y2=0
cc_544 N_RESET_B_c_613_n N_A_695_457#_c_830_n 0.00449896f $X=4.875 $Y=1.26 $X2=0
+ $Y2=0
cc_545 N_RESET_B_c_623_n N_A_695_457#_c_830_n 0.00353489f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_546 N_RESET_B_c_625_n N_A_695_457#_c_830_n 0.0084128f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_547 N_RESET_B_c_626_n N_A_695_457#_c_830_n 0.00351517f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_548 N_RESET_B_c_627_n N_A_695_457#_c_830_n 0.01951f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_549 N_RESET_B_c_631_n N_A_695_457#_c_830_n 0.00785354f $X=4.875 $Y=2.002
+ $X2=0 $Y2=0
cc_550 N_RESET_B_c_613_n N_A_695_457#_c_831_n 0.0103083f $X=4.875 $Y=1.26 $X2=0
+ $Y2=0
cc_551 N_RESET_B_c_625_n N_A_695_457#_c_831_n 0.00409962f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_552 N_RESET_B_c_618_n N_A_695_457#_c_837_n 0.00887731f $X=4.86 $Y=2.21 $X2=0
+ $Y2=0
cc_553 N_RESET_B_c_623_n N_A_695_457#_c_837_n 0.0041068f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_554 N_RESET_B_c_625_n N_A_695_457#_c_837_n 4.57663e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_555 N_RESET_B_c_626_n N_A_695_457#_c_837_n 0.00893467f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_556 N_RESET_B_c_627_n N_A_695_457#_c_837_n 0.0191542f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_557 N_RESET_B_c_631_n N_A_695_457#_c_837_n 0.00191227f $X=4.875 $Y=2.002
+ $X2=0 $Y2=0
cc_558 N_RESET_B_c_623_n N_A_695_457#_c_838_n 0.00693162f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_559 N_RESET_B_c_618_n N_A_695_457#_c_839_n 7.07248e-19 $X=4.86 $Y=2.21 $X2=0
+ $Y2=0
cc_560 N_RESET_B_c_623_n N_A_695_457#_c_839_n 0.00694709f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_561 N_RESET_B_c_618_n N_A_695_457#_c_875_n 0.00379552f $X=4.86 $Y=2.21 $X2=0
+ $Y2=0
cc_562 N_RESET_B_c_623_n N_A_306_96#_M1011_g 0.00818514f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_563 N_RESET_B_c_608_n N_A_306_96#_c_952_n 0.010267f $X=4.71 $Y=0.18 $X2=0
+ $Y2=0
cc_564 N_RESET_B_c_623_n N_A_306_96#_c_964_n 0.00258458f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_565 N_RESET_B_c_608_n N_A_306_96#_c_955_n 0.00526413f $X=4.71 $Y=0.18 $X2=0
+ $Y2=0
cc_566 N_RESET_B_c_623_n N_A_306_96#_M1019_g 0.00260456f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_567 N_RESET_B_c_618_n N_A_306_96#_c_969_n 0.00852675f $X=4.86 $Y=2.21 $X2=0
+ $Y2=0
cc_568 N_RESET_B_c_625_n N_A_306_96#_M1015_g 0.00898574f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_569 N_RESET_B_c_625_n N_A_306_96#_c_956_n 0.00802201f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_570 N_RESET_B_c_625_n N_A_306_96#_c_957_n 3.42215e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_571 N_RESET_B_M1008_g N_A_306_96#_c_959_n 0.00308278f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_572 N_RESET_B_c_608_n N_A_306_96#_c_959_n 0.00906252f $X=4.71 $Y=0.18 $X2=0
+ $Y2=0
cc_573 N_RESET_B_c_624_n N_A_306_96#_c_960_n 7.86393e-19 $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_574 N_RESET_B_c_614_n N_A_306_96#_c_960_n 0.0080451f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_575 N_RESET_B_c_615_n N_A_306_96#_c_960_n 0.0598064f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_576 N_RESET_B_M1008_g N_A_306_96#_c_961_n 0.00122712f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_577 N_RESET_B_c_615_n N_A_306_96#_c_961_n 8.29766e-19 $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_578 N_RESET_B_c_617_n N_A_306_96#_c_976_n 0.00234359f $X=0.945 $Y=2.375 $X2=0
+ $Y2=0
cc_579 N_RESET_B_c_623_n N_A_306_96#_c_976_n 0.0320911f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_580 N_RESET_B_c_624_n N_A_306_96#_c_976_n 0.00217735f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_581 N_RESET_B_c_615_n N_A_306_96#_c_976_n 0.0133824f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_582 N_RESET_B_c_630_n N_A_306_96#_c_976_n 0.00158946f $X=1.155 $Y=1.975 $X2=0
+ $Y2=0
cc_583 N_RESET_B_c_623_n N_A_306_96#_c_1035_n 0.00202299f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_584 N_RESET_B_M1028_g N_A_1518_203#_c_1149_n 0.00652196f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_585 N_RESET_B_c_621_n N_A_1518_203#_c_1150_n 0.022618f $X=8.26 $Y=2.39 $X2=0
+ $Y2=0
cc_586 N_RESET_B_c_625_n N_A_1518_203#_c_1150_n 0.00706641f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_587 N_RESET_B_c_628_n N_A_1518_203#_c_1150_n 0.00231702f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_588 N_RESET_B_c_632_n N_A_1518_203#_c_1150_n 0.00228452f $X=8.18 $Y=2.09
+ $X2=0 $Y2=0
cc_589 N_RESET_B_c_621_n N_A_1518_203#_c_1151_n 0.012219f $X=8.26 $Y=2.39 $X2=0
+ $Y2=0
cc_590 N_RESET_B_M1028_g N_A_1518_203#_M1014_g 0.0166359f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_591 N_RESET_B_M1028_g N_A_1518_203#_c_1142_n 0.0133984f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_592 N_RESET_B_M1028_g N_A_1518_203#_c_1143_n 0.0149634f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_593 N_RESET_B_M1028_g N_A_1518_203#_c_1144_n 0.00216035f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_594 N_RESET_B_M1028_g N_A_1518_203#_c_1154_n 0.00169886f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_595 N_RESET_B_c_621_n N_A_1518_203#_c_1154_n 6.9451e-19 $X=8.26 $Y=2.39 $X2=0
+ $Y2=0
cc_596 N_RESET_B_c_628_n N_A_1518_203#_c_1154_n 4.76192e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_597 N_RESET_B_c_632_n N_A_1518_203#_c_1154_n 0.00873148f $X=8.18 $Y=2.09
+ $X2=0 $Y2=0
cc_598 N_RESET_B_M1028_g N_A_1518_203#_c_1146_n 0.00118187f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_599 N_RESET_B_c_625_n N_A_1518_203#_c_1146_n 3.17521e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_600 N_RESET_B_M1028_g N_A_1518_203#_c_1147_n 0.021263f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_601 N_RESET_B_c_621_n N_A_1518_203#_c_1156_n 0.00637785f $X=8.26 $Y=2.39
+ $X2=0 $Y2=0
cc_602 N_RESET_B_c_632_n N_A_1518_203#_c_1156_n 0.00174345f $X=8.18 $Y=2.09
+ $X2=0 $Y2=0
cc_603 N_RESET_B_c_621_n N_A_1518_203#_c_1157_n 0.00534913f $X=8.26 $Y=2.39
+ $X2=0 $Y2=0
cc_604 N_RESET_B_c_628_n N_A_1518_203#_c_1157_n 5.01506e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_605 N_RESET_B_c_632_n N_A_1518_203#_c_1157_n 0.0175397f $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_606 N_RESET_B_c_625_n N_A_1266_74#_M1015_d 0.00283611f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_607 N_RESET_B_M1028_g N_A_1266_74#_M1017_g 0.0757442f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_608 N_RESET_B_M1028_g N_A_1266_74#_c_1274_n 0.00953304f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_609 N_RESET_B_c_621_n N_A_1266_74#_c_1274_n 0.0206573f $X=8.26 $Y=2.39 $X2=0
+ $Y2=0
cc_610 N_RESET_B_c_632_n N_A_1266_74#_c_1274_n 3.48207e-19 $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_611 N_RESET_B_c_621_n N_A_1266_74#_c_1275_n 0.00915627f $X=8.26 $Y=2.39 $X2=0
+ $Y2=0
cc_612 N_RESET_B_M1028_g N_A_1266_74#_c_1262_n 0.00996674f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_613 N_RESET_B_c_625_n N_A_1266_74#_c_1281_n 0.0174694f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_614 N_RESET_B_c_625_n N_A_1266_74#_c_1303_n 0.0206747f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_615 N_RESET_B_M1028_g N_A_1266_74#_c_1282_n 0.00109662f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_616 N_RESET_B_c_621_n N_A_1266_74#_c_1282_n 0.00116333f $X=8.26 $Y=2.39 $X2=0
+ $Y2=0
cc_617 N_RESET_B_c_625_n N_A_1266_74#_c_1282_n 0.0211228f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_618 N_RESET_B_c_628_n N_A_1266_74#_c_1282_n 0.00228452f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_619 N_RESET_B_c_632_n N_A_1266_74#_c_1282_n 0.0236542f $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_620 N_RESET_B_M1028_g N_A_1266_74#_c_1270_n 0.011972f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_621 N_RESET_B_c_621_n N_A_1266_74#_c_1270_n 0.00135016f $X=8.26 $Y=2.39 $X2=0
+ $Y2=0
cc_622 N_RESET_B_c_625_n N_A_1266_74#_c_1270_n 0.00476106f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_623 N_RESET_B_c_628_n N_A_1266_74#_c_1270_n 0.00823149f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_624 N_RESET_B_c_632_n N_A_1266_74#_c_1270_n 0.02904f $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_625 N_RESET_B_c_625_n N_A_1266_74#_c_1272_n 0.00599756f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_626 N_RESET_B_M1028_g N_A_1266_74#_c_1273_n 0.00110907f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_627 N_RESET_B_c_623_n N_VPWR_M1006_d 0.00582056f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_628 N_RESET_B_c_622_n N_VPWR_c_1478_n 0.0080317f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_629 N_RESET_B_c_618_n N_VPWR_c_1480_n 0.00274139f $X=4.86 $Y=2.21 $X2=0 $Y2=0
cc_630 N_RESET_B_c_618_n N_VPWR_c_1482_n 0.0078214f $X=4.86 $Y=2.21 $X2=0 $Y2=0
cc_631 N_RESET_B_c_611_n N_VPWR_c_1482_n 0.00126145f $X=4.875 $Y=1.795 $X2=0
+ $Y2=0
cc_632 N_RESET_B_c_625_n N_VPWR_c_1482_n 0.0317336f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_633 N_RESET_B_c_626_n N_VPWR_c_1482_n 5.51604e-19 $X=5.185 $Y=2.035 $X2=0
+ $Y2=0
cc_634 N_RESET_B_c_627_n N_VPWR_c_1482_n 0.023147f $X=5.04 $Y=2.035 $X2=0 $Y2=0
cc_635 N_RESET_B_c_631_n N_VPWR_c_1482_n 0.00289108f $X=4.875 $Y=2.002 $X2=0
+ $Y2=0
cc_636 N_RESET_B_c_621_n N_VPWR_c_1483_n 0.00888753f $X=8.26 $Y=2.39 $X2=0 $Y2=0
cc_637 N_RESET_B_c_628_n N_VPWR_c_1483_n 0.00171912f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_638 N_RESET_B_c_632_n N_VPWR_c_1483_n 0.0244512f $X=8.18 $Y=2.09 $X2=0 $Y2=0
cc_639 N_RESET_B_c_621_n N_VPWR_c_1484_n 0.00510653f $X=8.26 $Y=2.39 $X2=0 $Y2=0
cc_640 N_RESET_B_c_622_n N_VPWR_c_1488_n 0.00378953f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_641 N_RESET_B_c_618_n N_VPWR_c_1475_n 9.49986e-19 $X=4.86 $Y=2.21 $X2=0 $Y2=0
cc_642 N_RESET_B_c_621_n N_VPWR_c_1475_n 0.0052212f $X=8.26 $Y=2.39 $X2=0 $Y2=0
cc_643 N_RESET_B_c_622_n N_VPWR_c_1475_n 0.00369031f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_644 N_RESET_B_M1008_g N_A_30_78#_c_1624_n 0.00433444f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_645 N_RESET_B_c_622_n N_A_30_78#_c_1631_n 2.11957e-19 $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_646 N_RESET_B_M1008_g N_A_30_78#_c_1625_n 0.0089809f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_647 N_RESET_B_c_607_n N_A_30_78#_c_1625_n 0.0116119f $X=1.072 $Y=1.893 $X2=0
+ $Y2=0
cc_648 N_RESET_B_c_617_n N_A_30_78#_c_1625_n 0.00433638f $X=0.945 $Y=2.375 $X2=0
+ $Y2=0
cc_649 N_RESET_B_c_624_n N_A_30_78#_c_1625_n 0.00186952f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_650 N_RESET_B_c_614_n N_A_30_78#_c_1625_n 0.00558005f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_651 N_RESET_B_c_615_n N_A_30_78#_c_1625_n 0.069302f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_652 N_RESET_B_c_630_n N_A_30_78#_c_1625_n 0.00612462f $X=1.155 $Y=1.975 $X2=0
+ $Y2=0
cc_653 N_RESET_B_c_617_n N_A_30_78#_c_1633_n 0.0101591f $X=0.945 $Y=2.375 $X2=0
+ $Y2=0
cc_654 N_RESET_B_c_622_n N_A_30_78#_c_1633_n 0.0115083f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_655 N_RESET_B_c_623_n N_A_30_78#_c_1633_n 0.00550786f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_656 N_RESET_B_c_624_n N_A_30_78#_c_1633_n 0.0094643f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_657 N_RESET_B_c_615_n N_A_30_78#_c_1633_n 0.0173369f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_658 N_RESET_B_c_630_n N_A_30_78#_c_1633_n 0.003052f $X=1.155 $Y=1.975 $X2=0
+ $Y2=0
cc_659 N_RESET_B_c_623_n N_A_30_78#_c_1634_n 0.0033801f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_660 N_RESET_B_c_623_n N_A_30_78#_c_1635_n 0.0225207f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_661 N_RESET_B_c_623_n N_A_30_78#_c_1636_n 0.0101888f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_662 N_RESET_B_c_623_n N_A_30_78#_c_1627_n 0.0138311f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_663 N_RESET_B_M1008_g N_A_30_78#_c_1628_n 9.29579e-19 $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_664 N_RESET_B_c_617_n N_A_30_78#_c_1638_n 7.56365e-19 $X=0.945 $Y=2.375 $X2=0
+ $Y2=0
cc_665 N_RESET_B_c_622_n N_A_30_78#_c_1638_n 0.00246461f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_666 N_RESET_B_c_623_n N_A_30_78#_c_1639_n 0.00946737f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_667 N_RESET_B_c_623_n N_A_30_78#_c_1630_n 0.00584074f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_668 N_RESET_B_M1008_g N_VGND_c_1791_n 0.00257803f $X=0.9 $Y=0.6 $X2=0 $Y2=0
cc_669 N_RESET_B_c_608_n N_VGND_c_1791_n 0.0200565f $X=4.71 $Y=0.18 $X2=0 $Y2=0
cc_670 N_RESET_B_c_614_n N_VGND_c_1791_n 0.00181416f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_671 N_RESET_B_c_615_n N_VGND_c_1791_n 0.0144384f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_672 N_RESET_B_c_608_n N_VGND_c_1792_n 0.0257653f $X=4.71 $Y=0.18 $X2=0 $Y2=0
cc_673 N_RESET_B_M1028_g N_VGND_c_1793_n 0.0058325f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_674 N_RESET_B_c_609_n N_VGND_c_1797_n 0.00764766f $X=0.975 $Y=0.18 $X2=0
+ $Y2=0
cc_675 N_RESET_B_c_608_n N_VGND_c_1799_n 0.0221705f $X=4.71 $Y=0.18 $X2=0 $Y2=0
cc_676 N_RESET_B_c_608_n N_VGND_c_1800_n 0.0656472f $X=4.71 $Y=0.18 $X2=0 $Y2=0
cc_677 N_RESET_B_M1028_g N_VGND_c_1802_n 0.00552345f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_678 N_RESET_B_c_608_n N_VGND_c_1807_n 0.0939206f $X=4.71 $Y=0.18 $X2=0 $Y2=0
cc_679 N_RESET_B_c_609_n N_VGND_c_1807_n 0.0105042f $X=0.975 $Y=0.18 $X2=0 $Y2=0
cc_680 N_RESET_B_M1028_g N_VGND_c_1807_n 0.00534666f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_681 N_A_695_457#_c_838_n N_A_306_96#_c_965_n 0.00392476f $X=3.93 $Y=2.562
+ $X2=0 $Y2=0
cc_682 N_A_695_457#_c_827_n N_A_306_96#_c_955_n 6.61176e-19 $X=4.015 $Y=2.4
+ $X2=0 $Y2=0
cc_683 N_A_695_457#_c_832_n N_A_306_96#_c_955_n 0.00203911f $X=4.015 $Y=0.86
+ $X2=0 $Y2=0
cc_684 N_A_695_457#_c_827_n N_A_306_96#_M1019_g 0.00138382f $X=4.015 $Y=2.4
+ $X2=0 $Y2=0
cc_685 N_A_695_457#_c_838_n N_A_306_96#_M1019_g 0.0118268f $X=3.93 $Y=2.562
+ $X2=0 $Y2=0
cc_686 N_A_695_457#_c_833_n N_A_306_96#_c_969_n 0.0104018f $X=5.88 $Y=1.66 $X2=0
+ $Y2=0
cc_687 N_A_695_457#_c_861_n N_A_306_96#_c_969_n 0.00193774f $X=4.615 $Y=2.485
+ $X2=0 $Y2=0
cc_688 N_A_695_457#_c_837_n N_A_306_96#_c_969_n 0.00523168f $X=5.085 $Y=2.485
+ $X2=0 $Y2=0
cc_689 N_A_695_457#_c_838_n N_A_306_96#_c_969_n 0.00450392f $X=3.93 $Y=2.562
+ $X2=0 $Y2=0
cc_690 N_A_695_457#_c_875_n N_A_306_96#_c_969_n 0.001324f $X=4.7 $Y=2.445 $X2=0
+ $Y2=0
cc_691 N_A_695_457#_c_833_n N_A_306_96#_M1015_g 0.00888826f $X=5.88 $Y=1.66
+ $X2=0 $Y2=0
cc_692 N_A_695_457#_c_833_n N_A_306_96#_c_957_n 0.00427682f $X=5.88 $Y=1.66
+ $X2=0 $Y2=0
cc_693 N_A_695_457#_c_831_n N_A_306_96#_c_957_n 0.00245186f $X=5.485 $Y=1.41
+ $X2=0 $Y2=0
cc_694 N_A_695_457#_c_861_n N_VPWR_M1003_d 0.00582643f $X=4.615 $Y=2.485 $X2=0
+ $Y2=0
cc_695 N_A_695_457#_c_828_n N_VPWR_M1003_d 4.43648e-19 $X=4.7 $Y=2.32 $X2=0
+ $Y2=0
cc_696 N_A_695_457#_c_875_n N_VPWR_M1003_d 0.0021968f $X=4.7 $Y=2.445 $X2=0
+ $Y2=0
cc_697 N_A_695_457#_c_861_n N_VPWR_c_1480_n 0.0180683f $X=4.615 $Y=2.485 $X2=0
+ $Y2=0
cc_698 N_A_695_457#_c_875_n N_VPWR_c_1480_n 0.00862169f $X=4.7 $Y=2.445 $X2=0
+ $Y2=0
cc_699 N_A_695_457#_c_837_n N_VPWR_c_1481_n 0.00589153f $X=5.085 $Y=2.485 $X2=0
+ $Y2=0
cc_700 N_A_695_457#_c_875_n N_VPWR_c_1481_n 5.93009e-19 $X=4.7 $Y=2.445 $X2=0
+ $Y2=0
cc_701 N_A_695_457#_c_833_n N_VPWR_c_1482_n 0.0131452f $X=5.88 $Y=1.66 $X2=0
+ $Y2=0
cc_702 N_A_695_457#_c_830_n N_VPWR_c_1482_n 0.0133374f $X=5.485 $Y=1.41 $X2=0
+ $Y2=0
cc_703 N_A_695_457#_c_831_n N_VPWR_c_1482_n 0.00741213f $X=5.485 $Y=1.41 $X2=0
+ $Y2=0
cc_704 N_A_695_457#_c_837_n N_VPWR_c_1482_n 0.0177113f $X=5.085 $Y=2.485 $X2=0
+ $Y2=0
cc_705 N_A_695_457#_c_861_n N_VPWR_c_1490_n 0.00180774f $X=4.615 $Y=2.485 $X2=0
+ $Y2=0
cc_706 N_A_695_457#_c_838_n N_VPWR_c_1490_n 0.0146861f $X=3.93 $Y=2.562 $X2=0
+ $Y2=0
cc_707 N_A_695_457#_c_833_n N_VPWR_c_1475_n 9.14192e-19 $X=5.88 $Y=1.66 $X2=0
+ $Y2=0
cc_708 N_A_695_457#_c_861_n N_VPWR_c_1475_n 0.00449748f $X=4.615 $Y=2.485 $X2=0
+ $Y2=0
cc_709 N_A_695_457#_c_837_n N_VPWR_c_1475_n 0.0102762f $X=5.085 $Y=2.485 $X2=0
+ $Y2=0
cc_710 N_A_695_457#_c_838_n N_VPWR_c_1475_n 0.0191974f $X=3.93 $Y=2.562 $X2=0
+ $Y2=0
cc_711 N_A_695_457#_c_875_n N_VPWR_c_1475_n 0.0021032f $X=4.7 $Y=2.445 $X2=0
+ $Y2=0
cc_712 N_A_695_457#_c_827_n N_A_30_78#_c_1626_n 0.00500199f $X=4.015 $Y=2.4
+ $X2=0 $Y2=0
cc_713 N_A_695_457#_M1009_d N_A_30_78#_c_1636_n 0.00209257f $X=3.475 $Y=2.285
+ $X2=0 $Y2=0
cc_714 N_A_695_457#_c_827_n N_A_30_78#_c_1636_n 0.0108294f $X=4.015 $Y=2.4 $X2=0
+ $Y2=0
cc_715 N_A_695_457#_c_838_n N_A_30_78#_c_1636_n 0.0151296f $X=3.93 $Y=2.562
+ $X2=0 $Y2=0
cc_716 N_A_695_457#_c_827_n N_A_30_78#_c_1627_n 0.0550948f $X=4.015 $Y=2.4 $X2=0
+ $Y2=0
cc_717 N_A_695_457#_c_838_n N_A_30_78#_c_1639_n 0.0103876f $X=3.93 $Y=2.562
+ $X2=0 $Y2=0
cc_718 N_A_695_457#_c_832_n N_A_30_78#_c_1629_n 0.0144099f $X=4.015 $Y=0.86
+ $X2=0 $Y2=0
cc_719 N_A_695_457#_c_827_n N_A_30_78#_c_1630_n 0.0131435f $X=4.015 $Y=2.4 $X2=0
+ $Y2=0
cc_720 N_A_695_457#_c_832_n N_A_30_78#_c_1630_n 0.0101207f $X=4.015 $Y=0.86
+ $X2=0 $Y2=0
cc_721 N_A_695_457#_c_827_n A_785_457# 0.00168676f $X=4.015 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_722 N_A_695_457#_c_839_n A_785_457# 4.77189e-19 $X=4.215 $Y=2.562 $X2=-0.19
+ $Y2=-0.245
cc_723 N_A_695_457#_M1026_g N_VGND_c_1800_n 0.00178007f $X=5.44 $Y=0.74 $X2=0
+ $Y2=0
cc_724 N_A_695_457#_M1026_g N_VGND_c_1801_n 0.00309023f $X=5.44 $Y=0.74 $X2=0
+ $Y2=0
cc_725 N_A_695_457#_M1026_g N_VGND_c_1807_n 0.00390562f $X=5.44 $Y=0.74 $X2=0
+ $Y2=0
cc_726 N_A_306_96#_M1016_g N_A_1518_203#_M1014_g 0.0368892f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_727 N_A_306_96#_M1016_g N_A_1518_203#_c_1142_n 0.0235039f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_728 N_A_306_96#_M1016_g N_A_1518_203#_c_1146_n 3.81559e-19 $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_729 N_A_306_96#_M1016_g N_A_1518_203#_c_1147_n 0.0205557f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_730 N_A_306_96#_c_957_n N_A_1266_74#_c_1268_n 2.4837e-19 $X=6.475 $Y=1.66
+ $X2=0 $Y2=0
cc_731 N_A_306_96#_M1015_g N_A_1266_74#_c_1281_n 0.00801796f $X=6.385 $Y=2.385
+ $X2=0 $Y2=0
cc_732 N_A_306_96#_c_956_n N_A_1266_74#_c_1281_n 0.00695524f $X=7.23 $Y=1.66
+ $X2=0 $Y2=0
cc_733 N_A_306_96#_c_957_n N_A_1266_74#_c_1281_n 0.00199946f $X=6.475 $Y=1.66
+ $X2=0 $Y2=0
cc_734 N_A_306_96#_M1016_g N_A_1266_74#_c_1269_n 0.00507341f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_735 N_A_306_96#_c_956_n N_A_1266_74#_c_1282_n 3.51038e-19 $X=7.23 $Y=1.66
+ $X2=0 $Y2=0
cc_736 N_A_306_96#_M1016_g N_A_1266_74#_c_1271_n 0.00127921f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_737 N_A_306_96#_c_956_n N_A_1266_74#_c_1272_n 0.00490084f $X=7.23 $Y=1.66
+ $X2=0 $Y2=0
cc_738 N_A_306_96#_c_957_n N_A_1266_74#_c_1272_n 0.00528124f $X=6.475 $Y=1.66
+ $X2=0 $Y2=0
cc_739 N_A_306_96#_M1016_g N_A_1266_74#_c_1272_n 2.86702e-19 $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_740 N_A_306_96#_M1011_g N_VPWR_c_1479_n 0.0084462f $X=2.375 $Y=2.45 $X2=0
+ $Y2=0
cc_741 N_A_306_96#_c_964_n N_VPWR_c_1479_n 0.00157439f $X=2.885 $Y=3.075 $X2=0
+ $Y2=0
cc_742 N_A_306_96#_c_966_n N_VPWR_c_1479_n 0.00261603f $X=2.96 $Y=3.15 $X2=0
+ $Y2=0
cc_743 N_A_306_96#_M1019_g N_VPWR_c_1480_n 0.00671018f $X=3.85 $Y=2.495 $X2=0
+ $Y2=0
cc_744 N_A_306_96#_c_969_n N_VPWR_c_1480_n 0.0250293f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_745 N_A_306_96#_c_969_n N_VPWR_c_1481_n 0.0218819f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_746 N_A_306_96#_c_969_n N_VPWR_c_1482_n 0.0259878f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_747 N_A_306_96#_M1015_g N_VPWR_c_1482_n 0.00308789f $X=6.385 $Y=2.385 $X2=0
+ $Y2=0
cc_748 N_A_306_96#_c_974_n N_VPWR_c_1482_n 0.00312383f $X=6.385 $Y=3.15 $X2=0
+ $Y2=0
cc_749 N_A_306_96#_M1011_g N_VPWR_c_1490_n 0.00404449f $X=2.375 $Y=2.45 $X2=0
+ $Y2=0
cc_750 N_A_306_96#_c_966_n N_VPWR_c_1490_n 0.0424196f $X=2.96 $Y=3.15 $X2=0
+ $Y2=0
cc_751 N_A_306_96#_c_969_n N_VPWR_c_1491_n 0.0203278f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_752 N_A_306_96#_M1011_g N_VPWR_c_1475_n 0.00492022f $X=2.375 $Y=2.45 $X2=0
+ $Y2=0
cc_753 N_A_306_96#_c_965_n N_VPWR_c_1475_n 0.0237205f $X=3.775 $Y=3.15 $X2=0
+ $Y2=0
cc_754 N_A_306_96#_c_966_n N_VPWR_c_1475_n 0.00695678f $X=2.96 $Y=3.15 $X2=0
+ $Y2=0
cc_755 N_A_306_96#_c_969_n N_VPWR_c_1475_n 0.053457f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_756 N_A_306_96#_c_973_n N_VPWR_c_1475_n 0.00423956f $X=3.85 $Y=3.15 $X2=0
+ $Y2=0
cc_757 N_A_306_96#_c_974_n N_VPWR_c_1475_n 0.0128115f $X=6.385 $Y=3.15 $X2=0
+ $Y2=0
cc_758 N_A_306_96#_c_959_n N_A_30_78#_c_1625_n 0.00411959f $X=1.675 $Y=0.625
+ $X2=0 $Y2=0
cc_759 N_A_306_96#_c_961_n N_A_30_78#_c_1625_n 0.00499576f $X=1.647 $Y=1.055
+ $X2=0 $Y2=0
cc_760 N_A_306_96#_c_976_n N_A_30_78#_c_1633_n 0.00467759f $X=1.54 $Y=2.092
+ $X2=0 $Y2=0
cc_761 N_A_306_96#_M1006_s N_A_30_78#_c_1634_n 0.00895973f $X=1.54 $Y=1.95 $X2=0
+ $Y2=0
cc_762 N_A_306_96#_c_976_n N_A_30_78#_c_1634_n 0.017969f $X=1.54 $Y=2.092 $X2=0
+ $Y2=0
cc_763 N_A_306_96#_M1011_g N_A_30_78#_c_1635_n 0.0141403f $X=2.375 $Y=2.45 $X2=0
+ $Y2=0
cc_764 N_A_306_96#_c_964_n N_A_30_78#_c_1635_n 0.0147996f $X=2.885 $Y=3.075
+ $X2=0 $Y2=0
cc_765 N_A_306_96#_c_953_n N_A_30_78#_c_1626_n 0.00463589f $X=3.43 $Y=1.275
+ $X2=0 $Y2=0
cc_766 N_A_306_96#_c_955_n N_A_30_78#_c_1626_n 0.00459249f $X=3.505 $Y=1.2 $X2=0
+ $Y2=0
cc_767 N_A_306_96#_M1019_g N_A_30_78#_c_1636_n 0.00134037f $X=3.85 $Y=2.495
+ $X2=0 $Y2=0
cc_768 N_A_306_96#_c_954_n N_A_30_78#_c_1627_n 8.13937e-19 $X=3.095 $Y=1.275
+ $X2=0 $Y2=0
cc_769 N_A_306_96#_c_964_n N_A_30_78#_c_1639_n 0.0101189f $X=2.885 $Y=3.075
+ $X2=0 $Y2=0
cc_770 N_A_306_96#_c_965_n N_A_30_78#_c_1639_n 0.00467498f $X=3.775 $Y=3.15
+ $X2=0 $Y2=0
cc_771 N_A_306_96#_c_953_n N_A_30_78#_c_1629_n 0.00192283f $X=3.43 $Y=1.275
+ $X2=0 $Y2=0
cc_772 N_A_306_96#_c_955_n N_A_30_78#_c_1629_n 0.00435411f $X=3.505 $Y=1.2 $X2=0
+ $Y2=0
cc_773 N_A_306_96#_c_953_n N_A_30_78#_c_1630_n 0.013367f $X=3.43 $Y=1.275 $X2=0
+ $Y2=0
cc_774 N_A_306_96#_c_954_n N_A_30_78#_c_1630_n 2.85666e-19 $X=3.095 $Y=1.275
+ $X2=0 $Y2=0
cc_775 N_A_306_96#_c_989_n N_VGND_M1030_d 0.00726965f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_776 N_A_306_96#_c_959_n N_VGND_c_1791_n 0.0388156f $X=1.675 $Y=0.625 $X2=0
+ $Y2=0
cc_777 N_A_306_96#_c_952_n N_VGND_c_1792_n 0.00242994f $X=2.5 $Y=1.41 $X2=0
+ $Y2=0
cc_778 N_A_306_96#_c_959_n N_VGND_c_1792_n 0.0171529f $X=1.675 $Y=0.625 $X2=0
+ $Y2=0
cc_779 N_A_306_96#_c_989_n N_VGND_c_1792_n 0.0232685f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_780 N_A_306_96#_M1016_g N_VGND_c_1793_n 5.78056e-19 $X=7.305 $Y=0.615 $X2=0
+ $Y2=0
cc_781 N_A_306_96#_c_959_n N_VGND_c_1799_n 0.0170748f $X=1.675 $Y=0.625 $X2=0
+ $Y2=0
cc_782 N_A_306_96#_M1016_g N_VGND_c_1801_n 9.33926e-19 $X=7.305 $Y=0.615 $X2=0
+ $Y2=0
cc_783 N_A_306_96#_c_952_n N_VGND_c_1807_n 8.51577e-19 $X=2.5 $Y=1.41 $X2=0
+ $Y2=0
cc_784 N_A_306_96#_c_959_n N_VGND_c_1807_n 0.0126098f $X=1.675 $Y=0.625 $X2=0
+ $Y2=0
cc_785 N_A_1518_203#_c_1143_n N_A_1266_74#_M1017_g 0.0107164f $X=8.615 $Y=1.1
+ $X2=0 $Y2=0
cc_786 N_A_1518_203#_c_1144_n N_A_1266_74#_M1017_g 0.0159617f $X=8.78 $Y=0.615
+ $X2=0 $Y2=0
cc_787 N_A_1518_203#_c_1145_n N_A_1266_74#_M1017_g 0.00301146f $X=9.105 $Y=1.855
+ $X2=0 $Y2=0
cc_788 N_A_1518_203#_c_1148_n N_A_1266_74#_M1017_g 0.00389282f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_789 N_A_1518_203#_c_1153_n N_A_1266_74#_c_1274_n 0.0107968f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_790 N_A_1518_203#_c_1154_n N_A_1266_74#_c_1274_n 0.00310966f $X=8.685 $Y=1.94
+ $X2=0 $Y2=0
cc_791 N_A_1518_203#_c_1145_n N_A_1266_74#_c_1274_n 0.00343619f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_792 N_A_1518_203#_c_1157_n N_A_1266_74#_c_1274_n 0.00678514f $X=8.502
+ $Y=2.445 $X2=0 $Y2=0
cc_793 N_A_1518_203#_c_1156_n N_A_1266_74#_c_1275_n 0.006945f $X=8.485 $Y=2.675
+ $X2=0 $Y2=0
cc_794 N_A_1518_203#_c_1157_n N_A_1266_74#_c_1275_n 0.00313845f $X=8.502
+ $Y=2.445 $X2=0 $Y2=0
cc_795 N_A_1518_203#_c_1153_n N_A_1266_74#_c_1261_n 0.00354772f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_796 N_A_1518_203#_c_1145_n N_A_1266_74#_c_1261_n 0.0103302f $X=9.105 $Y=1.855
+ $X2=0 $Y2=0
cc_797 N_A_1518_203#_c_1148_n N_A_1266_74#_c_1261_n 0.00508985f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_798 N_A_1518_203#_c_1154_n N_A_1266_74#_c_1262_n 7.74206e-19 $X=8.685 $Y=1.94
+ $X2=0 $Y2=0
cc_799 N_A_1518_203#_c_1148_n N_A_1266_74#_c_1262_n 8.2291e-19 $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_800 N_A_1518_203#_c_1145_n N_A_1266_74#_c_1263_n 0.00511666f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_801 N_A_1518_203#_c_1148_n N_A_1266_74#_c_1263_n 0.00147647f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_802 N_A_1518_203#_c_1153_n N_A_1266_74#_c_1278_n 6.47767e-19 $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_803 N_A_1518_203#_c_1145_n N_A_1266_74#_c_1278_n 0.00358035f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_804 N_A_1518_203#_c_1153_n N_A_1266_74#_c_1279_n 0.00455214f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_805 N_A_1518_203#_c_1157_n N_A_1266_74#_c_1279_n 9.14342e-19 $X=8.502
+ $Y=2.445 $X2=0 $Y2=0
cc_806 N_A_1518_203#_c_1144_n N_A_1266_74#_c_1265_n 2.88416e-19 $X=8.78 $Y=0.615
+ $X2=0 $Y2=0
cc_807 N_A_1518_203#_c_1148_n N_A_1266_74#_c_1265_n 0.00670166f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_808 N_A_1518_203#_c_1144_n N_A_1266_74#_c_1266_n 0.00317724f $X=8.78 $Y=0.615
+ $X2=0 $Y2=0
cc_809 N_A_1518_203#_c_1145_n N_A_1266_74#_c_1267_n 0.00419613f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_810 N_A_1518_203#_c_1151_n N_A_1266_74#_c_1303_n 0.00757243f $X=7.685 $Y=2.39
+ $X2=0 $Y2=0
cc_811 N_A_1518_203#_c_1149_n N_A_1266_74#_c_1282_n 0.00331106f $X=7.685
+ $Y=1.835 $X2=0 $Y2=0
cc_812 N_A_1518_203#_c_1150_n N_A_1266_74#_c_1282_n 0.0103166f $X=7.685 $Y=2.3
+ $X2=0 $Y2=0
cc_813 N_A_1518_203#_c_1151_n N_A_1266_74#_c_1282_n 0.0046186f $X=7.685 $Y=2.39
+ $X2=0 $Y2=0
cc_814 N_A_1518_203#_c_1142_n N_A_1266_74#_c_1282_n 0.0015543f $X=7.685 $Y=1.745
+ $X2=0 $Y2=0
cc_815 N_A_1518_203#_c_1149_n N_A_1266_74#_c_1270_n 8.26265e-19 $X=7.685
+ $Y=1.835 $X2=0 $Y2=0
cc_816 N_A_1518_203#_c_1142_n N_A_1266_74#_c_1270_n 0.00762694f $X=7.685
+ $Y=1.745 $X2=0 $Y2=0
cc_817 N_A_1518_203#_c_1143_n N_A_1266_74#_c_1270_n 0.0272699f $X=8.615 $Y=1.1
+ $X2=0 $Y2=0
cc_818 N_A_1518_203#_c_1154_n N_A_1266_74#_c_1270_n 4.22281e-19 $X=8.685 $Y=1.94
+ $X2=0 $Y2=0
cc_819 N_A_1518_203#_c_1146_n N_A_1266_74#_c_1270_n 0.0204811f $X=7.755 $Y=1.1
+ $X2=0 $Y2=0
cc_820 N_A_1518_203#_c_1147_n N_A_1266_74#_c_1270_n 0.00111936f $X=7.755 $Y=1.18
+ $X2=0 $Y2=0
cc_821 N_A_1518_203#_c_1142_n N_A_1266_74#_c_1271_n 0.00211774f $X=7.685
+ $Y=1.745 $X2=0 $Y2=0
cc_822 N_A_1518_203#_c_1146_n N_A_1266_74#_c_1271_n 0.0034757f $X=7.755 $Y=1.1
+ $X2=0 $Y2=0
cc_823 N_A_1518_203#_c_1143_n N_A_1266_74#_c_1273_n 0.0242574f $X=8.615 $Y=1.1
+ $X2=0 $Y2=0
cc_824 N_A_1518_203#_c_1153_n N_A_1266_74#_c_1273_n 0.0118853f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_825 N_A_1518_203#_c_1154_n N_A_1266_74#_c_1273_n 0.0136054f $X=8.685 $Y=1.94
+ $X2=0 $Y2=0
cc_826 N_A_1518_203#_c_1145_n N_A_1266_74#_c_1273_n 0.0235661f $X=9.105 $Y=1.855
+ $X2=0 $Y2=0
cc_827 N_A_1518_203#_c_1145_n N_A_1864_409#_c_1422_n 2.38456e-19 $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_828 N_A_1518_203#_c_1153_n N_A_1864_409#_c_1429_n 0.0121572f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_829 N_A_1518_203#_c_1145_n N_A_1864_409#_c_1429_n 0.00900265f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_830 N_A_1518_203#_c_1144_n N_A_1864_409#_c_1424_n 0.00478045f $X=8.78
+ $Y=0.615 $X2=0 $Y2=0
cc_831 N_A_1518_203#_c_1145_n N_A_1864_409#_c_1424_n 0.0077671f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_832 N_A_1518_203#_c_1148_n N_A_1864_409#_c_1424_n 0.00665068f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_833 N_A_1518_203#_c_1145_n N_A_1864_409#_c_1425_n 0.0234089f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_834 N_A_1518_203#_c_1151_n N_VPWR_c_1483_n 0.00654507f $X=7.685 $Y=2.39 $X2=0
+ $Y2=0
cc_835 N_A_1518_203#_c_1156_n N_VPWR_c_1483_n 0.0178695f $X=8.485 $Y=2.675 $X2=0
+ $Y2=0
cc_836 N_A_1518_203#_c_1156_n N_VPWR_c_1484_n 0.0120785f $X=8.485 $Y=2.675 $X2=0
+ $Y2=0
cc_837 N_A_1518_203#_c_1153_n N_VPWR_c_1485_n 0.0259196f $X=9.02 $Y=1.94 $X2=0
+ $Y2=0
cc_838 N_A_1518_203#_c_1157_n N_VPWR_c_1485_n 0.0548082f $X=8.502 $Y=2.445 $X2=0
+ $Y2=0
cc_839 N_A_1518_203#_c_1151_n N_VPWR_c_1491_n 0.00501877f $X=7.685 $Y=2.39 $X2=0
+ $Y2=0
cc_840 N_A_1518_203#_c_1151_n N_VPWR_c_1475_n 0.0052212f $X=7.685 $Y=2.39 $X2=0
+ $Y2=0
cc_841 N_A_1518_203#_c_1156_n N_VPWR_c_1475_n 0.0126247f $X=8.485 $Y=2.675 $X2=0
+ $Y2=0
cc_842 N_A_1518_203#_M1014_g N_VGND_c_1793_n 0.0107187f $X=7.695 $Y=0.615 $X2=0
+ $Y2=0
cc_843 N_A_1518_203#_c_1143_n N_VGND_c_1793_n 0.0130069f $X=8.615 $Y=1.1 $X2=0
+ $Y2=0
cc_844 N_A_1518_203#_c_1144_n N_VGND_c_1793_n 0.00738736f $X=8.78 $Y=0.615 $X2=0
+ $Y2=0
cc_845 N_A_1518_203#_c_1146_n N_VGND_c_1793_n 0.0145528f $X=7.755 $Y=1.1 $X2=0
+ $Y2=0
cc_846 N_A_1518_203#_c_1147_n N_VGND_c_1793_n 0.0011793f $X=7.755 $Y=1.18 $X2=0
+ $Y2=0
cc_847 N_A_1518_203#_c_1144_n N_VGND_c_1794_n 0.0303742f $X=8.78 $Y=0.615 $X2=0
+ $Y2=0
cc_848 N_A_1518_203#_c_1148_n N_VGND_c_1794_n 0.00112954f $X=9.105 $Y=1.1 $X2=0
+ $Y2=0
cc_849 N_A_1518_203#_M1014_g N_VGND_c_1801_n 0.0045897f $X=7.695 $Y=0.615 $X2=0
+ $Y2=0
cc_850 N_A_1518_203#_c_1144_n N_VGND_c_1802_n 0.0126905f $X=8.78 $Y=0.615 $X2=0
+ $Y2=0
cc_851 N_A_1518_203#_M1014_g N_VGND_c_1807_n 0.0044912f $X=7.695 $Y=0.615 $X2=0
+ $Y2=0
cc_852 N_A_1518_203#_c_1144_n N_VGND_c_1807_n 0.0118012f $X=8.78 $Y=0.615 $X2=0
+ $Y2=0
cc_853 N_A_1266_74#_c_1264_n N_A_1864_409#_c_1422_n 0.00139534f $X=9.48 $Y=1.07
+ $X2=0 $Y2=0
cc_854 N_A_1266_74#_c_1267_n N_A_1864_409#_c_1422_n 0.0154815f $X=9.245 $Y=1.52
+ $X2=0 $Y2=0
cc_855 N_A_1266_74#_c_1278_n N_A_1864_409#_c_1429_n 0.00590965f $X=9.245 $Y=1.88
+ $X2=0 $Y2=0
cc_856 N_A_1266_74#_c_1279_n N_A_1864_409#_c_1429_n 0.0105256f $X=9.245 $Y=1.97
+ $X2=0 $Y2=0
cc_857 N_A_1266_74#_c_1263_n N_A_1864_409#_c_1424_n 0.00400367f $X=9.23 $Y=1.355
+ $X2=0 $Y2=0
cc_858 N_A_1266_74#_c_1264_n N_A_1864_409#_c_1424_n 0.00708838f $X=9.48 $Y=1.07
+ $X2=0 $Y2=0
cc_859 N_A_1266_74#_c_1266_n N_A_1864_409#_c_1424_n 0.0140899f $X=9.555 $Y=0.995
+ $X2=0 $Y2=0
cc_860 N_A_1266_74#_c_1267_n N_A_1864_409#_c_1424_n 7.91947e-19 $X=9.245 $Y=1.52
+ $X2=0 $Y2=0
cc_861 N_A_1266_74#_c_1264_n N_A_1864_409#_c_1425_n 0.0079216f $X=9.48 $Y=1.07
+ $X2=0 $Y2=0
cc_862 N_A_1266_74#_c_1267_n N_A_1864_409#_c_1425_n 0.00324958f $X=9.245 $Y=1.52
+ $X2=0 $Y2=0
cc_863 N_A_1266_74#_c_1282_n N_VPWR_c_1483_n 0.00177331f $X=7.55 $Y=2.475 $X2=0
+ $Y2=0
cc_864 N_A_1266_74#_c_1275_n N_VPWR_c_1484_n 0.00477303f $X=8.71 $Y=2.39 $X2=0
+ $Y2=0
cc_865 N_A_1266_74#_c_1274_n N_VPWR_c_1485_n 0.001714f $X=8.71 $Y=2.3 $X2=0
+ $Y2=0
cc_866 N_A_1266_74#_c_1275_n N_VPWR_c_1485_n 0.00744434f $X=8.71 $Y=2.39 $X2=0
+ $Y2=0
cc_867 N_A_1266_74#_c_1261_n N_VPWR_c_1485_n 3.97376e-19 $X=9.155 $Y=1.52 $X2=0
+ $Y2=0
cc_868 N_A_1266_74#_c_1279_n N_VPWR_c_1485_n 0.0126982f $X=9.245 $Y=1.97 $X2=0
+ $Y2=0
cc_869 N_A_1266_74#_c_1303_n N_VPWR_c_1491_n 0.0213832f $X=7.465 $Y=2.64 $X2=0
+ $Y2=0
cc_870 N_A_1266_74#_c_1404_p N_VPWR_c_1491_n 0.00379401f $X=6.65 $Y=2.64 $X2=0
+ $Y2=0
cc_871 N_A_1266_74#_c_1279_n N_VPWR_c_1492_n 0.00470366f $X=9.245 $Y=1.97 $X2=0
+ $Y2=0
cc_872 N_A_1266_74#_c_1275_n N_VPWR_c_1475_n 0.0052212f $X=8.71 $Y=2.39 $X2=0
+ $Y2=0
cc_873 N_A_1266_74#_c_1279_n N_VPWR_c_1475_n 0.00473388f $X=9.245 $Y=1.97 $X2=0
+ $Y2=0
cc_874 N_A_1266_74#_c_1303_n N_VPWR_c_1475_n 0.0313462f $X=7.465 $Y=2.64 $X2=0
+ $Y2=0
cc_875 N_A_1266_74#_c_1404_p N_VPWR_c_1475_n 0.00557315f $X=6.65 $Y=2.64 $X2=0
+ $Y2=0
cc_876 N_A_1266_74#_c_1303_n A_1468_493# 0.00358233f $X=7.465 $Y=2.64 $X2=-0.19
+ $Y2=-0.245
cc_877 N_A_1266_74#_c_1266_n N_Q_c_1761_n 0.00112501f $X=9.555 $Y=0.995 $X2=0
+ $Y2=0
cc_878 N_A_1266_74#_c_1264_n N_Q_c_1762_n 0.00112501f $X=9.48 $Y=1.07 $X2=0
+ $Y2=0
cc_879 N_A_1266_74#_c_1279_n Q 0.00322019f $X=9.245 $Y=1.97 $X2=0 $Y2=0
cc_880 N_A_1266_74#_M1017_g N_VGND_c_1794_n 0.00359522f $X=8.565 $Y=0.615 $X2=0
+ $Y2=0
cc_881 N_A_1266_74#_c_1265_n N_VGND_c_1794_n 0.0104251f $X=9.305 $Y=1.07 $X2=0
+ $Y2=0
cc_882 N_A_1266_74#_c_1266_n N_VGND_c_1794_n 0.0065091f $X=9.555 $Y=0.995 $X2=0
+ $Y2=0
cc_883 N_A_1266_74#_M1017_g N_VGND_c_1802_n 0.00527282f $X=8.565 $Y=0.615 $X2=0
+ $Y2=0
cc_884 N_A_1266_74#_c_1266_n N_VGND_c_1803_n 0.00434272f $X=9.555 $Y=0.995 $X2=0
+ $Y2=0
cc_885 N_A_1266_74#_M1017_g N_VGND_c_1807_n 0.00534666f $X=8.565 $Y=0.615 $X2=0
+ $Y2=0
cc_886 N_A_1266_74#_c_1266_n N_VGND_c_1807_n 0.00830282f $X=9.555 $Y=0.995 $X2=0
+ $Y2=0
cc_887 N_A_1864_409#_c_1429_n N_VPWR_c_1485_n 0.0462745f $X=9.47 $Y=2.19 $X2=0
+ $Y2=0
cc_888 N_A_1864_409#_c_1426_n N_VPWR_c_1487_n 0.0203918f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_889 N_A_1864_409#_c_1423_n N_VPWR_c_1487_n 8.22785e-19 $X=10.53 $Y=1.575
+ $X2=0 $Y2=0
cc_890 N_A_1864_409#_c_1426_n N_VPWR_c_1492_n 0.00429299f $X=10.53 $Y=1.765
+ $X2=0 $Y2=0
cc_891 N_A_1864_409#_c_1429_n N_VPWR_c_1492_n 0.00575213f $X=9.47 $Y=2.19 $X2=0
+ $Y2=0
cc_892 N_A_1864_409#_c_1426_n N_VPWR_c_1475_n 0.00852523f $X=10.53 $Y=1.765
+ $X2=0 $Y2=0
cc_893 N_A_1864_409#_c_1429_n N_VPWR_c_1475_n 0.00591657f $X=9.47 $Y=2.19 $X2=0
+ $Y2=0
cc_894 N_A_1864_409#_M1002_g N_Q_c_1761_n 0.00853833f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_895 N_A_1864_409#_c_1424_n N_Q_c_1761_n 0.0694074f $X=9.77 $Y=0.645 $X2=0
+ $Y2=0
cc_896 N_A_1864_409#_M1002_g N_Q_c_1762_n 0.00343176f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_897 N_A_1864_409#_c_1422_n N_Q_c_1762_n 0.00187014f $X=10.44 $Y=1.55 $X2=0
+ $Y2=0
cc_898 N_A_1864_409#_c_1422_n Q 0.0150903f $X=10.44 $Y=1.55 $X2=0 $Y2=0
cc_899 N_A_1864_409#_c_1429_n Q 0.0848083f $X=9.47 $Y=2.19 $X2=0 $Y2=0
cc_900 N_A_1864_409#_c_1425_n Q 0.017588f $X=9.77 $Y=1.55 $X2=0 $Y2=0
cc_901 N_A_1864_409#_c_1426_n N_Q_c_1763_n 0.00351033f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_902 N_A_1864_409#_M1002_g N_Q_c_1763_n 0.0104864f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_903 N_A_1864_409#_c_1422_n N_Q_c_1763_n 0.0395686f $X=10.44 $Y=1.55 $X2=0
+ $Y2=0
cc_904 N_A_1864_409#_c_1423_n N_Q_c_1763_n 0.00217631f $X=10.53 $Y=1.575 $X2=0
+ $Y2=0
cc_905 N_A_1864_409#_c_1429_n N_Q_c_1763_n 0.00535008f $X=9.47 $Y=2.19 $X2=0
+ $Y2=0
cc_906 N_A_1864_409#_c_1425_n N_Q_c_1763_n 0.0198451f $X=9.77 $Y=1.55 $X2=0
+ $Y2=0
cc_907 N_A_1864_409#_c_1424_n N_VGND_c_1794_n 0.0184694f $X=9.77 $Y=0.645 $X2=0
+ $Y2=0
cc_908 N_A_1864_409#_c_1425_n N_VGND_c_1794_n 0.00144181f $X=9.77 $Y=1.55 $X2=0
+ $Y2=0
cc_909 N_A_1864_409#_M1002_g N_VGND_c_1796_n 0.00647412f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_910 N_A_1864_409#_M1002_g N_VGND_c_1803_n 0.00434272f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_911 N_A_1864_409#_c_1424_n N_VGND_c_1803_n 0.0145639f $X=9.77 $Y=0.645 $X2=0
+ $Y2=0
cc_912 N_A_1864_409#_M1002_g N_VGND_c_1807_n 0.00828941f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_913 N_A_1864_409#_c_1424_n N_VGND_c_1807_n 0.0119984f $X=9.77 $Y=0.645 $X2=0
+ $Y2=0
cc_914 N_VPWR_c_1477_n N_A_30_78#_c_1631_n 0.0223613f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_915 N_VPWR_c_1478_n N_A_30_78#_c_1631_n 0.0101408f $X=1.145 $Y=2.815 $X2=0
+ $Y2=0
cc_916 N_VPWR_c_1488_n N_A_30_78#_c_1631_n 0.0110897f $X=0.98 $Y=3.33 $X2=0
+ $Y2=0
cc_917 N_VPWR_c_1475_n N_A_30_78#_c_1631_n 0.0092154f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_918 N_VPWR_M1000_d N_A_30_78#_c_1633_n 0.00225122f $X=1.005 $Y=2.54 $X2=0
+ $Y2=0
cc_919 N_VPWR_c_1478_n N_A_30_78#_c_1633_n 0.0213601f $X=1.145 $Y=2.815 $X2=0
+ $Y2=0
cc_920 N_VPWR_c_1489_n N_A_30_78#_c_1633_n 0.00196088f $X=1.985 $Y=3.33 $X2=0
+ $Y2=0
cc_921 N_VPWR_c_1475_n N_A_30_78#_c_1633_n 0.0119186f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_922 N_VPWR_c_1489_n N_A_30_78#_c_1634_n 0.00530811f $X=1.985 $Y=3.33 $X2=0
+ $Y2=0
cc_923 N_VPWR_c_1475_n N_A_30_78#_c_1634_n 0.0105073f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_924 N_VPWR_M1006_d N_A_30_78#_c_1635_n 0.00511413f $X=2 $Y=1.95 $X2=0 $Y2=0
cc_925 N_VPWR_c_1479_n N_A_30_78#_c_1635_n 0.0168112f $X=2.15 $Y=2.825 $X2=0
+ $Y2=0
cc_926 N_VPWR_c_1489_n N_A_30_78#_c_1635_n 7.38795e-19 $X=1.985 $Y=3.33 $X2=0
+ $Y2=0
cc_927 N_VPWR_c_1490_n N_A_30_78#_c_1635_n 0.00886008f $X=4.385 $Y=3.33 $X2=0
+ $Y2=0
cc_928 N_VPWR_c_1475_n N_A_30_78#_c_1635_n 0.01976f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_929 N_VPWR_c_1477_n N_A_30_78#_c_1638_n 0.00821798f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_930 N_VPWR_c_1488_n N_A_30_78#_c_1638_n 2.18842e-19 $X=0.98 $Y=3.33 $X2=0
+ $Y2=0
cc_931 N_VPWR_c_1475_n N_A_30_78#_c_1638_n 0.00139524f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_932 N_VPWR_c_1490_n N_A_30_78#_c_1639_n 0.00592793f $X=4.385 $Y=3.33 $X2=0
+ $Y2=0
cc_933 N_VPWR_c_1475_n N_A_30_78#_c_1639_n 0.00748882f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_934 N_VPWR_c_1485_n Q 0.00265735f $X=9.02 $Y=2.36 $X2=0 $Y2=0
cc_935 N_VPWR_c_1492_n Q 0.0311454f $X=10.595 $Y=3.33 $X2=0 $Y2=0
cc_936 N_VPWR_c_1475_n Q 0.0257795f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_937 N_VPWR_c_1487_n N_Q_c_1763_n 0.045174f $X=10.76 $Y=1.985 $X2=0 $Y2=0
cc_938 N_A_30_78#_c_1624_n A_117_78# 0.00231141f $X=0.685 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_939 N_A_30_78#_c_1624_n N_VGND_c_1791_n 0.00719261f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_940 N_A_30_78#_c_1628_n N_VGND_c_1791_n 0.00436551f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_941 N_A_30_78#_c_1624_n N_VGND_c_1797_n 0.00570266f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_942 N_A_30_78#_c_1628_n N_VGND_c_1797_n 0.0131067f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_943 N_A_30_78#_c_1624_n N_VGND_c_1807_n 0.0110739f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_944 N_A_30_78#_c_1628_n N_VGND_c_1807_n 0.0117869f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_945 N_Q_c_1761_n N_VGND_c_1796_n 0.0293763f $X=10.33 $Y=0.515 $X2=0 $Y2=0
cc_946 N_Q_c_1761_n N_VGND_c_1803_n 0.0145639f $X=10.33 $Y=0.515 $X2=0 $Y2=0
cc_947 N_Q_c_1761_n N_VGND_c_1807_n 0.0119984f $X=10.33 $Y=0.515 $X2=0 $Y2=0
