* File: sky130_fd_sc_ls__a211o_2.pex.spice
* Created: Fri Aug 28 12:49:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A211O_2%A_85_270# 1 2 3 11 12 14 17 19 21 24 29 30
+ 31 32 33 36 38 40 42 46 49 51 53 59
c128 49 0 2.02221e-19 $X=1.17 $Y=1.515
c129 24 0 9.24433e-20 $X=1.11 $Y=0.74
r130 58 59 27.1946 $w=2.57e-07 $l=1.45e-07 $layer=POLY_cond $X=0.965 $Y=1.557
+ $X2=1.11 $Y2=1.557
r131 50 59 11.2529 $w=2.57e-07 $l=6e-08 $layer=POLY_cond $X=1.17 $Y=1.557
+ $X2=1.11 $Y2=1.557
r132 49 52 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.17 $Y=1.515
+ $X2=1.17 $Y2=1.68
r133 49 51 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.17 $Y=1.515
+ $X2=1.17 $Y2=1.35
r134 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.515 $X2=1.17 $Y2=1.515
r135 44 46 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=3.615 $Y=0.92
+ $X2=3.615 $Y2=0.515
r136 40 55 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=2.12 $X2=3.57
+ $Y2=2.035
r137 40 42 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.57 $Y=2.12
+ $X2=3.57 $Y2=2.815
r138 39 53 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.7 $Y=1.005
+ $X2=2.515 $Y2=1.005
r139 38 44 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.49 $Y=1.005
+ $X2=3.615 $Y2=0.92
r140 38 39 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.49 $Y=1.005
+ $X2=2.7 $Y2=1.005
r141 34 53 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=0.92
+ $X2=2.515 $Y2=1.005
r142 34 36 12.6146 $w=3.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.515 $Y=0.92
+ $X2=2.515 $Y2=0.515
r143 32 55 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=2.035
+ $X2=3.57 $Y2=2.035
r144 32 33 135.048 $w=1.68e-07 $l=2.07e-06 $layer=LI1_cond $X=3.405 $Y=2.035
+ $X2=1.335 $Y2=2.035
r145 30 53 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.33 $Y=1.005
+ $X2=2.515 $Y2=1.005
r146 30 31 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=2.33 $Y=1.005
+ $X2=1.335 $Y2=1.005
r147 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.25 $Y=1.95
+ $X2=1.335 $Y2=2.035
r148 29 52 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.25 $Y=1.95
+ $X2=1.25 $Y2=1.68
r149 26 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.25 $Y=1.09
+ $X2=1.335 $Y2=1.005
r150 26 51 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.25 $Y=1.09
+ $X2=1.25 $Y2=1.35
r151 22 59 15.359 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.11 $Y=1.35
+ $X2=1.11 $Y2=1.557
r152 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.11 $Y=1.35
+ $X2=1.11 $Y2=0.74
r153 19 58 15.359 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.765
+ $X2=0.965 $Y2=1.557
r154 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.965 $Y=1.765
+ $X2=0.965 $Y2=2.4
r155 15 58 53.4514 $w=2.57e-07 $l=3.7446e-07 $layer=POLY_cond $X=0.68 $Y=1.35
+ $X2=0.965 $Y2=1.557
r156 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.68 $Y=1.35
+ $X2=0.68 $Y2=0.74
r157 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.515 $Y=1.765
+ $X2=0.515 $Y2=2.4
r158 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.515 $Y=1.675
+ $X2=0.515 $Y2=1.765
r159 10 15 30.9455 $w=2.57e-07 $l=2.2798e-07 $layer=POLY_cond $X=0.515 $Y=1.5
+ $X2=0.68 $Y2=1.35
r160 10 11 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=0.515 $Y=1.5
+ $X2=0.515 $Y2=1.675
r161 3 55 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.96 $X2=3.57 $Y2=2.115
r162 3 42 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.96 $X2=3.57 $Y2=2.815
r163 2 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.435
+ $Y=0.37 $X2=3.575 $Y2=0.515
r164 1 36 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=2.355
+ $Y=0.37 $X2=2.515 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_2%A2 3 7 9 10 11 15 17
c44 15 0 2.19694e-19 $X=1.71 $Y=1.425
c45 10 0 7.65662e-20 $X=1.935 $Y=1.73
r46 14 17 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.71 $Y=1.425
+ $X2=1.92 $Y2=1.425
r47 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.425 $X2=1.71 $Y2=1.425
r48 11 15 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.425
r49 7 10 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=1.935 $Y=1.885
+ $X2=1.935 $Y2=1.73
r50 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.935 $Y=1.885
+ $X2=1.935 $Y2=2.46
r51 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.59
+ $X2=1.92 $Y2=1.425
r52 5 10 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=1.92 $Y=1.59 $X2=1.92
+ $Y2=1.73
r53 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.26
+ $X2=1.92 $Y2=1.425
r54 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.92 $Y=1.26 $X2=1.92
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_2%A1 3 7 9 10 11 14 15
c46 10 0 1.27251e-19 $X=2.475 $Y=1.73
c47 3 0 1.02299e-19 $X=2.28 $Y=0.74
r48 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.37 $Y=1.425
+ $X2=2.37 $Y2=1.59
r49 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.37 $Y=1.425
+ $X2=2.37 $Y2=1.26
r50 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.37
+ $Y=1.425 $X2=2.37 $Y2=1.425
r51 11 15 5.85834 $w=4.88e-07 $l=2.4e-07 $layer=LI1_cond $X=2.29 $Y=1.665
+ $X2=2.29 $Y2=1.425
r52 10 17 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.46 $Y=1.73
+ $X2=2.46 $Y2=1.59
r53 7 10 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=2.475 $Y=1.885
+ $X2=2.475 $Y2=1.73
r54 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.475 $Y=1.885
+ $X2=2.475 $Y2=2.46
r55 3 16 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.28 $Y=0.74 $X2=2.28
+ $Y2=1.26
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_2%B1 3 6 7 9 10 13 14
c40 13 0 1.08088e-19 $X=2.91 $Y=1.425
c41 6 0 1.39721e-19 $X=2.925 $Y=1.795
r42 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.91 $Y=1.425
+ $X2=2.91 $Y2=1.59
r43 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.91 $Y=1.425
+ $X2=2.91 $Y2=1.26
r44 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.91
+ $Y=1.425 $X2=2.91 $Y2=1.425
r45 10 14 5.85834 $w=4.88e-07 $l=2.4e-07 $layer=LI1_cond $X=2.99 $Y=1.665
+ $X2=2.99 $Y2=1.425
r46 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.925 $Y=1.885
+ $X2=2.925 $Y2=2.46
r47 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.925 $Y=1.795 $X2=2.925
+ $Y2=1.885
r48 6 16 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=2.925 $Y=1.795
+ $X2=2.925 $Y2=1.59
r49 3 15 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.82 $Y=0.74 $X2=2.82
+ $Y2=1.26
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_2%C1 1 3 6 8
c27 8 0 2.47809e-19 $X=3.6 $Y=1.665
r28 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.615 $X2=3.57 $Y2=1.615
r29 4 11 39.3587 $w=3.88e-07 $l=2.22486e-07 $layer=POLY_cond $X=3.36 $Y=1.45
+ $X2=3.495 $Y2=1.615
r30 4 6 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.36 $Y=1.45 $X2=3.36
+ $Y2=0.74
r31 1 11 52.4025 $w=3.88e-07 $l=3.36749e-07 $layer=POLY_cond $X=3.345 $Y=1.885
+ $X2=3.495 $Y2=1.615
r32 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.345 $Y=1.885
+ $X2=3.345 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_2%VPWR 1 2 3 10 12 18 22 24 26 31 41 42 48 51
r51 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r53 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r55 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r56 39 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 38 41 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r58 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 36 51 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.22 $Y2=3.33
r60 36 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r62 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 32 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=3.33
+ $X2=1.19 $Y2=3.33
r64 32 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.355 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 31 51 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.075 $Y=3.33
+ $X2=2.22 $Y2=3.33
r66 31 34 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.075 $Y=3.33
+ $X2=1.68 $Y2=3.33
r67 30 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 30 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r69 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r70 27 45 3.99677 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=3.33
+ $X2=0.187 $Y2=3.33
r71 27 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.375 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 26 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=1.19 $Y2=3.33
r73 26 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=0.72 $Y2=3.33
r74 24 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r75 24 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r76 20 51 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=3.245
+ $X2=2.22 $Y2=3.33
r77 20 22 17.4853 $w=2.88e-07 $l=4.4e-07 $layer=LI1_cond $X=2.22 $Y=3.245
+ $X2=2.22 $Y2=2.805
r78 16 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=3.33
r79 16 18 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=2.455
r80 12 15 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.25 $Y=1.985
+ $X2=0.25 $Y2=2.815
r81 10 45 3.14639 $w=2.5e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.25 $Y=3.245
+ $X2=0.187 $Y2=3.33
r82 10 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.25 $Y=3.245
+ $X2=0.25 $Y2=2.815
r83 3 22 600 $w=1.7e-07 $l=9.26107e-07 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.96 $X2=2.18 $Y2=2.805
r84 2 18 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=1.84 $X2=1.19 $Y2=2.455
r85 1 15 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.84 $X2=0.29 $Y2=2.815
r86 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.84 $X2=0.29 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_2%X 1 2 9 14 16 17 18 19 20
r28 19 20 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=2.405
+ $X2=0.705 $Y2=2.775
r29 18 19 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=0.705 $Y=1.985
+ $X2=0.705 $Y2=2.405
r30 17 18 14.1839 $w=2.58e-07 $l=3.2e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.985
r31 16 17 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=1.295
+ $X2=0.705 $Y2=1.665
r32 12 16 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=0.705 $Y=1.18
+ $X2=0.705 $Y2=1.295
r33 12 14 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.705 $Y=1.095
+ $X2=0.895 $Y2=1.095
r34 7 14 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=1.01
+ $X2=0.895 $Y2=1.095
r35 7 9 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=0.895 $Y=1.01
+ $X2=0.895 $Y2=0.515
r36 2 20 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.84 $X2=0.74 $Y2=2.815
r37 2 18 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.84 $X2=0.74 $Y2=1.985
r38 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.755
+ $Y=0.37 $X2=0.895 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_2%A_317_392# 1 2 9 14 16
r26 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=2.375
+ $X2=1.71 $Y2=2.375
r27 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=2.375
+ $X2=2.7 $Y2=2.375
r28 9 10 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.535 $Y=2.375
+ $X2=1.875 $Y2=2.375
r29 2 16 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=2.55
+ $Y=1.96 $X2=2.7 $Y2=2.455
r30 1 14 300 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=2 $X=1.585
+ $Y=1.96 $X2=1.71 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__A211O_2%VGND 1 2 3 12 14 17 18 20 23 24 25 27 28 32
+ 34 47 48 51
c60 32 0 1.02299e-19 $X=3.09 $Y=0.55
c61 18 0 1.25655e-19 $X=1.33 $Y=0.55
r62 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r63 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r64 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r65 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r66 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r67 41 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r68 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r69 39 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.33 $Y=0 $X2=1.245
+ $Y2=0
r70 39 41 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.33 $Y=0 $X2=1.68
+ $Y2=0
r71 38 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r72 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r73 34 45 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r74 34 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r75 29 32 3.8895 $w=3.98e-07 $l=1.35e-07 $layer=LI1_cond $X=2.955 $Y=0.55
+ $X2=3.09 $Y2=0.55
r76 27 44 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=2.64
+ $Y2=0
r77 27 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=0 $X2=2.955
+ $Y2=0
r78 26 47 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=3.6
+ $Y2=0
r79 26 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=0 $X2=2.955
+ $Y2=0
r80 24 37 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=0.3 $Y=0 $X2=0.24 $Y2=0
r81 24 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.3 $Y=0 $X2=0.465
+ $Y2=0
r82 23 29 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.955 $Y=0.35 $X2=2.955
+ $Y2=0.55
r83 22 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=0.085
+ $X2=2.955 $Y2=0
r84 22 23 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.955 $Y=0.085
+ $X2=2.955 $Y2=0.35
r85 18 20 10.8042 $w=3.98e-07 $l=3.75e-07 $layer=LI1_cond $X=1.33 $Y=0.55
+ $X2=1.705 $Y2=0.55
r86 17 18 8.37092 $w=4e-07 $l=2.38747e-07 $layer=LI1_cond $X=1.245 $Y=0.35
+ $X2=1.33 $Y2=0.55
r87 16 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0
r88 16 17 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0.35
r89 15 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.465
+ $Y2=0
r90 14 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=0 $X2=1.245
+ $Y2=0
r91 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.16 $Y=0 $X2=0.63
+ $Y2=0
r92 10 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.465 $Y=0.085
+ $X2=0.465 $Y2=0
r93 10 12 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.465 $Y=0.085
+ $X2=0.465 $Y2=0.595
r94 3 32 182 $w=1.7e-07 $l=2.70416e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.37 $X2=3.09 $Y2=0.55
r95 2 20 91 $w=1.7e-07 $l=6.03324e-07 $layer=licon1_NDIFF $count=2 $X=1.185
+ $Y=0.37 $X2=1.705 $Y2=0.55
r96 1 12 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.34
+ $Y=0.37 $X2=0.465 $Y2=0.595
.ends

