* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_31_368# a_803_323# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VPWR B1_N a_803_323# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 a_31_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 a_31_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X4 a_46_74# A1 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 VGND A2 a_46_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 a_46_74# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 a_31_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 VGND A2 a_46_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 VGND a_803_323# Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X10 a_31_368# a_803_323# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 Y a_803_323# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 a_803_323# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 VGND a_803_323# Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X14 VGND B1_N a_803_323# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 a_31_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X16 Y A1 a_46_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 Y a_803_323# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 VPWR A2 a_31_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X19 Y a_803_323# a_31_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X20 a_46_74# A1 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 VPWR A2 a_31_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X22 VPWR A1 a_31_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X23 VPWR A1 a_31_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X24 Y A1 a_46_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X25 a_46_74# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X26 Y a_803_323# a_31_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
.ends
