* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_507_368# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VGND A1 a_225_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 a_225_74# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_225_74# a_27_74# Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 VPWR a_27_74# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X5 Y a_27_74# a_225_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 Y A2 a_507_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 VPWR A1 a_507_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 Y a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 VGND A2 a_225_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X10 a_225_74# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X11 a_27_74# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_27_74# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_507_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
.ends
