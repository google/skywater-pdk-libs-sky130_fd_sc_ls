* File: sky130_fd_sc_ls__dlrtp_2.pxi.spice
* Created: Fri Aug 28 13:19:17 2020
* 
x_PM_SKY130_FD_SC_LS__DLRTP_2%D N_D_c_139_n N_D_M1012_g N_D_M1006_g D
+ N_D_c_141_n PM_SKY130_FD_SC_LS__DLRTP_2%D
x_PM_SKY130_FD_SC_LS__DLRTP_2%GATE N_GATE_M1019_g N_GATE_c_167_n N_GATE_c_172_n
+ N_GATE_M1009_g GATE N_GATE_c_169_n N_GATE_c_170_n
+ PM_SKY130_FD_SC_LS__DLRTP_2%GATE
x_PM_SKY130_FD_SC_LS__DLRTP_2%A_235_74# N_A_235_74#_M1019_d N_A_235_74#_M1009_d
+ N_A_235_74#_c_210_n N_A_235_74#_M1017_g N_A_235_74#_M1021_g
+ N_A_235_74#_c_226_n N_A_235_74#_M1008_g N_A_235_74#_c_212_n
+ N_A_235_74#_c_213_n N_A_235_74#_M1015_g N_A_235_74#_c_215_n
+ N_A_235_74#_c_216_n N_A_235_74#_c_230_n N_A_235_74#_c_217_n
+ N_A_235_74#_c_257_p N_A_235_74#_c_218_n N_A_235_74#_c_219_n
+ N_A_235_74#_c_220_n N_A_235_74#_c_231_n N_A_235_74#_c_221_n
+ N_A_235_74#_c_222_n N_A_235_74#_c_223_n N_A_235_74#_c_224_n
+ PM_SKY130_FD_SC_LS__DLRTP_2%A_235_74#
x_PM_SKY130_FD_SC_LS__DLRTP_2%A_27_392# N_A_27_392#_M1006_s N_A_27_392#_M1012_s
+ N_A_27_392#_c_361_n N_A_27_392#_M1010_g N_A_27_392#_M1000_g
+ N_A_27_392#_c_363_n N_A_27_392#_c_364_n N_A_27_392#_c_365_n
+ N_A_27_392#_c_366_n N_A_27_392#_c_370_n N_A_27_392#_c_371_n
+ N_A_27_392#_c_372_n N_A_27_392#_c_367_n PM_SKY130_FD_SC_LS__DLRTP_2%A_27_392#
x_PM_SKY130_FD_SC_LS__DLRTP_2%A_347_98# N_A_347_98#_M1021_s N_A_347_98#_M1017_s
+ N_A_347_98#_M1001_g N_A_347_98#_c_464_n N_A_347_98#_M1018_g
+ N_A_347_98#_c_458_n N_A_347_98#_c_459_n N_A_347_98#_c_516_n
+ N_A_347_98#_c_460_n N_A_347_98#_c_467_n N_A_347_98#_c_468_n
+ N_A_347_98#_c_469_n N_A_347_98#_c_461_n N_A_347_98#_c_470_n
+ N_A_347_98#_c_471_n N_A_347_98#_c_462_n N_A_347_98#_c_463_n
+ N_A_347_98#_c_472_n PM_SKY130_FD_SC_LS__DLRTP_2%A_347_98#
x_PM_SKY130_FD_SC_LS__DLRTP_2%A_832_55# N_A_832_55#_M1011_s N_A_832_55#_M1007_d
+ N_A_832_55#_c_573_n N_A_832_55#_M1016_g N_A_832_55#_c_574_n
+ N_A_832_55#_c_584_n N_A_832_55#_M1005_g N_A_832_55#_c_585_n
+ N_A_832_55#_M1002_g N_A_832_55#_M1004_g N_A_832_55#_M1013_g
+ N_A_832_55#_c_586_n N_A_832_55#_M1020_g N_A_832_55#_c_577_n
+ N_A_832_55#_c_587_n N_A_832_55#_c_578_n N_A_832_55#_c_588_n
+ N_A_832_55#_c_589_n N_A_832_55#_c_579_n N_A_832_55#_c_670_p
+ N_A_832_55#_c_580_n N_A_832_55#_c_591_n N_A_832_55#_c_581_n
+ N_A_832_55#_c_582_n PM_SKY130_FD_SC_LS__DLRTP_2%A_832_55#
x_PM_SKY130_FD_SC_LS__DLRTP_2%A_646_74# N_A_646_74#_M1001_d N_A_646_74#_M1008_d
+ N_A_646_74#_c_710_n N_A_646_74#_M1007_g N_A_646_74#_M1011_g
+ N_A_646_74#_c_705_n N_A_646_74#_c_706_n N_A_646_74#_c_707_n
+ N_A_646_74#_c_708_n N_A_646_74#_c_713_n N_A_646_74#_c_709_n
+ N_A_646_74#_c_715_n N_A_646_74#_c_716_n N_A_646_74#_c_717_n
+ PM_SKY130_FD_SC_LS__DLRTP_2%A_646_74#
x_PM_SKY130_FD_SC_LS__DLRTP_2%RESET_B N_RESET_B_c_793_n N_RESET_B_M1003_g
+ N_RESET_B_c_794_n N_RESET_B_M1014_g RESET_B N_RESET_B_c_795_n
+ PM_SKY130_FD_SC_LS__DLRTP_2%RESET_B
x_PM_SKY130_FD_SC_LS__DLRTP_2%VPWR N_VPWR_M1012_d N_VPWR_M1017_d N_VPWR_M1005_d
+ N_VPWR_M1014_d N_VPWR_M1020_s N_VPWR_c_829_n N_VPWR_c_830_n N_VPWR_c_831_n
+ N_VPWR_c_832_n N_VPWR_c_833_n N_VPWR_c_834_n N_VPWR_c_835_n VPWR
+ N_VPWR_c_836_n N_VPWR_c_837_n N_VPWR_c_838_n N_VPWR_c_839_n N_VPWR_c_840_n
+ N_VPWR_c_841_n N_VPWR_c_828_n PM_SKY130_FD_SC_LS__DLRTP_2%VPWR
x_PM_SKY130_FD_SC_LS__DLRTP_2%Q N_Q_M1004_d N_Q_M1002_d N_Q_c_917_n N_Q_c_921_n
+ N_Q_c_922_n N_Q_c_918_n N_Q_c_919_n N_Q_c_923_n Q
+ PM_SKY130_FD_SC_LS__DLRTP_2%Q
x_PM_SKY130_FD_SC_LS__DLRTP_2%VGND N_VGND_M1006_d N_VGND_M1021_d N_VGND_M1016_d
+ N_VGND_M1003_d N_VGND_M1013_s N_VGND_c_961_n N_VGND_c_962_n N_VGND_c_963_n
+ N_VGND_c_964_n N_VGND_c_965_n N_VGND_c_966_n N_VGND_c_967_n VGND
+ N_VGND_c_968_n N_VGND_c_969_n N_VGND_c_970_n N_VGND_c_971_n N_VGND_c_972_n
+ N_VGND_c_973_n N_VGND_c_974_n PM_SKY130_FD_SC_LS__DLRTP_2%VGND
cc_1 VNB N_D_c_139_n 0.0248281f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_2 VNB N_D_M1006_g 0.0403394f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.835
cc_3 VNB N_D_c_141_n 0.00925599f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_4 VNB N_GATE_c_167_n 0.00704352f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.835
cc_5 VNB GATE 0.00262154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_GATE_c_169_n 0.0370731f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_7 VNB N_GATE_c_170_n 0.0227676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_235_74#_c_210_n 0.0118411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_235_74#_M1021_g 0.025926f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_10 VNB N_A_235_74#_c_212_n 0.0166873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_235_74#_c_213_n 0.00208209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_235_74#_M1015_g 0.0368511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_235_74#_c_215_n 0.0292038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_235_74#_c_216_n 0.00718515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_235_74#_c_217_n 0.00368649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_235_74#_c_218_n 0.00878693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_235_74#_c_219_n 9.77433e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_235_74#_c_220_n 0.0149319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_235_74#_c_221_n 0.00217878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_235_74#_c_222_n 0.0013407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_235_74#_c_223_n 0.0379701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_235_74#_c_224_n 0.00850203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_392#_c_361_n 0.0223813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_392#_M1000_g 0.0340105f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_25 VNB N_A_27_392#_c_363_n 0.025219f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_26 VNB N_A_27_392#_c_364_n 0.00531987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_392#_c_365_n 0.00984315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_392#_c_366_n 0.00700458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_392#_c_367_n 0.00174573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_347_98#_c_458_n 0.00308891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_347_98#_c_459_n 0.0253554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_347_98#_c_460_n 0.0031413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_347_98#_c_461_n 0.00262021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_347_98#_c_462_n 0.0330043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_347_98#_c_463_n 0.0180454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_832_55#_c_573_n 0.0165761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_832_55#_c_574_n 0.0356667f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_38 VNB N_A_832_55#_M1004_g 0.0229601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_832_55#_M1013_g 0.0226634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_832_55#_c_577_n 0.0231996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_832_55#_c_578_n 0.00819495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_832_55#_c_579_n 0.00254477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_832_55#_c_580_n 0.00550664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_832_55#_c_581_n 0.00318073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_832_55#_c_582_n 0.0567986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_646_74#_M1011_g 0.0266145f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_47 VNB N_A_646_74#_c_705_n 0.031895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_646_74#_c_706_n 0.0133901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_646_74#_c_707_n 8.48194e-19 $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_50 VNB N_A_646_74#_c_708_n 0.011705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_646_74#_c_709_n 0.00819016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_RESET_B_c_793_n 0.0183889f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_53 VNB N_RESET_B_c_794_n 0.033804f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.45
cc_54 VNB N_RESET_B_c_795_n 0.013192f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_55 VNB N_VPWR_c_828_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_Q_c_917_n 0.00248769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_Q_c_918_n 0.00893082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_Q_c_919_n 0.00236567f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_59 VNB Q 0.0266172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_961_n 0.0168478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_962_n 0.0203039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_963_n 0.00913215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_964_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_965_n 0.0289884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_966_n 0.0175013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_967_n 0.0350547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_968_n 0.039317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_969_n 0.0329481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_970_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_971_n 0.0274122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_972_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_973_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_974_n 0.414379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VPB N_D_c_139_n 0.0476472f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_75 VPB N_D_c_141_n 0.00541046f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_76 VPB N_GATE_c_167_n 0.00874321f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.835
cc_77 VPB N_GATE_c_172_n 0.0274537f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.835
cc_78 VPB N_A_235_74#_c_210_n 0.0326134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_235_74#_c_226_n 0.0148923f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_235_74#_c_212_n 0.0366005f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_235_74#_c_213_n 0.0115319f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_235_74#_c_215_n 0.0201498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_235_74#_c_230_n 0.00456571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_235_74#_c_231_n 0.0119485f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_235_74#_c_221_n 0.00119273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_235_74#_c_223_n 0.00741039f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_27_392#_c_361_n 0.0361325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_27_392#_c_366_n 0.00623345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_27_392#_c_370_n 0.00871078f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_27_392#_c_371_n 0.00142025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_27_392#_c_372_n 0.0431375f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_347_98#_c_464_n 0.0165629f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.615
cc_93 VPB N_A_347_98#_c_458_n 0.00227525f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_347_98#_c_460_n 0.00221225f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_347_98#_c_467_n 0.00654345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_347_98#_c_468_n 0.00214892f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_347_98#_c_469_n 0.00176728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_347_98#_c_470_n 0.00256782f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_347_98#_c_471_n 0.00574392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_347_98#_c_472_n 0.0516286f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_832_55#_c_574_n 0.0285625f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_102 VPB N_A_832_55#_c_584_n 0.057088f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_103 VPB N_A_832_55#_c_585_n 0.0162631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_832_55#_c_586_n 0.0165709f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_832_55#_c_587_n 0.00653784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_832_55#_c_588_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_832_55#_c_589_n 0.00807721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_832_55#_c_579_n 8.97934e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_832_55#_c_591_n 0.00757242f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_832_55#_c_581_n 2.97853e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_832_55#_c_582_n 0.0133109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_646_74#_c_710_n 0.017194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_646_74#_c_705_n 0.013969f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_646_74#_c_706_n 0.00652232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_646_74#_c_713_n 0.0307003f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_646_74#_c_709_n 0.00129873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_646_74#_c_715_n 8.46624e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_646_74#_c_716_n 0.00663645f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_646_74#_c_717_n 0.00339684f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_RESET_B_c_794_n 0.0226672f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.45
cc_121 VPB N_VPWR_c_829_n 0.0204215f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_830_n 0.0142301f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_831_n 0.00830446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_832_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_833_n 0.0442244f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_834_n 0.036437f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_835_n 0.00631927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_836_n 0.0467908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_837_n 0.0187266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_838_n 0.018682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_839_n 0.0264984f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_840_n 0.0210825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_841_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_828_n 0.0973179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_Q_c_921_n 0.00129357f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_136 VPB N_Q_c_922_n 0.00290132f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_137 VPB N_Q_c_923_n 0.00882548f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB Q 0.00708423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 N_D_c_139_n N_GATE_c_167_n 0.0064837f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_140 N_D_c_139_n N_GATE_c_172_n 0.0210224f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_141 N_D_M1006_g N_GATE_c_169_n 0.00782333f $X=0.52 $Y=0.835 $X2=0 $Y2=0
cc_142 N_D_M1006_g N_GATE_c_170_n 0.0163764f $X=0.52 $Y=0.835 $X2=0 $Y2=0
cc_143 N_D_M1006_g N_A_235_74#_c_220_n 4.146e-19 $X=0.52 $Y=0.835 $X2=0 $Y2=0
cc_144 N_D_c_139_n N_A_235_74#_c_231_n 2.43556e-19 $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_145 N_D_M1006_g N_A_27_392#_c_363_n 0.0116684f $X=0.52 $Y=0.835 $X2=0 $Y2=0
cc_146 N_D_M1006_g N_A_27_392#_c_364_n 0.0124006f $X=0.52 $Y=0.835 $X2=0 $Y2=0
cc_147 N_D_c_141_n N_A_27_392#_c_364_n 0.00317967f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_148 N_D_c_139_n N_A_27_392#_c_365_n 0.00532044f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_149 N_D_M1006_g N_A_27_392#_c_365_n 0.00417698f $X=0.52 $Y=0.835 $X2=0 $Y2=0
cc_150 N_D_c_141_n N_A_27_392#_c_365_n 0.0280475f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_151 N_D_c_139_n N_A_27_392#_c_366_n 0.00156941f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_152 N_D_M1006_g N_A_27_392#_c_366_n 0.00987116f $X=0.52 $Y=0.835 $X2=0 $Y2=0
cc_153 N_D_c_141_n N_A_27_392#_c_366_n 0.0250891f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_154 N_D_c_139_n N_A_27_392#_c_372_n 0.0382168f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_155 N_D_c_141_n N_A_27_392#_c_372_n 0.0328854f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_156 N_D_c_139_n N_VPWR_c_829_n 0.00357566f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_157 N_D_c_139_n N_VPWR_c_839_n 0.00365184f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_158 N_D_c_139_n N_VPWR_c_828_n 0.0049649f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_159 N_D_M1006_g N_VGND_c_961_n 0.00567863f $X=0.52 $Y=0.835 $X2=0 $Y2=0
cc_160 N_D_M1006_g N_VGND_c_971_n 0.0043356f $X=0.52 $Y=0.835 $X2=0 $Y2=0
cc_161 N_D_M1006_g N_VGND_c_974_n 0.00487769f $X=0.52 $Y=0.835 $X2=0 $Y2=0
cc_162 N_GATE_c_167_n N_A_235_74#_c_215_n 0.00632258f $X=1.125 $Y=1.795 $X2=0
+ $Y2=0
cc_163 N_GATE_c_169_n N_A_235_74#_c_215_n 0.00685518f $X=1.155 $Y=1.385 $X2=0
+ $Y2=0
cc_164 GATE N_A_235_74#_c_216_n 0.0178735f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_165 N_GATE_c_169_n N_A_235_74#_c_216_n 0.00467249f $X=1.155 $Y=1.385 $X2=0
+ $Y2=0
cc_166 N_GATE_c_170_n N_A_235_74#_c_216_n 0.00346505f $X=1.155 $Y=1.22 $X2=0
+ $Y2=0
cc_167 N_GATE_c_167_n N_A_235_74#_c_230_n 0.0029667f $X=1.125 $Y=1.795 $X2=0
+ $Y2=0
cc_168 N_GATE_c_172_n N_A_235_74#_c_230_n 0.00114122f $X=1.125 $Y=1.885 $X2=0
+ $Y2=0
cc_169 GATE N_A_235_74#_c_220_n 0.00888881f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_170 N_GATE_c_169_n N_A_235_74#_c_220_n 0.00212432f $X=1.155 $Y=1.385 $X2=0
+ $Y2=0
cc_171 N_GATE_c_170_n N_A_235_74#_c_220_n 0.00859891f $X=1.155 $Y=1.22 $X2=0
+ $Y2=0
cc_172 N_GATE_c_172_n N_A_235_74#_c_231_n 0.00586241f $X=1.125 $Y=1.885 $X2=0
+ $Y2=0
cc_173 GATE N_A_235_74#_c_231_n 0.00420322f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_174 N_GATE_c_169_n N_A_235_74#_c_231_n 0.00159251f $X=1.155 $Y=1.385 $X2=0
+ $Y2=0
cc_175 N_GATE_c_167_n N_A_235_74#_c_221_n 0.0021511f $X=1.125 $Y=1.795 $X2=0
+ $Y2=0
cc_176 GATE N_A_235_74#_c_221_n 0.0103132f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_177 N_GATE_c_169_n N_A_235_74#_c_221_n 8.58045e-19 $X=1.155 $Y=1.385 $X2=0
+ $Y2=0
cc_178 N_GATE_c_170_n N_A_27_392#_c_363_n 8.51597e-19 $X=1.155 $Y=1.22 $X2=0
+ $Y2=0
cc_179 GATE N_A_27_392#_c_364_n 0.00829681f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_180 N_GATE_c_169_n N_A_27_392#_c_364_n 5.43244e-19 $X=1.155 $Y=1.385 $X2=0
+ $Y2=0
cc_181 N_GATE_c_170_n N_A_27_392#_c_364_n 0.00128853f $X=1.155 $Y=1.22 $X2=0
+ $Y2=0
cc_182 N_GATE_c_167_n N_A_27_392#_c_366_n 0.00384357f $X=1.125 $Y=1.795 $X2=0
+ $Y2=0
cc_183 N_GATE_c_172_n N_A_27_392#_c_366_n 7.09582e-19 $X=1.125 $Y=1.885 $X2=0
+ $Y2=0
cc_184 GATE N_A_27_392#_c_366_n 0.0198903f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_185 N_GATE_c_169_n N_A_27_392#_c_366_n 0.00219339f $X=1.155 $Y=1.385 $X2=0
+ $Y2=0
cc_186 N_GATE_c_172_n N_A_27_392#_c_370_n 0.0187913f $X=1.125 $Y=1.885 $X2=0
+ $Y2=0
cc_187 N_GATE_c_172_n N_A_27_392#_c_372_n 0.0089078f $X=1.125 $Y=1.885 $X2=0
+ $Y2=0
cc_188 N_GATE_c_172_n N_A_347_98#_c_470_n 4.84431e-19 $X=1.125 $Y=1.885 $X2=0
+ $Y2=0
cc_189 N_GATE_c_172_n N_VPWR_c_829_n 0.00432851f $X=1.125 $Y=1.885 $X2=0 $Y2=0
cc_190 N_GATE_c_172_n N_VPWR_c_834_n 0.00366846f $X=1.125 $Y=1.885 $X2=0 $Y2=0
cc_191 N_GATE_c_172_n N_VPWR_c_828_n 0.0049649f $X=1.125 $Y=1.885 $X2=0 $Y2=0
cc_192 N_GATE_c_170_n N_VGND_c_961_n 0.00941074f $X=1.155 $Y=1.22 $X2=0 $Y2=0
cc_193 N_GATE_c_170_n N_VGND_c_967_n 0.00434272f $X=1.155 $Y=1.22 $X2=0 $Y2=0
cc_194 N_GATE_c_170_n N_VGND_c_974_n 0.00830058f $X=1.155 $Y=1.22 $X2=0 $Y2=0
cc_195 N_A_235_74#_c_210_n N_A_27_392#_c_361_n 0.0405505f $X=2.135 $Y=1.885
+ $X2=0 $Y2=0
cc_196 N_A_235_74#_c_226_n N_A_27_392#_c_361_n 0.0466055f $X=3.17 $Y=1.885 $X2=0
+ $Y2=0
cc_197 N_A_235_74#_c_213_n N_A_27_392#_c_361_n 0.0117039f $X=3.26 $Y=1.735 $X2=0
+ $Y2=0
cc_198 N_A_235_74#_M1021_g N_A_27_392#_M1000_g 0.029484f $X=2.175 $Y=0.86 $X2=0
+ $Y2=0
cc_199 N_A_235_74#_c_217_n N_A_27_392#_M1000_g 0.0113271f $X=2.805 $Y=0.665
+ $X2=0 $Y2=0
cc_200 N_A_235_74#_c_257_p N_A_27_392#_M1000_g 0.00400332f $X=2.89 $Y=0.58 $X2=0
+ $Y2=0
cc_201 N_A_235_74#_c_219_n N_A_27_392#_M1000_g 0.00401328f $X=2.975 $Y=0.34
+ $X2=0 $Y2=0
cc_202 N_A_235_74#_c_216_n N_A_27_392#_c_364_n 0.00243787f $X=1.54 $Y=1.42 $X2=0
+ $Y2=0
cc_203 N_A_235_74#_c_230_n N_A_27_392#_c_366_n 0.00589115f $X=1.54 $Y=1.94 $X2=0
+ $Y2=0
cc_204 N_A_235_74#_c_231_n N_A_27_392#_c_366_n 3.9843e-19 $X=1.54 $Y=2.105 $X2=0
+ $Y2=0
cc_205 N_A_235_74#_c_221_n N_A_27_392#_c_366_n 0.00665224f $X=1.725 $Y=1.585
+ $X2=0 $Y2=0
cc_206 N_A_235_74#_M1009_d N_A_27_392#_c_370_n 0.00814605f $X=1.2 $Y=1.96 $X2=0
+ $Y2=0
cc_207 N_A_235_74#_c_210_n N_A_27_392#_c_370_n 0.0146141f $X=2.135 $Y=1.885
+ $X2=0 $Y2=0
cc_208 N_A_235_74#_c_215_n N_A_27_392#_c_370_n 0.00456949f $X=2.045 $Y=1.585
+ $X2=0 $Y2=0
cc_209 N_A_235_74#_c_231_n N_A_27_392#_c_370_n 0.0295292f $X=1.54 $Y=2.105 $X2=0
+ $Y2=0
cc_210 N_A_235_74#_c_210_n N_A_27_392#_c_371_n 0.00508288f $X=2.135 $Y=1.885
+ $X2=0 $Y2=0
cc_211 N_A_235_74#_c_226_n N_A_27_392#_c_371_n 2.99642e-19 $X=3.17 $Y=1.885
+ $X2=0 $Y2=0
cc_212 N_A_235_74#_c_231_n N_A_27_392#_c_372_n 0.0162024f $X=1.54 $Y=2.105 $X2=0
+ $Y2=0
cc_213 N_A_235_74#_c_210_n N_A_27_392#_c_367_n 8.2736e-19 $X=2.135 $Y=1.885
+ $X2=0 $Y2=0
cc_214 N_A_235_74#_c_217_n N_A_347_98#_M1021_s 0.0102425f $X=2.805 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_215 N_A_235_74#_c_226_n N_A_347_98#_c_464_n 0.0128379f $X=3.17 $Y=1.885 $X2=0
+ $Y2=0
cc_216 N_A_235_74#_c_210_n N_A_347_98#_c_458_n 0.0190775f $X=2.135 $Y=1.885
+ $X2=0 $Y2=0
cc_217 N_A_235_74#_M1021_g N_A_347_98#_c_458_n 0.00750041f $X=2.175 $Y=0.86
+ $X2=0 $Y2=0
cc_218 N_A_235_74#_c_216_n N_A_347_98#_c_458_n 0.0066868f $X=1.54 $Y=1.42 $X2=0
+ $Y2=0
cc_219 N_A_235_74#_c_230_n N_A_347_98#_c_458_n 0.00673003f $X=1.54 $Y=1.94 $X2=0
+ $Y2=0
cc_220 N_A_235_74#_c_221_n N_A_347_98#_c_458_n 0.0240774f $X=1.725 $Y=1.585
+ $X2=0 $Y2=0
cc_221 N_A_235_74#_M1021_g N_A_347_98#_c_459_n 0.00417341f $X=2.175 $Y=0.86
+ $X2=0 $Y2=0
cc_222 N_A_235_74#_c_213_n N_A_347_98#_c_459_n 6.53802e-19 $X=3.26 $Y=1.735
+ $X2=0 $Y2=0
cc_223 N_A_235_74#_c_217_n N_A_347_98#_c_459_n 0.0282239f $X=2.805 $Y=0.665
+ $X2=0 $Y2=0
cc_224 N_A_235_74#_c_218_n N_A_347_98#_c_459_n 0.00532848f $X=3.92 $Y=0.34 $X2=0
+ $Y2=0
cc_225 N_A_235_74#_c_226_n N_A_347_98#_c_460_n 0.00154626f $X=3.17 $Y=1.885
+ $X2=0 $Y2=0
cc_226 N_A_235_74#_c_213_n N_A_347_98#_c_460_n 0.00796956f $X=3.26 $Y=1.735
+ $X2=0 $Y2=0
cc_227 N_A_235_74#_c_226_n N_A_347_98#_c_467_n 0.0132479f $X=3.17 $Y=1.885 $X2=0
+ $Y2=0
cc_228 N_A_235_74#_c_226_n N_A_347_98#_c_469_n 4.82699e-19 $X=3.17 $Y=1.885
+ $X2=0 $Y2=0
cc_229 N_A_235_74#_M1021_g N_A_347_98#_c_461_n 0.0155579f $X=2.175 $Y=0.86 $X2=0
+ $Y2=0
cc_230 N_A_235_74#_c_215_n N_A_347_98#_c_461_n 0.00908545f $X=2.045 $Y=1.585
+ $X2=0 $Y2=0
cc_231 N_A_235_74#_c_217_n N_A_347_98#_c_461_n 0.0282363f $X=2.805 $Y=0.665
+ $X2=0 $Y2=0
cc_232 N_A_235_74#_c_220_n N_A_347_98#_c_461_n 0.0272269f $X=1.315 $Y=0.515
+ $X2=0 $Y2=0
cc_233 N_A_235_74#_c_221_n N_A_347_98#_c_461_n 0.00751825f $X=1.725 $Y=1.585
+ $X2=0 $Y2=0
cc_234 N_A_235_74#_c_210_n N_A_347_98#_c_470_n 0.0107038f $X=2.135 $Y=1.885
+ $X2=0 $Y2=0
cc_235 N_A_235_74#_c_215_n N_A_347_98#_c_470_n 0.00757595f $X=2.045 $Y=1.585
+ $X2=0 $Y2=0
cc_236 N_A_235_74#_c_231_n N_A_347_98#_c_470_n 0.0249765f $X=1.54 $Y=2.105 $X2=0
+ $Y2=0
cc_237 N_A_235_74#_c_221_n N_A_347_98#_c_470_n 0.00473243f $X=1.725 $Y=1.585
+ $X2=0 $Y2=0
cc_238 N_A_235_74#_c_226_n N_A_347_98#_c_471_n 0.0101667f $X=3.17 $Y=1.885 $X2=0
+ $Y2=0
cc_239 N_A_235_74#_c_213_n N_A_347_98#_c_462_n 0.0195624f $X=3.26 $Y=1.735 $X2=0
+ $Y2=0
cc_240 N_A_235_74#_M1015_g N_A_347_98#_c_462_n 0.00321247f $X=3.845 $Y=0.615
+ $X2=0 $Y2=0
cc_241 N_A_235_74#_c_223_n N_A_347_98#_c_462_n 0.00481586f $X=3.925 $Y=1.425
+ $X2=0 $Y2=0
cc_242 N_A_235_74#_M1015_g N_A_347_98#_c_463_n 0.0138977f $X=3.845 $Y=0.615
+ $X2=0 $Y2=0
cc_243 N_A_235_74#_c_217_n N_A_347_98#_c_463_n 0.00168224f $X=2.805 $Y=0.665
+ $X2=0 $Y2=0
cc_244 N_A_235_74#_c_257_p N_A_347_98#_c_463_n 0.00336012f $X=2.89 $Y=0.58 $X2=0
+ $Y2=0
cc_245 N_A_235_74#_c_218_n N_A_347_98#_c_463_n 0.0119273f $X=3.92 $Y=0.34 $X2=0
+ $Y2=0
cc_246 N_A_235_74#_c_226_n N_A_347_98#_c_472_n 0.00937594f $X=3.17 $Y=1.885
+ $X2=0 $Y2=0
cc_247 N_A_235_74#_c_212_n N_A_347_98#_c_472_n 0.015892f $X=3.76 $Y=1.735 $X2=0
+ $Y2=0
cc_248 N_A_235_74#_c_223_n N_A_347_98#_c_472_n 0.00309466f $X=3.925 $Y=1.425
+ $X2=0 $Y2=0
cc_249 N_A_235_74#_M1015_g N_A_832_55#_c_573_n 0.0347794f $X=3.845 $Y=0.615
+ $X2=0 $Y2=0
cc_250 N_A_235_74#_c_218_n N_A_832_55#_c_573_n 0.00117076f $X=3.92 $Y=0.34 $X2=0
+ $Y2=0
cc_251 N_A_235_74#_c_224_n N_A_832_55#_c_573_n 0.00754794f $X=3.957 $Y=1.26
+ $X2=0 $Y2=0
cc_252 N_A_235_74#_M1015_g N_A_832_55#_c_574_n 0.00477445f $X=3.845 $Y=0.615
+ $X2=0 $Y2=0
cc_253 N_A_235_74#_c_222_n N_A_832_55#_c_574_n 0.00153666f $X=3.925 $Y=1.425
+ $X2=0 $Y2=0
cc_254 N_A_235_74#_c_223_n N_A_832_55#_c_574_n 0.0281443f $X=3.925 $Y=1.425
+ $X2=0 $Y2=0
cc_255 N_A_235_74#_c_224_n N_A_832_55#_c_574_n 0.00431668f $X=3.957 $Y=1.26
+ $X2=0 $Y2=0
cc_256 N_A_235_74#_c_218_n N_A_646_74#_M1001_d 0.00478265f $X=3.92 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_257 N_A_235_74#_M1015_g N_A_646_74#_c_707_n 0.00190538f $X=3.845 $Y=0.615
+ $X2=0 $Y2=0
cc_258 N_A_235_74#_c_217_n N_A_646_74#_c_707_n 0.0104267f $X=2.805 $Y=0.665
+ $X2=0 $Y2=0
cc_259 N_A_235_74#_c_218_n N_A_646_74#_c_707_n 0.0325532f $X=3.92 $Y=0.34 $X2=0
+ $Y2=0
cc_260 N_A_235_74#_c_224_n N_A_646_74#_c_707_n 0.00137358f $X=3.957 $Y=1.26
+ $X2=0 $Y2=0
cc_261 N_A_235_74#_c_212_n N_A_646_74#_c_708_n 0.00914778f $X=3.76 $Y=1.735
+ $X2=0 $Y2=0
cc_262 N_A_235_74#_M1015_g N_A_646_74#_c_708_n 0.00399052f $X=3.845 $Y=0.615
+ $X2=0 $Y2=0
cc_263 N_A_235_74#_c_222_n N_A_646_74#_c_708_n 0.0243903f $X=3.925 $Y=1.425
+ $X2=0 $Y2=0
cc_264 N_A_235_74#_c_223_n N_A_646_74#_c_708_n 0.00756358f $X=3.925 $Y=1.425
+ $X2=0 $Y2=0
cc_265 N_A_235_74#_c_224_n N_A_646_74#_c_708_n 0.0226172f $X=3.957 $Y=1.26 $X2=0
+ $Y2=0
cc_266 N_A_235_74#_c_212_n N_A_646_74#_c_713_n 0.00494965f $X=3.76 $Y=1.735
+ $X2=0 $Y2=0
cc_267 N_A_235_74#_c_222_n N_A_646_74#_c_713_n 0.0202911f $X=3.925 $Y=1.425
+ $X2=0 $Y2=0
cc_268 N_A_235_74#_c_223_n N_A_646_74#_c_713_n 0.0070896f $X=3.925 $Y=1.425
+ $X2=0 $Y2=0
cc_269 N_A_235_74#_c_222_n N_A_646_74#_c_709_n 0.00641528f $X=3.925 $Y=1.425
+ $X2=0 $Y2=0
cc_270 N_A_235_74#_c_226_n N_A_646_74#_c_715_n 0.00390285f $X=3.17 $Y=1.885
+ $X2=0 $Y2=0
cc_271 N_A_235_74#_c_212_n N_A_646_74#_c_715_n 0.00254916f $X=3.76 $Y=1.735
+ $X2=0 $Y2=0
cc_272 N_A_235_74#_c_226_n N_A_646_74#_c_716_n 0.00521023f $X=3.17 $Y=1.885
+ $X2=0 $Y2=0
cc_273 N_A_235_74#_c_226_n N_A_646_74#_c_717_n 9.08877e-19 $X=3.17 $Y=1.885
+ $X2=0 $Y2=0
cc_274 N_A_235_74#_c_212_n N_A_646_74#_c_717_n 0.0114093f $X=3.76 $Y=1.735 $X2=0
+ $Y2=0
cc_275 N_A_235_74#_c_213_n N_A_646_74#_c_717_n 0.00162887f $X=3.26 $Y=1.735
+ $X2=0 $Y2=0
cc_276 N_A_235_74#_c_210_n N_VPWR_c_830_n 0.00432032f $X=2.135 $Y=1.885 $X2=0
+ $Y2=0
cc_277 N_A_235_74#_c_210_n N_VPWR_c_834_n 0.00366846f $X=2.135 $Y=1.885 $X2=0
+ $Y2=0
cc_278 N_A_235_74#_c_226_n N_VPWR_c_836_n 0.00278271f $X=3.17 $Y=1.885 $X2=0
+ $Y2=0
cc_279 N_A_235_74#_c_210_n N_VPWR_c_828_n 0.0049649f $X=2.135 $Y=1.885 $X2=0
+ $Y2=0
cc_280 N_A_235_74#_c_226_n N_VPWR_c_828_n 0.00354422f $X=3.17 $Y=1.885 $X2=0
+ $Y2=0
cc_281 N_A_235_74#_c_217_n N_VGND_M1021_d 0.0086219f $X=2.805 $Y=0.665 $X2=0
+ $Y2=0
cc_282 N_A_235_74#_c_220_n N_VGND_c_961_n 0.024197f $X=1.315 $Y=0.515 $X2=0
+ $Y2=0
cc_283 N_A_235_74#_c_218_n N_VGND_c_962_n 0.0129787f $X=3.92 $Y=0.34 $X2=0 $Y2=0
cc_284 N_A_235_74#_c_224_n N_VGND_c_962_n 0.0278898f $X=3.957 $Y=1.26 $X2=0
+ $Y2=0
cc_285 N_A_235_74#_M1021_g N_VGND_c_966_n 0.0014541f $X=2.175 $Y=0.86 $X2=0
+ $Y2=0
cc_286 N_A_235_74#_c_217_n N_VGND_c_966_n 0.0244722f $X=2.805 $Y=0.665 $X2=0
+ $Y2=0
cc_287 N_A_235_74#_c_219_n N_VGND_c_966_n 0.0112922f $X=2.975 $Y=0.34 $X2=0
+ $Y2=0
cc_288 N_A_235_74#_M1021_g N_VGND_c_967_n 0.00374721f $X=2.175 $Y=0.86 $X2=0
+ $Y2=0
cc_289 N_A_235_74#_c_217_n N_VGND_c_967_n 0.0124277f $X=2.805 $Y=0.665 $X2=0
+ $Y2=0
cc_290 N_A_235_74#_c_220_n N_VGND_c_967_n 0.0210047f $X=1.315 $Y=0.515 $X2=0
+ $Y2=0
cc_291 N_A_235_74#_M1015_g N_VGND_c_968_n 9.35083e-19 $X=3.845 $Y=0.615 $X2=0
+ $Y2=0
cc_292 N_A_235_74#_c_217_n N_VGND_c_968_n 0.00275846f $X=2.805 $Y=0.665 $X2=0
+ $Y2=0
cc_293 N_A_235_74#_c_218_n N_VGND_c_968_n 0.0725671f $X=3.92 $Y=0.34 $X2=0 $Y2=0
cc_294 N_A_235_74#_c_219_n N_VGND_c_968_n 0.0117819f $X=2.975 $Y=0.34 $X2=0
+ $Y2=0
cc_295 N_A_235_74#_M1021_g N_VGND_c_974_n 0.00508379f $X=2.175 $Y=0.86 $X2=0
+ $Y2=0
cc_296 N_A_235_74#_c_217_n N_VGND_c_974_n 0.0263281f $X=2.805 $Y=0.665 $X2=0
+ $Y2=0
cc_297 N_A_235_74#_c_218_n N_VGND_c_974_n 0.0414485f $X=3.92 $Y=0.34 $X2=0 $Y2=0
cc_298 N_A_235_74#_c_219_n N_VGND_c_974_n 0.0063954f $X=2.975 $Y=0.34 $X2=0
+ $Y2=0
cc_299 N_A_235_74#_c_220_n N_VGND_c_974_n 0.0173423f $X=1.315 $Y=0.515 $X2=0
+ $Y2=0
cc_300 N_A_235_74#_c_217_n A_568_74# 0.00286327f $X=2.805 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_301 N_A_235_74#_c_257_p A_568_74# 0.00171077f $X=2.89 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_302 N_A_235_74#_c_218_n A_568_74# 9.80156e-19 $X=3.92 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_303 N_A_235_74#_c_224_n A_784_81# 0.00479806f $X=3.957 $Y=1.26 $X2=-0.19
+ $Y2=-0.245
cc_304 N_A_27_392#_c_370_n N_A_347_98#_M1017_s 0.00845913f $X=2.51 $Y=2.525
+ $X2=0 $Y2=0
cc_305 N_A_27_392#_c_361_n N_A_347_98#_c_458_n 0.00216731f $X=2.75 $Y=1.885
+ $X2=0 $Y2=0
cc_306 N_A_27_392#_M1000_g N_A_347_98#_c_458_n 0.00102671f $X=2.765 $Y=0.69
+ $X2=0 $Y2=0
cc_307 N_A_27_392#_c_367_n N_A_347_98#_c_458_n 0.0256095f $X=2.675 $Y=1.605
+ $X2=0 $Y2=0
cc_308 N_A_27_392#_c_361_n N_A_347_98#_c_459_n 0.00123009f $X=2.75 $Y=1.885
+ $X2=0 $Y2=0
cc_309 N_A_27_392#_M1000_g N_A_347_98#_c_459_n 0.0130896f $X=2.765 $Y=0.69 $X2=0
+ $Y2=0
cc_310 N_A_27_392#_c_367_n N_A_347_98#_c_459_n 0.0440002f $X=2.675 $Y=1.605
+ $X2=0 $Y2=0
cc_311 N_A_27_392#_c_361_n N_A_347_98#_c_516_n 0.00865258f $X=2.75 $Y=1.885
+ $X2=0 $Y2=0
cc_312 N_A_27_392#_c_370_n N_A_347_98#_c_516_n 0.0113396f $X=2.51 $Y=2.525 $X2=0
+ $Y2=0
cc_313 N_A_27_392#_c_371_n N_A_347_98#_c_516_n 0.0196638f $X=2.595 $Y=2.44 $X2=0
+ $Y2=0
cc_314 N_A_27_392#_c_361_n N_A_347_98#_c_460_n 0.00637387f $X=2.75 $Y=1.885
+ $X2=0 $Y2=0
cc_315 N_A_27_392#_c_371_n N_A_347_98#_c_460_n 0.00677755f $X=2.595 $Y=2.44
+ $X2=0 $Y2=0
cc_316 N_A_27_392#_c_361_n N_A_347_98#_c_468_n 0.00168766f $X=2.75 $Y=1.885
+ $X2=0 $Y2=0
cc_317 N_A_27_392#_M1000_g N_A_347_98#_c_461_n 8.55919e-19 $X=2.765 $Y=0.69
+ $X2=0 $Y2=0
cc_318 N_A_27_392#_c_361_n N_A_347_98#_c_470_n 2.5705e-19 $X=2.75 $Y=1.885 $X2=0
+ $Y2=0
cc_319 N_A_27_392#_c_370_n N_A_347_98#_c_470_n 0.0242436f $X=2.51 $Y=2.525 $X2=0
+ $Y2=0
cc_320 N_A_27_392#_c_371_n N_A_347_98#_c_470_n 0.00884827f $X=2.595 $Y=2.44
+ $X2=0 $Y2=0
cc_321 N_A_27_392#_c_361_n N_A_347_98#_c_471_n 0.00131666f $X=2.75 $Y=1.885
+ $X2=0 $Y2=0
cc_322 N_A_27_392#_c_371_n N_A_347_98#_c_471_n 0.0106432f $X=2.595 $Y=2.44 $X2=0
+ $Y2=0
cc_323 N_A_27_392#_M1000_g N_A_347_98#_c_462_n 0.0211809f $X=2.765 $Y=0.69 $X2=0
+ $Y2=0
cc_324 N_A_27_392#_M1000_g N_A_347_98#_c_463_n 0.0464649f $X=2.765 $Y=0.69 $X2=0
+ $Y2=0
cc_325 N_A_27_392#_M1000_g N_A_646_74#_c_707_n 5.95138e-19 $X=2.765 $Y=0.69
+ $X2=0 $Y2=0
cc_326 N_A_27_392#_c_370_n N_VPWR_M1012_d 0.0068796f $X=2.51 $Y=2.525 $X2=-0.19
+ $Y2=-0.245
cc_327 N_A_27_392#_c_372_n N_VPWR_M1012_d 0.0118348f $X=0.28 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_328 N_A_27_392#_c_370_n N_VPWR_M1017_d 0.0140367f $X=2.51 $Y=2.525 $X2=0
+ $Y2=0
cc_329 N_A_27_392#_c_371_n N_VPWR_M1017_d 0.00551492f $X=2.595 $Y=2.44 $X2=0
+ $Y2=0
cc_330 N_A_27_392#_c_370_n N_VPWR_c_829_n 0.00965353f $X=2.51 $Y=2.525 $X2=0
+ $Y2=0
cc_331 N_A_27_392#_c_372_n N_VPWR_c_829_n 0.0203314f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_332 N_A_27_392#_c_361_n N_VPWR_c_830_n 0.00574461f $X=2.75 $Y=1.885 $X2=0
+ $Y2=0
cc_333 N_A_27_392#_c_370_n N_VPWR_c_830_n 0.0263592f $X=2.51 $Y=2.525 $X2=0
+ $Y2=0
cc_334 N_A_27_392#_c_370_n N_VPWR_c_834_n 0.0172927f $X=2.51 $Y=2.525 $X2=0
+ $Y2=0
cc_335 N_A_27_392#_c_361_n N_VPWR_c_836_n 0.00457248f $X=2.75 $Y=1.885 $X2=0
+ $Y2=0
cc_336 N_A_27_392#_c_370_n N_VPWR_c_836_n 6.37789e-19 $X=2.51 $Y=2.525 $X2=0
+ $Y2=0
cc_337 N_A_27_392#_c_372_n N_VPWR_c_839_n 0.0115119f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_338 N_A_27_392#_c_361_n N_VPWR_c_828_n 0.00897726f $X=2.75 $Y=1.885 $X2=0
+ $Y2=0
cc_339 N_A_27_392#_c_370_n N_VPWR_c_828_n 0.038311f $X=2.51 $Y=2.525 $X2=0 $Y2=0
cc_340 N_A_27_392#_c_372_n N_VPWR_c_828_n 0.0175462f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_341 N_A_27_392#_c_364_n N_VGND_M1006_d 0.00188126f $X=0.685 $Y=1.195
+ $X2=-0.19 $Y2=-0.245
cc_342 N_A_27_392#_c_363_n N_VGND_c_961_n 0.0150958f $X=0.305 $Y=0.835 $X2=0
+ $Y2=0
cc_343 N_A_27_392#_c_364_n N_VGND_c_961_n 0.0180563f $X=0.685 $Y=1.195 $X2=0
+ $Y2=0
cc_344 N_A_27_392#_M1000_g N_VGND_c_966_n 0.00328112f $X=2.765 $Y=0.69 $X2=0
+ $Y2=0
cc_345 N_A_27_392#_M1000_g N_VGND_c_968_n 0.00310328f $X=2.765 $Y=0.69 $X2=0
+ $Y2=0
cc_346 N_A_27_392#_c_363_n N_VGND_c_971_n 0.0081488f $X=0.305 $Y=0.835 $X2=0
+ $Y2=0
cc_347 N_A_27_392#_M1000_g N_VGND_c_974_n 0.00393394f $X=2.765 $Y=0.69 $X2=0
+ $Y2=0
cc_348 N_A_27_392#_c_363_n N_VGND_c_974_n 0.0106395f $X=0.305 $Y=0.835 $X2=0
+ $Y2=0
cc_349 N_A_347_98#_c_464_n N_A_832_55#_c_584_n 0.00984643f $X=3.705 $Y=2.465
+ $X2=0 $Y2=0
cc_350 N_A_347_98#_c_467_n N_A_832_55#_c_584_n 0.00177437f $X=3.73 $Y=2.99 $X2=0
+ $Y2=0
cc_351 N_A_347_98#_c_469_n N_A_832_55#_c_584_n 0.00913042f $X=3.895 $Y=2.215
+ $X2=0 $Y2=0
cc_352 N_A_347_98#_c_472_n N_A_832_55#_c_584_n 0.0201499f $X=3.705 $Y=2.257
+ $X2=0 $Y2=0
cc_353 N_A_347_98#_c_469_n N_A_832_55#_c_587_n 0.016823f $X=3.895 $Y=2.215 $X2=0
+ $Y2=0
cc_354 N_A_347_98#_c_472_n N_A_832_55#_c_587_n 0.00108126f $X=3.705 $Y=2.257
+ $X2=0 $Y2=0
cc_355 N_A_347_98#_c_467_n N_A_646_74#_M1008_d 0.00334086f $X=3.73 $Y=2.99 $X2=0
+ $Y2=0
cc_356 N_A_347_98#_c_459_n N_A_646_74#_c_707_n 0.00514946f $X=3.05 $Y=1.165
+ $X2=0 $Y2=0
cc_357 N_A_347_98#_c_462_n N_A_646_74#_c_707_n 0.00268414f $X=3.215 $Y=1.285
+ $X2=0 $Y2=0
cc_358 N_A_347_98#_c_463_n N_A_646_74#_c_707_n 0.00859693f $X=3.215 $Y=1.12
+ $X2=0 $Y2=0
cc_359 N_A_347_98#_c_459_n N_A_646_74#_c_708_n 0.027507f $X=3.05 $Y=1.165 $X2=0
+ $Y2=0
cc_360 N_A_347_98#_c_460_n N_A_646_74#_c_708_n 0.0163151f $X=3.135 $Y=1.94 $X2=0
+ $Y2=0
cc_361 N_A_347_98#_c_462_n N_A_646_74#_c_708_n 0.00280153f $X=3.215 $Y=1.285
+ $X2=0 $Y2=0
cc_362 N_A_347_98#_c_463_n N_A_646_74#_c_708_n 0.00500291f $X=3.215 $Y=1.12
+ $X2=0 $Y2=0
cc_363 N_A_347_98#_c_469_n N_A_646_74#_c_713_n 0.0262108f $X=3.895 $Y=2.215
+ $X2=0 $Y2=0
cc_364 N_A_347_98#_c_472_n N_A_646_74#_c_713_n 0.00427327f $X=3.705 $Y=2.257
+ $X2=0 $Y2=0
cc_365 N_A_347_98#_c_464_n N_A_646_74#_c_715_n 0.00229161f $X=3.705 $Y=2.465
+ $X2=0 $Y2=0
cc_366 N_A_347_98#_c_467_n N_A_646_74#_c_715_n 0.0201163f $X=3.73 $Y=2.99 $X2=0
+ $Y2=0
cc_367 N_A_347_98#_c_460_n N_A_646_74#_c_716_n 6.77588e-19 $X=3.135 $Y=1.94
+ $X2=0 $Y2=0
cc_368 N_A_347_98#_c_469_n N_A_646_74#_c_716_n 0.0486637f $X=3.895 $Y=2.215
+ $X2=0 $Y2=0
cc_369 N_A_347_98#_c_471_n N_A_646_74#_c_716_n 0.0124923f $X=3.135 $Y=2.025
+ $X2=0 $Y2=0
cc_370 N_A_347_98#_c_472_n N_A_646_74#_c_716_n 0.00476054f $X=3.705 $Y=2.257
+ $X2=0 $Y2=0
cc_371 N_A_347_98#_c_460_n N_A_646_74#_c_717_n 0.0134563f $X=3.135 $Y=1.94 $X2=0
+ $Y2=0
cc_372 N_A_347_98#_c_472_n N_A_646_74#_c_717_n 0.00117204f $X=3.705 $Y=2.257
+ $X2=0 $Y2=0
cc_373 N_A_347_98#_c_516_n N_VPWR_c_830_n 0.00658881f $X=2.975 $Y=2.905 $X2=0
+ $Y2=0
cc_374 N_A_347_98#_c_468_n N_VPWR_c_830_n 0.0104027f $X=3.06 $Y=2.99 $X2=0 $Y2=0
cc_375 N_A_347_98#_c_464_n N_VPWR_c_836_n 0.00278223f $X=3.705 $Y=2.465 $X2=0
+ $Y2=0
cc_376 N_A_347_98#_c_467_n N_VPWR_c_836_n 0.0658254f $X=3.73 $Y=2.99 $X2=0 $Y2=0
cc_377 N_A_347_98#_c_468_n N_VPWR_c_836_n 0.0121867f $X=3.06 $Y=2.99 $X2=0 $Y2=0
cc_378 N_A_347_98#_c_464_n N_VPWR_c_840_n 3.91083e-19 $X=3.705 $Y=2.465 $X2=0
+ $Y2=0
cc_379 N_A_347_98#_c_467_n N_VPWR_c_840_n 0.00796543f $X=3.73 $Y=2.99 $X2=0
+ $Y2=0
cc_380 N_A_347_98#_c_469_n N_VPWR_c_840_n 0.0109461f $X=3.895 $Y=2.215 $X2=0
+ $Y2=0
cc_381 N_A_347_98#_c_464_n N_VPWR_c_828_n 0.00356419f $X=3.705 $Y=2.465 $X2=0
+ $Y2=0
cc_382 N_A_347_98#_c_467_n N_VPWR_c_828_n 0.0366416f $X=3.73 $Y=2.99 $X2=0 $Y2=0
cc_383 N_A_347_98#_c_468_n N_VPWR_c_828_n 0.00660921f $X=3.06 $Y=2.99 $X2=0
+ $Y2=0
cc_384 N_A_347_98#_c_516_n A_565_392# 0.0119697f $X=2.975 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_385 N_A_347_98#_c_468_n A_565_392# 6.47146e-19 $X=3.06 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_386 N_A_347_98#_c_471_n A_565_392# 0.00189564f $X=3.135 $Y=2.025 $X2=-0.19
+ $Y2=-0.245
cc_387 N_A_347_98#_c_467_n A_756_508# 0.00100794f $X=3.73 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_388 N_A_347_98#_c_469_n A_756_508# 0.00646594f $X=3.895 $Y=2.215 $X2=-0.19
+ $Y2=-0.245
cc_389 N_A_347_98#_c_459_n N_VGND_M1021_d 0.00337951f $X=3.05 $Y=1.165 $X2=0
+ $Y2=0
cc_390 N_A_347_98#_c_463_n N_VGND_c_968_n 0.00278271f $X=3.215 $Y=1.12 $X2=0
+ $Y2=0
cc_391 N_A_347_98#_c_463_n N_VGND_c_974_n 0.00358137f $X=3.215 $Y=1.12 $X2=0
+ $Y2=0
cc_392 N_A_832_55#_c_574_n N_A_646_74#_c_710_n 0.00317977f $X=4.375 $Y=2.05
+ $X2=0 $Y2=0
cc_393 N_A_832_55#_c_584_n N_A_646_74#_c_710_n 0.0174329f $X=4.39 $Y=2.465 $X2=0
+ $Y2=0
cc_394 N_A_832_55#_c_588_n N_A_646_74#_c_710_n 0.0154137f $X=5.42 $Y=2.815 $X2=0
+ $Y2=0
cc_395 N_A_832_55#_c_591_n N_A_646_74#_c_710_n 0.0222468f $X=5.34 $Y=1.805 $X2=0
+ $Y2=0
cc_396 N_A_832_55#_c_577_n N_A_646_74#_M1011_g 0.00374527f $X=4.375 $Y=0.975
+ $X2=0 $Y2=0
cc_397 N_A_832_55#_c_578_n N_A_646_74#_M1011_g 0.0155425f $X=5.01 $Y=0.515 $X2=0
+ $Y2=0
cc_398 N_A_832_55#_c_580_n N_A_646_74#_M1011_g 0.00534707f $X=5.055 $Y=1.13
+ $X2=0 $Y2=0
cc_399 N_A_832_55#_c_581_n N_A_646_74#_M1011_g 0.00636408f $X=5.34 $Y=1.72 $X2=0
+ $Y2=0
cc_400 N_A_832_55#_c_574_n N_A_646_74#_c_705_n 0.0216901f $X=4.375 $Y=2.05 $X2=0
+ $Y2=0
cc_401 N_A_832_55#_c_587_n N_A_646_74#_c_705_n 0.00581447f $X=5.095 $Y=2.24
+ $X2=0 $Y2=0
cc_402 N_A_832_55#_c_580_n N_A_646_74#_c_705_n 0.00779936f $X=5.055 $Y=1.13
+ $X2=0 $Y2=0
cc_403 N_A_832_55#_c_581_n N_A_646_74#_c_705_n 0.005029f $X=5.34 $Y=1.72 $X2=0
+ $Y2=0
cc_404 N_A_832_55#_c_574_n N_A_646_74#_c_706_n 8.98488e-19 $X=4.375 $Y=2.05
+ $X2=0 $Y2=0
cc_405 N_A_832_55#_c_591_n N_A_646_74#_c_706_n 0.00413813f $X=5.34 $Y=1.805
+ $X2=0 $Y2=0
cc_406 N_A_832_55#_c_581_n N_A_646_74#_c_706_n 0.0102417f $X=5.34 $Y=1.72 $X2=0
+ $Y2=0
cc_407 N_A_832_55#_c_574_n N_A_646_74#_c_708_n 3.76298e-19 $X=4.375 $Y=2.05
+ $X2=0 $Y2=0
cc_408 N_A_832_55#_c_574_n N_A_646_74#_c_713_n 0.0177403f $X=4.375 $Y=2.05 $X2=0
+ $Y2=0
cc_409 N_A_832_55#_c_584_n N_A_646_74#_c_713_n 0.0043602f $X=4.39 $Y=2.465 $X2=0
+ $Y2=0
cc_410 N_A_832_55#_c_587_n N_A_646_74#_c_713_n 0.0488981f $X=5.095 $Y=2.24 $X2=0
+ $Y2=0
cc_411 N_A_832_55#_c_591_n N_A_646_74#_c_713_n 0.0112763f $X=5.34 $Y=1.805 $X2=0
+ $Y2=0
cc_412 N_A_832_55#_c_574_n N_A_646_74#_c_709_n 0.0034961f $X=4.375 $Y=2.05 $X2=0
+ $Y2=0
cc_413 N_A_832_55#_c_580_n N_A_646_74#_c_709_n 0.00565954f $X=5.055 $Y=1.13
+ $X2=0 $Y2=0
cc_414 N_A_832_55#_c_581_n N_A_646_74#_c_709_n 0.0295736f $X=5.34 $Y=1.72 $X2=0
+ $Y2=0
cc_415 N_A_832_55#_M1004_g N_RESET_B_c_793_n 0.0196532f $X=6.205 $Y=0.74
+ $X2=-0.19 $Y2=-0.245
cc_416 N_A_832_55#_c_578_n N_RESET_B_c_793_n 0.00328558f $X=5.01 $Y=0.515
+ $X2=-0.19 $Y2=-0.245
cc_417 N_A_832_55#_c_585_n N_RESET_B_c_794_n 0.0292706f $X=6.195 $Y=1.765 $X2=0
+ $Y2=0
cc_418 N_A_832_55#_M1004_g N_RESET_B_c_794_n 0.00317376f $X=6.205 $Y=0.74 $X2=0
+ $Y2=0
cc_419 N_A_832_55#_c_588_n N_RESET_B_c_794_n 0.00643705f $X=5.42 $Y=2.815 $X2=0
+ $Y2=0
cc_420 N_A_832_55#_c_589_n N_RESET_B_c_794_n 0.0155076f $X=6.05 $Y=1.805 $X2=0
+ $Y2=0
cc_421 N_A_832_55#_c_579_n N_RESET_B_c_794_n 0.00259866f $X=6.22 $Y=1.465 $X2=0
+ $Y2=0
cc_422 N_A_832_55#_c_591_n N_RESET_B_c_794_n 0.0109253f $X=5.34 $Y=1.805 $X2=0
+ $Y2=0
cc_423 N_A_832_55#_c_581_n N_RESET_B_c_794_n 0.00138999f $X=5.34 $Y=1.72 $X2=0
+ $Y2=0
cc_424 N_A_832_55#_c_582_n N_RESET_B_c_794_n 0.0242766f $X=6.645 $Y=1.532 $X2=0
+ $Y2=0
cc_425 N_A_832_55#_M1004_g N_RESET_B_c_795_n 0.00137679f $X=6.205 $Y=0.74 $X2=0
+ $Y2=0
cc_426 N_A_832_55#_c_589_n N_RESET_B_c_795_n 0.0187724f $X=6.05 $Y=1.805 $X2=0
+ $Y2=0
cc_427 N_A_832_55#_c_579_n N_RESET_B_c_795_n 0.0153318f $X=6.22 $Y=1.465 $X2=0
+ $Y2=0
cc_428 N_A_832_55#_c_591_n N_RESET_B_c_795_n 0.0128485f $X=5.34 $Y=1.805 $X2=0
+ $Y2=0
cc_429 N_A_832_55#_c_581_n N_RESET_B_c_795_n 0.0283699f $X=5.34 $Y=1.72 $X2=0
+ $Y2=0
cc_430 N_A_832_55#_c_582_n N_RESET_B_c_795_n 9.94568e-19 $X=6.645 $Y=1.532 $X2=0
+ $Y2=0
cc_431 N_A_832_55#_c_587_n N_VPWR_M1005_d 0.00682474f $X=5.095 $Y=2.24 $X2=0
+ $Y2=0
cc_432 N_A_832_55#_c_589_n N_VPWR_M1014_d 0.00304484f $X=6.05 $Y=1.805 $X2=0
+ $Y2=0
cc_433 N_A_832_55#_c_579_n N_VPWR_M1014_d 2.57397e-19 $X=6.22 $Y=1.465 $X2=0
+ $Y2=0
cc_434 N_A_832_55#_c_585_n N_VPWR_c_831_n 0.00735548f $X=6.195 $Y=1.765 $X2=0
+ $Y2=0
cc_435 N_A_832_55#_c_589_n N_VPWR_c_831_n 0.0222109f $X=6.05 $Y=1.805 $X2=0
+ $Y2=0
cc_436 N_A_832_55#_c_579_n N_VPWR_c_831_n 0.00107067f $X=6.22 $Y=1.465 $X2=0
+ $Y2=0
cc_437 N_A_832_55#_c_591_n N_VPWR_c_831_n 0.0360219f $X=5.34 $Y=1.805 $X2=0
+ $Y2=0
cc_438 N_A_832_55#_c_586_n N_VPWR_c_833_n 0.00622993f $X=6.66 $Y=1.765 $X2=0
+ $Y2=0
cc_439 N_A_832_55#_c_584_n N_VPWR_c_836_n 0.00415318f $X=4.39 $Y=2.465 $X2=0
+ $Y2=0
cc_440 N_A_832_55#_c_588_n N_VPWR_c_837_n 0.014552f $X=5.42 $Y=2.815 $X2=0 $Y2=0
cc_441 N_A_832_55#_c_585_n N_VPWR_c_838_n 0.00445602f $X=6.195 $Y=1.765 $X2=0
+ $Y2=0
cc_442 N_A_832_55#_c_586_n N_VPWR_c_838_n 0.00461464f $X=6.66 $Y=1.765 $X2=0
+ $Y2=0
cc_443 N_A_832_55#_c_584_n N_VPWR_c_840_n 0.019118f $X=4.39 $Y=2.465 $X2=0 $Y2=0
cc_444 N_A_832_55#_c_587_n N_VPWR_c_840_n 0.0346382f $X=5.095 $Y=2.24 $X2=0
+ $Y2=0
cc_445 N_A_832_55#_c_588_n N_VPWR_c_840_n 0.013255f $X=5.42 $Y=2.815 $X2=0 $Y2=0
cc_446 N_A_832_55#_c_584_n N_VPWR_c_828_n 0.00857361f $X=4.39 $Y=2.465 $X2=0
+ $Y2=0
cc_447 N_A_832_55#_c_585_n N_VPWR_c_828_n 0.00857968f $X=6.195 $Y=1.765 $X2=0
+ $Y2=0
cc_448 N_A_832_55#_c_586_n N_VPWR_c_828_n 0.00911691f $X=6.66 $Y=1.765 $X2=0
+ $Y2=0
cc_449 N_A_832_55#_c_588_n N_VPWR_c_828_n 0.0119791f $X=5.42 $Y=2.815 $X2=0
+ $Y2=0
cc_450 N_A_832_55#_M1004_g N_Q_c_917_n 0.00751183f $X=6.205 $Y=0.74 $X2=0 $Y2=0
cc_451 N_A_832_55#_M1013_g N_Q_c_917_n 0.0126887f $X=6.645 $Y=0.74 $X2=0 $Y2=0
cc_452 N_A_832_55#_c_585_n N_Q_c_921_n 0.00639588f $X=6.195 $Y=1.765 $X2=0 $Y2=0
cc_453 N_A_832_55#_c_586_n N_Q_c_921_n 0.00128588f $X=6.66 $Y=1.765 $X2=0 $Y2=0
cc_454 N_A_832_55#_c_579_n N_Q_c_921_n 0.00644559f $X=6.22 $Y=1.465 $X2=0 $Y2=0
cc_455 N_A_832_55#_c_670_p N_Q_c_921_n 0.0194426f $X=6.555 $Y=1.465 $X2=0 $Y2=0
cc_456 N_A_832_55#_c_582_n N_Q_c_921_n 0.00708538f $X=6.645 $Y=1.532 $X2=0 $Y2=0
cc_457 N_A_832_55#_c_585_n N_Q_c_922_n 0.00759627f $X=6.195 $Y=1.765 $X2=0 $Y2=0
cc_458 N_A_832_55#_M1013_g N_Q_c_918_n 0.014059f $X=6.645 $Y=0.74 $X2=0 $Y2=0
cc_459 N_A_832_55#_c_670_p N_Q_c_918_n 0.00639324f $X=6.555 $Y=1.465 $X2=0 $Y2=0
cc_460 N_A_832_55#_c_582_n N_Q_c_918_n 6.97142e-19 $X=6.645 $Y=1.532 $X2=0 $Y2=0
cc_461 N_A_832_55#_M1004_g N_Q_c_919_n 0.00380194f $X=6.205 $Y=0.74 $X2=0 $Y2=0
cc_462 N_A_832_55#_M1013_g N_Q_c_919_n 6.77247e-19 $X=6.645 $Y=0.74 $X2=0 $Y2=0
cc_463 N_A_832_55#_c_670_p N_Q_c_919_n 0.0276532f $X=6.555 $Y=1.465 $X2=0 $Y2=0
cc_464 N_A_832_55#_c_582_n N_Q_c_919_n 0.00256252f $X=6.645 $Y=1.532 $X2=0 $Y2=0
cc_465 N_A_832_55#_c_586_n N_Q_c_923_n 0.0152824f $X=6.66 $Y=1.765 $X2=0 $Y2=0
cc_466 N_A_832_55#_c_670_p N_Q_c_923_n 0.00639324f $X=6.555 $Y=1.465 $X2=0 $Y2=0
cc_467 N_A_832_55#_c_582_n N_Q_c_923_n 4.77499e-19 $X=6.645 $Y=1.532 $X2=0 $Y2=0
cc_468 N_A_832_55#_M1013_g Q 0.0112569f $X=6.645 $Y=0.74 $X2=0 $Y2=0
cc_469 N_A_832_55#_c_586_n Q 8.88262e-19 $X=6.66 $Y=1.765 $X2=0 $Y2=0
cc_470 N_A_832_55#_c_579_n Q 0.00463998f $X=6.22 $Y=1.465 $X2=0 $Y2=0
cc_471 N_A_832_55#_c_670_p Q 0.0259734f $X=6.555 $Y=1.465 $X2=0 $Y2=0
cc_472 N_A_832_55#_c_582_n Q 0.00802566f $X=6.645 $Y=1.532 $X2=0 $Y2=0
cc_473 N_A_832_55#_c_573_n N_VGND_c_962_n 0.0113457f $X=4.235 $Y=0.9 $X2=0 $Y2=0
cc_474 N_A_832_55#_c_577_n N_VGND_c_962_n 0.00767933f $X=4.375 $Y=0.975 $X2=0
+ $Y2=0
cc_475 N_A_832_55#_c_578_n N_VGND_c_962_n 0.0339917f $X=5.01 $Y=0.515 $X2=0
+ $Y2=0
cc_476 N_A_832_55#_M1004_g N_VGND_c_963_n 0.0060582f $X=6.205 $Y=0.74 $X2=0
+ $Y2=0
cc_477 N_A_832_55#_c_578_n N_VGND_c_963_n 0.0228983f $X=5.01 $Y=0.515 $X2=0
+ $Y2=0
cc_478 N_A_832_55#_c_579_n N_VGND_c_963_n 0.00155541f $X=6.22 $Y=1.465 $X2=0
+ $Y2=0
cc_479 N_A_832_55#_c_582_n N_VGND_c_963_n 2.01415e-19 $X=6.645 $Y=1.532 $X2=0
+ $Y2=0
cc_480 N_A_832_55#_M1013_g N_VGND_c_965_n 0.0119854f $X=6.645 $Y=0.74 $X2=0
+ $Y2=0
cc_481 N_A_832_55#_c_573_n N_VGND_c_968_n 0.0045897f $X=4.235 $Y=0.9 $X2=0 $Y2=0
cc_482 N_A_832_55#_c_578_n N_VGND_c_969_n 0.0183108f $X=5.01 $Y=0.515 $X2=0
+ $Y2=0
cc_483 N_A_832_55#_M1004_g N_VGND_c_970_n 0.00434272f $X=6.205 $Y=0.74 $X2=0
+ $Y2=0
cc_484 N_A_832_55#_M1013_g N_VGND_c_970_n 0.00445602f $X=6.645 $Y=0.74 $X2=0
+ $Y2=0
cc_485 N_A_832_55#_c_573_n N_VGND_c_974_n 0.0044912f $X=4.235 $Y=0.9 $X2=0 $Y2=0
cc_486 N_A_832_55#_M1004_g N_VGND_c_974_n 0.00821554f $X=6.205 $Y=0.74 $X2=0
+ $Y2=0
cc_487 N_A_832_55#_M1013_g N_VGND_c_974_n 0.00860469f $X=6.645 $Y=0.74 $X2=0
+ $Y2=0
cc_488 N_A_832_55#_c_578_n N_VGND_c_974_n 0.0148883f $X=5.01 $Y=0.515 $X2=0
+ $Y2=0
cc_489 N_A_646_74#_M1011_g N_RESET_B_c_793_n 0.0488418f $X=5.225 $Y=0.74
+ $X2=-0.19 $Y2=-0.245
cc_490 N_A_646_74#_c_710_n N_RESET_B_c_794_n 0.0101951f $X=5.195 $Y=1.765 $X2=0
+ $Y2=0
cc_491 N_A_646_74#_M1011_g N_RESET_B_c_794_n 0.0174252f $X=5.225 $Y=0.74 $X2=0
+ $Y2=0
cc_492 N_A_646_74#_c_706_n N_RESET_B_c_794_n 0.0139508f $X=5.105 $Y=1.35 $X2=0
+ $Y2=0
cc_493 N_A_646_74#_M1011_g N_RESET_B_c_795_n 0.00197031f $X=5.225 $Y=0.74 $X2=0
+ $Y2=0
cc_494 N_A_646_74#_c_706_n N_RESET_B_c_795_n 3.30164e-19 $X=5.105 $Y=1.35 $X2=0
+ $Y2=0
cc_495 N_A_646_74#_c_713_n N_VPWR_M1005_d 0.00182387f $X=4.66 $Y=1.845 $X2=0
+ $Y2=0
cc_496 N_A_646_74#_c_710_n N_VPWR_c_837_n 0.00445602f $X=5.195 $Y=1.765 $X2=0
+ $Y2=0
cc_497 N_A_646_74#_c_710_n N_VPWR_c_840_n 0.00527389f $X=5.195 $Y=1.765 $X2=0
+ $Y2=0
cc_498 N_A_646_74#_c_710_n N_VPWR_c_828_n 0.00859441f $X=5.195 $Y=1.765 $X2=0
+ $Y2=0
cc_499 N_A_646_74#_M1011_g N_VGND_c_962_n 0.00376858f $X=5.225 $Y=0.74 $X2=0
+ $Y2=0
cc_500 N_A_646_74#_M1011_g N_VGND_c_969_n 0.00332301f $X=5.225 $Y=0.74 $X2=0
+ $Y2=0
cc_501 N_A_646_74#_M1011_g N_VGND_c_974_n 0.00495797f $X=5.225 $Y=0.74 $X2=0
+ $Y2=0
cc_502 N_RESET_B_c_794_n N_VPWR_c_831_n 0.00735548f $X=5.645 $Y=1.765 $X2=0
+ $Y2=0
cc_503 N_RESET_B_c_794_n N_VPWR_c_837_n 0.00445602f $X=5.645 $Y=1.765 $X2=0
+ $Y2=0
cc_504 N_RESET_B_c_794_n N_VPWR_c_828_n 0.00857909f $X=5.645 $Y=1.765 $X2=0
+ $Y2=0
cc_505 N_RESET_B_c_793_n N_Q_c_919_n 5.47188e-19 $X=5.615 $Y=1.22 $X2=0 $Y2=0
cc_506 N_RESET_B_c_793_n N_VGND_c_963_n 0.0123659f $X=5.615 $Y=1.22 $X2=0 $Y2=0
cc_507 N_RESET_B_c_794_n N_VGND_c_963_n 5.97749e-19 $X=5.645 $Y=1.765 $X2=0
+ $Y2=0
cc_508 N_RESET_B_c_795_n N_VGND_c_963_n 0.00734321f $X=5.675 $Y=1.385 $X2=0
+ $Y2=0
cc_509 N_RESET_B_c_793_n N_VGND_c_969_n 0.00461464f $X=5.615 $Y=1.22 $X2=0 $Y2=0
cc_510 N_RESET_B_c_793_n N_VGND_c_974_n 0.00909661f $X=5.615 $Y=1.22 $X2=0 $Y2=0
cc_511 N_VPWR_c_831_n N_Q_c_922_n 0.0290824f $X=5.92 $Y=2.145 $X2=0 $Y2=0
cc_512 N_VPWR_c_833_n N_Q_c_922_n 0.0321183f $X=6.92 $Y=2.305 $X2=0 $Y2=0
cc_513 N_VPWR_c_838_n N_Q_c_922_n 0.0145938f $X=6.755 $Y=3.33 $X2=0 $Y2=0
cc_514 N_VPWR_c_828_n N_Q_c_922_n 0.0120466f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_515 N_VPWR_M1020_s N_Q_c_923_n 0.00406667f $X=6.735 $Y=1.84 $X2=0 $Y2=0
cc_516 N_VPWR_c_833_n N_Q_c_923_n 0.0250012f $X=6.92 $Y=2.305 $X2=0 $Y2=0
cc_517 N_Q_c_918_n N_VGND_M1013_s 0.00451672f $X=6.845 $Y=1.045 $X2=0 $Y2=0
cc_518 N_Q_c_917_n N_VGND_c_963_n 0.0236416f $X=6.42 $Y=0.515 $X2=0 $Y2=0
cc_519 N_Q_c_917_n N_VGND_c_965_n 0.0173003f $X=6.42 $Y=0.515 $X2=0 $Y2=0
cc_520 N_Q_c_918_n N_VGND_c_965_n 0.0262685f $X=6.845 $Y=1.045 $X2=0 $Y2=0
cc_521 N_Q_c_917_n N_VGND_c_970_n 0.0145221f $X=6.42 $Y=0.515 $X2=0 $Y2=0
cc_522 N_Q_c_917_n N_VGND_c_974_n 0.0119308f $X=6.42 $Y=0.515 $X2=0 $Y2=0
