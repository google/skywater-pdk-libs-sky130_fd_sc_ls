* NGSPICE file created from sky130_fd_sc_ls__dlygate4sd3_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dlygate4sd3_1 A VGND VNB VPB VPWR X
M1000 VGND a_289_74# a_405_138# VNB nshort w=420000u l=500000u
+  ad=3.935e+11p pd=3.79e+06u as=1.092e+11p ps=1.36e+06u
M1001 VPWR a_289_74# a_405_138# VPB phighvt w=1e+06u l=500000u
+  ad=6.905e+11p pd=5.7e+06u as=2.6e+11p ps=2.52e+06u
M1002 VPWR A a_28_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1003 a_289_74# a_28_74# VPWR VPB phighvt w=1e+06u l=500000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1004 X a_405_138# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1005 VGND A a_28_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1006 X a_405_138# VGND VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1007 a_289_74# a_28_74# VGND VNB nshort w=420000u l=500000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
.ends

