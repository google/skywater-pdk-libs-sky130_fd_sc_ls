* File: sky130_fd_sc_ls__o2bb2a_2.spice
* Created: Fri Aug 28 13:50:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o2bb2a_2.pex.spice"
.subckt sky130_fd_sc_ls__o2bb2a_2  VNB VPB B1 B2 A2_N A1_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1_N	A1_N
* A2_N	A2_N
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_B1_M1011_g N_A_27_74#_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1012 N_A_27_74#_M1012_d N_B2_M1012_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1009 N_A_201_392#_M1009_d N_A_270_48#_M1009_g N_A_27_74#_M1012_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1
+ R=4.93333 SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 A_500_74# N_A2_N_M1006_g N_A_270_48#_M1006_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1010 N_VGND_M1010_d N_A1_N_M1010_g A_500_74# VNB NSHORT L=0.15 W=0.64
+ AD=0.134771 AS=0.0768 PD=1.0713 PS=0.88 NRD=3.744 NRS=12.18 M=1 R=4.26667
+ SA=75000.6 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1003 N_X_M1003_d N_A_201_392#_M1003_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.155829 PD=1.02 PS=1.2387 NRD=0 NRS=18.648 M=1 R=4.93333
+ SA=75001 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1003_d N_A_201_392#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 A_117_392# N_B1_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1001 N_A_201_392#_M1001_d N_B2_M1001_g A_117_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.18 AS=0.135 PD=1.36 PS=1.27 NRD=13.7703 NRS=15.7403 M=1 R=6.66667
+ SA=75000.6 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A_270_48#_M1002_g N_A_201_392#_M1001_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.275367 AS=0.18 PD=1.71739 PS=1.36 NRD=21.6503 NRS=1.9503 M=1
+ R=6.66667 SA=75001.1 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_270_48#_M1000_d N_A2_N_M1000_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1638 AS=0.231308 PD=1.23 PS=1.44261 NRD=12.8838 NRS=51.6731 M=1
+ R=5.6 SA=75001.8 SB=75001.9 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_A1_N_M1004_g N_A_270_48#_M1000_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.274746 AS=0.1638 PD=1.53857 PS=1.23 NRD=63.8083 NRS=12.8838 M=1
+ R=5.6 SA=75002.3 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1005 N_X_M1005_d N_A_201_392#_M1005_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.366329 PD=1.42 PS=2.05143 NRD=1.7533 NRS=28.1316 M=1 R=7.46667
+ SA=75002.4 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1008 N_X_M1005_d N_A_201_392#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.8 SB=75000.2 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__o2bb2a_2.pxi.spice"
*
.ends
*
*
