# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__mux2i_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__mux2i_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.180000 1.315000 1.550000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 1.430000 3.235000 1.775000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.804000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.430000 4.675000 1.840000 ;
        RECT 4.350000 1.840000 5.810000 2.010000 ;
        RECT 5.480000 1.350000 5.810000 1.840000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  2.040950 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 2.910000 0.425000 ;
        RECT 0.085000 0.425000 0.450000 1.010000 ;
        RECT 0.085000 1.010000 0.255000 1.820000 ;
        RECT 0.085000 1.820000 0.445000 1.945000 ;
        RECT 0.085000 1.945000 2.845000 2.115000 ;
        RECT 0.085000 2.115000 0.445000 2.980000 ;
        RECT 2.580000 0.425000 2.910000 0.580000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.615000  2.285000 4.005000 2.340000 ;
      RECT 0.615000  2.340000 3.185000 2.455000 ;
      RECT 0.615000  2.455000 0.945000 2.980000 ;
      RECT 0.640000  0.595000 2.410000 0.750000 ;
      RECT 0.640000  0.750000 5.115000 0.765000 ;
      RECT 0.640000  0.765000 0.970000 1.010000 ;
      RECT 1.685000  2.625000 5.090000 2.680000 ;
      RECT 1.685000  2.680000 3.525000 2.795000 ;
      RECT 1.685000  2.795000 2.395000 2.955000 ;
      RECT 1.740000  0.935000 2.070000 1.090000 ;
      RECT 1.740000  1.090000 4.030000 1.260000 ;
      RECT 2.240000  0.765000 5.115000 0.830000 ;
      RECT 2.240000  0.830000 3.250000 0.920000 ;
      RECT 3.015000  2.010000 4.005000 2.285000 ;
      RECT 3.075000  2.965000 3.470000 3.245000 ;
      RECT 3.080000  0.660000 5.115000 0.750000 ;
      RECT 3.140000  0.085000 3.470000 0.490000 ;
      RECT 3.355000  2.510000 5.090000 2.625000 ;
      RECT 3.650000  1.000000 4.030000 1.090000 ;
      RECT 4.210000  0.085000 4.555000 0.490000 ;
      RECT 4.210000  2.850000 4.555000 3.245000 ;
      RECT 4.735000  0.500000 5.115000 0.660000 ;
      RECT 4.760000  2.180000 5.090000 2.510000 ;
      RECT 4.760000  2.680000 5.090000 2.980000 ;
      RECT 4.910000  1.010000 6.150000 1.180000 ;
      RECT 4.910000  1.180000 5.240000 1.670000 ;
      RECT 5.260000  2.180000 5.590000 3.245000 ;
      RECT 5.285000  0.085000 5.615000 0.840000 ;
      RECT 5.795000  0.570000 6.150000 1.010000 ;
      RECT 5.795000  2.180000 6.150000 2.860000 ;
      RECT 5.980000  1.180000 6.150000 2.180000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_ls__mux2i_2
END LIBRARY
