* File: sky130_fd_sc_ls__buf_2.spice
* Created: Wed Sep  2 10:56:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__buf_2.pex.spice"
.subckt sky130_fd_sc_ls__buf_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_21_260#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A_21_260#_M1005_g N_X_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.166607 AS=0.1036 PD=1.25478 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1003 N_A_21_260#_M1003_d N_A_M1003_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1824 AS=0.144093 PD=1.85 PS=1.08522 NRD=0 NRS=14.988 M=1 R=4.26667
+ SA=75001.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_X_M1000_d N_A_21_260#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.756 PD=1.42 PS=3.59 NRD=1.7533 NRS=46.3147 M=1 R=7.46667
+ SA=75000.6 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1002 N_X_M1000_d N_A_21_260#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.222098 PD=1.42 PS=1.59019 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1004 N_A_21_260#_M1004_d N_A_M1004_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.32 AS=0.198302 PD=2.64 PS=1.41981 NRD=3.9203 NRS=19.6803 M=1 R=6.66667
+ SA=75001.6 SB=75000.2 A=0.15 P=2.3 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_ls__buf_2.pxi.spice"
*
.ends
*
*
