* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_313_74# A1 a_441_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 X a_441_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 VPWR A1 a_27_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_441_74# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 VPWR A3 a_27_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND A4 a_121_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 a_27_392# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_121_74# A3 a_199_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 X a_441_74# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 VPWR a_441_74# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X10 a_199_74# A2 a_313_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X11 a_27_392# B1 a_441_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND a_441_74# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 a_27_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends
