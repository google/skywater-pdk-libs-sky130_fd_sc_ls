* NGSPICE file created from sky130_fd_sc_ls__a22o_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 VPWR A2 a_388_368# VPB phighvt w=1e+06u l=150000u
+  ad=1.0048e+12p pd=8.36e+06u as=6.7e+11p ps=5.34e+06u
M1001 a_81_48# B1 a_388_368# VPB phighvt w=1e+06u l=150000u
+  ad=3.5e+11p pd=2.7e+06u as=0p ps=0u
M1002 X a_81_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1003 a_388_368# B2 a_81_48# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_304_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=4.218e+11p pd=4.1e+06u as=6.808e+11p ps=6.28e+06u
M1005 VPWR a_81_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_491_74# B1 a_81_48# VNB nshort w=740000u l=150000u
+  ad=1.85e+11p pd=1.98e+06u as=2.59e+11p ps=2.18e+06u
M1007 a_81_48# A1 a_304_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_81_48# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1009 a_388_368# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B2 a_491_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_81_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

