* File: sky130_fd_sc_ls__einvp_4.pxi.spice
* Created: Wed Sep  2 11:07:18 2020
* 
x_PM_SKY130_FD_SC_LS__EINVP_4%A N_A_M1002_g N_A_c_120_n N_A_M1000_g N_A_M1005_g
+ N_A_c_121_n N_A_M1008_g N_A_c_122_n N_A_M1009_g N_A_M1014_g N_A_c_114_n
+ N_A_c_115_n N_A_c_116_n N_A_c_125_n N_A_M1013_g N_A_M1016_g N_A_c_118_n A A A
+ N_A_c_119_n PM_SKY130_FD_SC_LS__EINVP_4%A
x_PM_SKY130_FD_SC_LS__EINVP_4%A_473_323# N_A_473_323#_M1015_s
+ N_A_473_323#_M1004_s N_A_473_323#_c_216_n N_A_473_323#_M1003_g
+ N_A_473_323#_c_204_n N_A_473_323#_c_205_n N_A_473_323#_c_219_n
+ N_A_473_323#_M1007_g N_A_473_323#_c_206_n N_A_473_323#_c_221_n
+ N_A_473_323#_M1011_g N_A_473_323#_c_207_n N_A_473_323#_c_223_n
+ N_A_473_323#_M1012_g N_A_473_323#_c_208_n N_A_473_323#_c_209_n
+ N_A_473_323#_c_210_n N_A_473_323#_c_211_n N_A_473_323#_c_212_n
+ N_A_473_323#_c_213_n N_A_473_323#_c_228_n N_A_473_323#_c_214_n
+ N_A_473_323#_c_215_n PM_SKY130_FD_SC_LS__EINVP_4%A_473_323#
x_PM_SKY130_FD_SC_LS__EINVP_4%TE N_TE_c_317_n N_TE_M1001_g N_TE_c_318_n
+ N_TE_c_319_n N_TE_c_320_n N_TE_M1006_g N_TE_c_321_n N_TE_c_322_n N_TE_M1010_g
+ N_TE_c_323_n N_TE_c_324_n N_TE_M1017_g N_TE_c_325_n N_TE_c_326_n N_TE_M1015_g
+ N_TE_c_333_n N_TE_M1004_g N_TE_c_327_n N_TE_c_328_n N_TE_c_329_n TE
+ N_TE_c_331_n N_TE_c_332_n PM_SKY130_FD_SC_LS__EINVP_4%TE
x_PM_SKY130_FD_SC_LS__EINVP_4%A_27_368# N_A_27_368#_M1000_d N_A_27_368#_M1008_d
+ N_A_27_368#_M1013_d N_A_27_368#_M1007_s N_A_27_368#_M1012_s
+ N_A_27_368#_c_418_n N_A_27_368#_c_419_n N_A_27_368#_c_420_n
+ N_A_27_368#_c_477_p N_A_27_368#_c_421_n N_A_27_368#_c_422_n
+ N_A_27_368#_c_423_n N_A_27_368#_c_417_n N_A_27_368#_c_425_n
+ N_A_27_368#_c_426_n N_A_27_368#_c_427_n N_A_27_368#_c_428_n
+ N_A_27_368#_c_467_n PM_SKY130_FD_SC_LS__EINVP_4%A_27_368#
x_PM_SKY130_FD_SC_LS__EINVP_4%Z N_Z_M1002_s N_Z_M1014_s N_Z_M1000_s N_Z_M1009_s
+ N_Z_c_513_n N_Z_c_508_n N_Z_c_509_n N_Z_c_523_n N_Z_c_527_n N_Z_c_510_n
+ N_Z_c_537_n N_Z_c_541_n N_Z_c_511_n Z PM_SKY130_FD_SC_LS__EINVP_4%Z
x_PM_SKY130_FD_SC_LS__EINVP_4%VPWR N_VPWR_M1003_d N_VPWR_M1011_d N_VPWR_M1004_d
+ N_VPWR_c_570_n N_VPWR_c_571_n N_VPWR_c_572_n N_VPWR_c_573_n VPWR
+ N_VPWR_c_574_n N_VPWR_c_575_n N_VPWR_c_576_n N_VPWR_c_577_n N_VPWR_c_578_n
+ N_VPWR_c_569_n PM_SKY130_FD_SC_LS__EINVP_4%VPWR
x_PM_SKY130_FD_SC_LS__EINVP_4%A_27_74# N_A_27_74#_M1002_d N_A_27_74#_M1005_d
+ N_A_27_74#_M1016_d N_A_27_74#_M1006_s N_A_27_74#_M1017_s N_A_27_74#_c_631_n
+ N_A_27_74#_c_632_n N_A_27_74#_c_633_n N_A_27_74#_c_701_n N_A_27_74#_c_634_n
+ N_A_27_74#_c_635_n N_A_27_74#_c_636_n N_A_27_74#_c_637_n N_A_27_74#_c_638_n
+ N_A_27_74#_c_639_n N_A_27_74#_c_640_n N_A_27_74#_c_641_n N_A_27_74#_c_642_n
+ PM_SKY130_FD_SC_LS__EINVP_4%A_27_74#
x_PM_SKY130_FD_SC_LS__EINVP_4%VGND N_VGND_M1001_d N_VGND_M1010_d N_VGND_M1015_d
+ N_VGND_c_727_n N_VGND_c_728_n N_VGND_c_729_n N_VGND_c_730_n N_VGND_c_731_n
+ N_VGND_c_732_n VGND N_VGND_c_733_n N_VGND_c_734_n N_VGND_c_735_n
+ N_VGND_c_736_n PM_SKY130_FD_SC_LS__EINVP_4%VGND
cc_1 VNB N_A_M1002_g 0.0326264f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_M1005_g 0.0244962f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_A_M1014_g 0.0240943f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.74
cc_4 VNB N_A_c_114_n 0.0109911f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.425
cc_5 VNB N_A_c_115_n 0.0589745f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.425
cc_6 VNB N_A_c_116_n 0.0114766f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.675
cc_7 VNB N_A_M1016_g 0.0243622f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_8 VNB N_A_c_118_n 0.00907757f $X=-0.19 $Y=-0.245 $X2=1.967 $Y2=1.425
cc_9 VNB N_A_c_119_n 0.016914f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_10 VNB N_A_473_323#_c_204_n 0.00778029f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_11 VNB N_A_473_323#_c_205_n 0.00498537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_473_323#_c_206_n 0.00674479f $X=-0.19 $Y=-0.245 $X2=1.505
+ $Y2=1.765
cc_13 VNB N_A_473_323#_c_207_n 0.00696655f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.74
cc_14 VNB N_A_473_323#_c_208_n 0.0177303f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.675
cc_15 VNB N_A_473_323#_c_209_n 0.00344292f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_16 VNB N_A_473_323#_c_210_n 0.00344284f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_17 VNB N_A_473_323#_c_211_n 0.00344292f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=1.35
cc_18 VNB N_A_473_323#_c_212_n 0.00909917f $X=-0.19 $Y=-0.245 $X2=1.967
+ $Y2=1.425
cc_19 VNB N_A_473_323#_c_213_n 0.00914505f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_20 VNB N_A_473_323#_c_214_n 2.54189e-19 $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.515
cc_21 VNB N_A_473_323#_c_215_n 0.00653231f $X=-0.19 $Y=-0.245 $X2=1.265
+ $Y2=1.557
cc_22 VNB N_TE_c_317_n 0.018325f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_23 VNB N_TE_c_318_n 0.0166678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_TE_c_319_n 0.00643851f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.765
cc_25 VNB N_TE_c_320_n 0.0180464f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_26 VNB N_TE_c_321_n 0.0105119f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_27 VNB N_TE_c_322_n 0.0180464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_TE_c_323_n 0.0166678f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_29 VNB N_TE_c_324_n 0.0232894f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.4
cc_30 VNB N_TE_c_325_n 0.0497754f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.74
cc_31 VNB N_TE_c_326_n 0.0245033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_TE_c_327_n 0.00411221f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_33 VNB N_TE_c_328_n 0.00411221f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_34 VNB N_TE_c_329_n 0.00411221f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=1.35
cc_35 VNB TE 0.0246417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_TE_c_331_n 0.0794645f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_37 VNB N_TE_c_332_n 0.00245723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_368#_c_417_n 0.00443147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Z_c_508_n 0.00388917f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.74
cc_40 VNB N_Z_c_509_n 0.00320239f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.74
cc_41 VNB N_Z_c_510_n 0.00363957f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_42 VNB N_Z_c_511_n 9.85474e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_43 VNB N_VPWR_c_569_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_44 VNB N_A_27_74#_c_631_n 0.0302158f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.35
cc_45 VNB N_A_27_74#_c_632_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.74
cc_46 VNB N_A_27_74#_c_633_n 0.00971634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_74#_c_634_n 0.00484762f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.765
cc_48 VNB N_A_27_74#_c_635_n 0.00195492f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_49 VNB N_A_27_74#_c_636_n 0.00396969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_27_74#_c_637_n 0.00466188f $X=-0.19 $Y=-0.245 $X2=1.967 $Y2=1.425
cc_51 VNB N_A_27_74#_c_638_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_52 VNB N_A_27_74#_c_639_n 0.0078054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_27_74#_c_640_n 0.00962339f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.557
cc_54 VNB N_A_27_74#_c_641_n 0.00244677f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_55 VNB N_A_27_74#_c_642_n 0.00200315f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.557
cc_56 VNB N_VGND_c_727_n 0.011008f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.765
cc_57 VNB N_VGND_c_728_n 0.0114288f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.4
cc_58 VNB N_VGND_c_729_n 0.0166826f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.35
cc_59 VNB N_VGND_c_730_n 0.0377021f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.74
cc_60 VNB N_VGND_c_731_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.425
cc_61 VNB N_VGND_c_732_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.5
cc_62 VNB N_VGND_c_733_n 0.0627368f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_63 VNB N_VGND_c_734_n 0.0334841f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_64 VNB N_VGND_c_735_n 0.00634377f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_65 VNB N_VGND_c_736_n 0.330625f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_66 VPB N_A_c_120_n 0.0189957f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_67 VPB N_A_c_121_n 0.0153915f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_68 VPB N_A_c_122_n 0.0150747f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=1.765
cc_69 VPB N_A_c_115_n 0.0378309f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.425
cc_70 VPB N_A_c_116_n 7.31788e-19 $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.675
cc_71 VPB N_A_c_125_n 0.0208846f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.765
cc_72 VPB N_A_c_119_n 0.0155975f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_73 VPB N_A_473_323#_c_216_n 0.0154576f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_74 VPB N_A_473_323#_c_204_n 0.00874663f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_75 VPB N_A_473_323#_c_205_n 0.00382842f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_473_323#_c_219_n 0.0154531f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_77 VPB N_A_473_323#_c_206_n 0.00675749f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=1.765
cc_78 VPB N_A_473_323#_c_221_n 0.014779f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=2.4
cc_79 VPB N_A_473_323#_c_207_n 0.00715532f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=0.74
cc_80 VPB N_A_473_323#_c_223_n 0.0185103f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=1.425
cc_81 VPB N_A_473_323#_c_208_n 0.0209585f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.675
cc_82 VPB N_A_473_323#_c_209_n 0.00167153f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_83 VPB N_A_473_323#_c_210_n 0.00167153f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_84 VPB N_A_473_323#_c_211_n 0.00167153f $X=-0.19 $Y=1.66 $X2=1.995 $Y2=1.35
cc_85 VPB N_A_473_323#_c_228_n 0.0990623f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_473_323#_c_214_n 0.0226371f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_87 VPB N_TE_c_333_n 0.0211109f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.5
cc_88 VPB N_TE_c_331_n 0.0107883f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_89 VPB N_A_27_368#_c_418_n 0.0366851f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=1.35
cc_90 VPB N_A_27_368#_c_419_n 0.00269852f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=1.425
cc_91 VPB N_A_27_368#_c_420_n 0.00988933f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.425
cc_92 VPB N_A_27_368#_c_421_n 0.0051269f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_93 VPB N_A_27_368#_c_422_n 2.81009e-19 $X=-0.19 $Y=1.66 $X2=1.967 $Y2=1.425
cc_94 VPB N_A_27_368#_c_423_n 0.00577788f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_95 VPB N_A_27_368#_c_417_n 0.0014986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_27_368#_c_425_n 0.00241809f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_97 VPB N_A_27_368#_c_426_n 0.00701f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_98 VPB N_A_27_368#_c_427_n 0.00237617f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_99 VPB N_A_27_368#_c_428_n 0.00181992f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_100 VPB N_Z_c_510_n 0.00151522f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_101 VPB N_VPWR_c_570_n 0.00777124f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_102 VPB N_VPWR_c_571_n 0.00525442f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=1.35
cc_103 VPB N_VPWR_c_572_n 0.0106521f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=1.425
cc_104 VPB N_VPWR_c_573_n 0.0560624f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.5
cc_105 VPB N_VPWR_c_574_n 0.061632f $X=-0.19 $Y=1.66 $X2=1.995 $Y2=0.74
cc_106 VPB N_VPWR_c_575_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_107 VPB N_VPWR_c_576_n 0.0448319f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_108 VPB N_VPWR_c_577_n 0.0047791f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_109 VPB N_VPWR_c_578_n 0.00479483f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_110 VPB N_VPWR_c_569_n 0.0888383f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_111 N_A_c_125_n N_A_473_323#_c_216_n 0.0217109f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_112 N_A_c_116_n N_A_473_323#_c_205_n 0.00536472f $X=1.955 $Y=1.675 $X2=0
+ $Y2=0
cc_113 N_A_M1016_g N_TE_c_317_n 0.0114134f $X=1.995 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_114 N_A_c_118_n N_TE_c_319_n 0.0114134f $X=1.967 $Y=1.425 $X2=0 $Y2=0
cc_115 N_A_c_120_n N_A_27_368#_c_418_n 0.0106095f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_116 N_A_c_121_n N_A_27_368#_c_418_n 6.12807e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A_c_119_n N_A_27_368#_c_418_n 0.025553f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_118 N_A_c_120_n N_A_27_368#_c_419_n 0.0114142f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A_c_121_n N_A_27_368#_c_419_n 0.0141012f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A_c_120_n N_A_27_368#_c_420_n 0.00253309f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A_c_122_n N_A_27_368#_c_421_n 0.0130187f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A_c_125_n N_A_27_368#_c_421_n 0.013793f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A_c_125_n N_A_27_368#_c_422_n 0.00592136f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A_c_116_n N_A_27_368#_c_417_n 0.00117873f $X=1.955 $Y=1.675 $X2=0 $Y2=0
cc_125 N_A_c_125_n N_A_27_368#_c_417_n 4.15888e-19 $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A_c_118_n N_A_27_368#_c_417_n 2.49919e-19 $X=1.967 $Y=1.425 $X2=0 $Y2=0
cc_127 N_A_M1005_g N_Z_c_513_n 0.00602688f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A_M1014_g N_Z_c_513_n 6.18096e-19 $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A_M1005_g N_Z_c_508_n 0.00952207f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_M1014_g N_Z_c_508_n 0.0176613f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A_c_115_n N_Z_c_508_n 0.00437201f $X=1.595 $Y=1.425 $X2=0 $Y2=0
cc_132 N_A_c_119_n N_Z_c_508_n 0.0367038f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A_M1002_g N_Z_c_509_n 0.00234945f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A_M1005_g N_Z_c_509_n 0.0026663f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_c_115_n N_Z_c_509_n 0.0039232f $X=1.595 $Y=1.425 $X2=0 $Y2=0
cc_136 N_A_c_119_n N_Z_c_509_n 0.0276331f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A_c_121_n N_Z_c_523_n 0.0122806f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A_c_122_n N_Z_c_523_n 0.0163732f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A_c_115_n N_Z_c_523_n 0.00158442f $X=1.595 $Y=1.425 $X2=0 $Y2=0
cc_140 N_A_c_119_n N_Z_c_523_n 0.0335539f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A_M1016_g N_Z_c_527_n 0.00395262f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A_c_122_n N_Z_c_510_n 0.0017463f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A_M1014_g N_Z_c_510_n 0.00474402f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A_c_114_n N_Z_c_510_n 0.0112863f $X=1.865 $Y=1.425 $X2=0 $Y2=0
cc_145 N_A_c_115_n N_Z_c_510_n 0.00247436f $X=1.595 $Y=1.425 $X2=0 $Y2=0
cc_146 N_A_c_116_n N_Z_c_510_n 0.00743471f $X=1.955 $Y=1.675 $X2=0 $Y2=0
cc_147 N_A_c_125_n N_Z_c_510_n 0.00473315f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A_M1016_g N_Z_c_510_n 0.00156994f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_c_118_n N_Z_c_510_n 0.00294268f $X=1.967 $Y=1.425 $X2=0 $Y2=0
cc_150 N_A_c_119_n N_Z_c_510_n 0.0326257f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_151 N_A_c_121_n N_Z_c_537_n 0.0102998f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A_c_122_n N_Z_c_537_n 5.483e-19 $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A_c_115_n N_Z_c_537_n 0.00166699f $X=1.595 $Y=1.425 $X2=0 $Y2=0
cc_154 N_A_c_119_n N_Z_c_537_n 0.0252536f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_155 N_A_c_122_n N_Z_c_541_n 9.50925e-19 $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_156 N_A_c_125_n N_Z_c_541_n 0.00162804f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A_M1016_g N_Z_c_511_n 0.00512787f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A_c_121_n Z 6.34207e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A_c_122_n Z 0.0103018f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A_c_125_n Z 0.00846074f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A_c_120_n N_VPWR_c_574_n 0.00278262f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A_c_121_n N_VPWR_c_574_n 0.00278271f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_c_122_n N_VPWR_c_574_n 0.00278271f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A_c_125_n N_VPWR_c_574_n 0.00278271f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A_c_120_n N_VPWR_c_569_n 0.0035775f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A_c_121_n N_VPWR_c_569_n 0.00354701f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A_c_122_n N_VPWR_c_569_n 0.00354284f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A_c_125_n N_VPWR_c_569_n 0.00354337f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_169 N_A_M1002_g N_A_27_74#_c_631_n 0.0114672f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A_M1005_g N_A_27_74#_c_631_n 8.28548e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A_c_119_n N_A_27_74#_c_631_n 0.023775f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_172 N_A_M1002_g N_A_27_74#_c_632_n 0.0104643f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A_M1005_g N_A_27_74#_c_632_n 0.0118001f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A_M1002_g N_A_27_74#_c_633_n 0.00282152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A_M1014_g N_A_27_74#_c_634_n 0.00938114f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_M1016_g N_A_27_74#_c_634_n 0.0136901f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A_M1016_g N_A_27_74#_c_635_n 0.0052852f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A_M1016_g N_A_27_74#_c_637_n 0.00392472f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A_M1014_g N_A_27_74#_c_641_n 0.00255335f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A_M1002_g N_VGND_c_733_n 0.00278247f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A_M1005_g N_VGND_c_733_n 0.00278271f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A_M1014_g N_VGND_c_733_n 0.00278271f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A_M1016_g N_VGND_c_733_n 0.00278271f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A_M1002_g N_VGND_c_736_n 0.00357743f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A_M1005_g N_VGND_c_736_n 0.00354959f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_186 N_A_M1014_g N_VGND_c_736_n 0.00354734f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A_M1016_g N_VGND_c_736_n 0.00354573f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A_473_323#_c_204_n N_TE_c_318_n 0.0155566f $X=2.88 $Y=1.69 $X2=0 $Y2=0
cc_189 N_A_473_323#_c_205_n N_TE_c_319_n 0.0155566f $X=2.53 $Y=1.69 $X2=0 $Y2=0
cc_190 N_A_473_323#_c_206_n N_TE_c_321_n 0.0155566f $X=3.33 $Y=1.69 $X2=0 $Y2=0
cc_191 N_A_473_323#_c_207_n N_TE_c_323_n 0.0155566f $X=3.79 $Y=1.69 $X2=0 $Y2=0
cc_192 N_A_473_323#_c_212_n N_TE_c_324_n 0.00176266f $X=4.84 $Y=0.515 $X2=0
+ $Y2=0
cc_193 N_A_473_323#_c_208_n N_TE_c_325_n 0.0155566f $X=4.395 $Y=1.69 $X2=0 $Y2=0
cc_194 N_A_473_323#_c_213_n N_TE_c_325_n 0.0141663f $X=4.7 $Y=1.64 $X2=0 $Y2=0
cc_195 N_A_473_323#_c_214_n N_TE_c_325_n 0.00755084f $X=5.03 $Y=2.815 $X2=0
+ $Y2=0
cc_196 N_A_473_323#_c_215_n N_TE_c_325_n 0.00468311f $X=4.81 $Y=1.13 $X2=0 $Y2=0
cc_197 N_A_473_323#_c_212_n N_TE_c_326_n 0.00812744f $X=4.84 $Y=0.515 $X2=0
+ $Y2=0
cc_198 N_A_473_323#_c_213_n N_TE_c_326_n 0.00267162f $X=4.7 $Y=1.64 $X2=0 $Y2=0
cc_199 N_A_473_323#_c_215_n N_TE_c_326_n 0.00684687f $X=4.81 $Y=1.13 $X2=0 $Y2=0
cc_200 N_A_473_323#_c_228_n N_TE_c_333_n 0.0155957f $X=4.56 $Y=1.805 $X2=0 $Y2=0
cc_201 N_A_473_323#_c_214_n N_TE_c_333_n 0.0155434f $X=5.03 $Y=2.815 $X2=0 $Y2=0
cc_202 N_A_473_323#_c_209_n N_TE_c_327_n 0.0155566f $X=2.955 $Y=1.69 $X2=0 $Y2=0
cc_203 N_A_473_323#_c_210_n N_TE_c_328_n 0.0155566f $X=3.405 $Y=1.69 $X2=0 $Y2=0
cc_204 N_A_473_323#_c_211_n N_TE_c_329_n 0.0155566f $X=3.865 $Y=1.69 $X2=0 $Y2=0
cc_205 N_A_473_323#_c_213_n TE 0.00316442f $X=4.7 $Y=1.64 $X2=0 $Y2=0
cc_206 N_A_473_323#_c_208_n N_TE_c_331_n 0.00388748f $X=4.395 $Y=1.69 $X2=0
+ $Y2=0
cc_207 N_A_473_323#_c_213_n N_TE_c_331_n 0.00182782f $X=4.7 $Y=1.64 $X2=0 $Y2=0
cc_208 N_A_473_323#_c_214_n N_TE_c_331_n 0.00787301f $X=5.03 $Y=2.815 $X2=0
+ $Y2=0
cc_209 N_A_473_323#_c_213_n N_TE_c_332_n 0.0233109f $X=4.7 $Y=1.64 $X2=0 $Y2=0
cc_210 N_A_473_323#_c_214_n N_TE_c_332_n 0.0166084f $X=5.03 $Y=2.815 $X2=0 $Y2=0
cc_211 N_A_473_323#_c_215_n N_TE_c_332_n 0.00191579f $X=4.81 $Y=1.13 $X2=0 $Y2=0
cc_212 N_A_473_323#_c_216_n N_A_27_368#_c_421_n 0.00330015f $X=2.455 $Y=1.765
+ $X2=0 $Y2=0
cc_213 N_A_473_323#_c_216_n N_A_27_368#_c_422_n 0.0128998f $X=2.455 $Y=1.765
+ $X2=0 $Y2=0
cc_214 N_A_473_323#_c_219_n N_A_27_368#_c_422_n 6.58456e-19 $X=2.955 $Y=1.765
+ $X2=0 $Y2=0
cc_215 N_A_473_323#_c_216_n N_A_27_368#_c_423_n 0.00708357f $X=2.455 $Y=1.765
+ $X2=0 $Y2=0
cc_216 N_A_473_323#_c_204_n N_A_27_368#_c_423_n 0.00835418f $X=2.88 $Y=1.69
+ $X2=0 $Y2=0
cc_217 N_A_473_323#_c_205_n N_A_27_368#_c_423_n 0.00225485f $X=2.53 $Y=1.69
+ $X2=0 $Y2=0
cc_218 N_A_473_323#_c_219_n N_A_27_368#_c_423_n 0.00708357f $X=2.955 $Y=1.765
+ $X2=0 $Y2=0
cc_219 N_A_473_323#_c_209_n N_A_27_368#_c_423_n 0.00224311f $X=2.955 $Y=1.69
+ $X2=0 $Y2=0
cc_220 N_A_473_323#_c_216_n N_A_27_368#_c_417_n 5.97842e-19 $X=2.455 $Y=1.765
+ $X2=0 $Y2=0
cc_221 N_A_473_323#_c_205_n N_A_27_368#_c_417_n 0.00229368f $X=2.53 $Y=1.69
+ $X2=0 $Y2=0
cc_222 N_A_473_323#_c_216_n N_A_27_368#_c_425_n 7.85528e-19 $X=2.455 $Y=1.765
+ $X2=0 $Y2=0
cc_223 N_A_473_323#_c_219_n N_A_27_368#_c_425_n 0.0144649f $X=2.955 $Y=1.765
+ $X2=0 $Y2=0
cc_224 N_A_473_323#_c_221_n N_A_27_368#_c_425_n 0.00546622f $X=3.405 $Y=1.765
+ $X2=0 $Y2=0
cc_225 N_A_473_323#_c_206_n N_A_27_368#_c_426_n 0.0010532f $X=3.33 $Y=1.69 $X2=0
+ $Y2=0
cc_226 N_A_473_323#_c_221_n N_A_27_368#_c_426_n 0.00790338f $X=3.405 $Y=1.765
+ $X2=0 $Y2=0
cc_227 N_A_473_323#_c_207_n N_A_27_368#_c_426_n 0.00708959f $X=3.79 $Y=1.69
+ $X2=0 $Y2=0
cc_228 N_A_473_323#_c_223_n N_A_27_368#_c_426_n 0.00764928f $X=3.865 $Y=1.765
+ $X2=0 $Y2=0
cc_229 N_A_473_323#_c_208_n N_A_27_368#_c_426_n 0.00947624f $X=4.395 $Y=1.69
+ $X2=0 $Y2=0
cc_230 N_A_473_323#_c_210_n N_A_27_368#_c_426_n 0.00250839f $X=3.405 $Y=1.69
+ $X2=0 $Y2=0
cc_231 N_A_473_323#_c_211_n N_A_27_368#_c_426_n 0.00249483f $X=3.865 $Y=1.69
+ $X2=0 $Y2=0
cc_232 N_A_473_323#_c_228_n N_A_27_368#_c_426_n 2.10193e-19 $X=4.56 $Y=1.805
+ $X2=0 $Y2=0
cc_233 N_A_473_323#_c_214_n N_A_27_368#_c_426_n 0.0113878f $X=5.03 $Y=2.815
+ $X2=0 $Y2=0
cc_234 N_A_473_323#_c_221_n N_A_27_368#_c_427_n 7.609e-19 $X=3.405 $Y=1.765
+ $X2=0 $Y2=0
cc_235 N_A_473_323#_c_223_n N_A_27_368#_c_427_n 0.0147409f $X=3.865 $Y=1.765
+ $X2=0 $Y2=0
cc_236 N_A_473_323#_c_228_n N_A_27_368#_c_427_n 0.00461458f $X=4.56 $Y=1.805
+ $X2=0 $Y2=0
cc_237 N_A_473_323#_c_214_n N_A_27_368#_c_427_n 0.0774029f $X=5.03 $Y=2.815
+ $X2=0 $Y2=0
cc_238 N_A_473_323#_c_219_n N_A_27_368#_c_467_n 6.19113e-19 $X=2.955 $Y=1.765
+ $X2=0 $Y2=0
cc_239 N_A_473_323#_c_206_n N_A_27_368#_c_467_n 0.00681422f $X=3.33 $Y=1.69
+ $X2=0 $Y2=0
cc_240 N_A_473_323#_c_209_n N_A_27_368#_c_467_n 2.51714e-19 $X=2.955 $Y=1.69
+ $X2=0 $Y2=0
cc_241 N_A_473_323#_c_205_n N_Z_c_510_n 2.19962e-19 $X=2.53 $Y=1.69 $X2=0 $Y2=0
cc_242 N_A_473_323#_c_216_n N_VPWR_c_570_n 0.00657293f $X=2.455 $Y=1.765 $X2=0
+ $Y2=0
cc_243 N_A_473_323#_c_204_n N_VPWR_c_570_n 0.0012088f $X=2.88 $Y=1.69 $X2=0
+ $Y2=0
cc_244 N_A_473_323#_c_219_n N_VPWR_c_570_n 0.00510303f $X=2.955 $Y=1.765 $X2=0
+ $Y2=0
cc_245 N_A_473_323#_c_219_n N_VPWR_c_571_n 6.7385e-19 $X=2.955 $Y=1.765 $X2=0
+ $Y2=0
cc_246 N_A_473_323#_c_221_n N_VPWR_c_571_n 0.0139706f $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_247 N_A_473_323#_c_207_n N_VPWR_c_571_n 9.24379e-19 $X=3.79 $Y=1.69 $X2=0
+ $Y2=0
cc_248 N_A_473_323#_c_223_n N_VPWR_c_571_n 0.00628007f $X=3.865 $Y=1.765 $X2=0
+ $Y2=0
cc_249 N_A_473_323#_c_214_n N_VPWR_c_571_n 2.73444e-19 $X=5.03 $Y=2.815 $X2=0
+ $Y2=0
cc_250 N_A_473_323#_c_214_n N_VPWR_c_573_n 0.0829771f $X=5.03 $Y=2.815 $X2=0
+ $Y2=0
cc_251 N_A_473_323#_c_216_n N_VPWR_c_574_n 0.0044313f $X=2.455 $Y=1.765 $X2=0
+ $Y2=0
cc_252 N_A_473_323#_c_219_n N_VPWR_c_575_n 0.00445602f $X=2.955 $Y=1.765 $X2=0
+ $Y2=0
cc_253 N_A_473_323#_c_221_n N_VPWR_c_575_n 0.00413917f $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_254 N_A_473_323#_c_223_n N_VPWR_c_576_n 0.00445602f $X=3.865 $Y=1.765 $X2=0
+ $Y2=0
cc_255 N_A_473_323#_c_228_n N_VPWR_c_576_n 0.00188351f $X=4.56 $Y=1.805 $X2=0
+ $Y2=0
cc_256 N_A_473_323#_c_214_n N_VPWR_c_576_n 0.0353756f $X=5.03 $Y=2.815 $X2=0
+ $Y2=0
cc_257 N_A_473_323#_c_216_n N_VPWR_c_569_n 0.00853664f $X=2.455 $Y=1.765 $X2=0
+ $Y2=0
cc_258 N_A_473_323#_c_219_n N_VPWR_c_569_n 0.0085805f $X=2.955 $Y=1.765 $X2=0
+ $Y2=0
cc_259 N_A_473_323#_c_221_n N_VPWR_c_569_n 0.00817726f $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_260 N_A_473_323#_c_223_n N_VPWR_c_569_n 0.00862487f $X=3.865 $Y=1.765 $X2=0
+ $Y2=0
cc_261 N_A_473_323#_c_214_n N_VPWR_c_569_n 0.0292986f $X=5.03 $Y=2.815 $X2=0
+ $Y2=0
cc_262 N_A_473_323#_c_205_n N_A_27_74#_c_636_n 0.00422967f $X=2.53 $Y=1.69 $X2=0
+ $Y2=0
cc_263 N_A_473_323#_c_205_n N_A_27_74#_c_637_n 0.00162016f $X=2.53 $Y=1.69 $X2=0
+ $Y2=0
cc_264 N_A_473_323#_c_208_n N_A_27_74#_c_639_n 0.00700874f $X=4.395 $Y=1.69
+ $X2=0 $Y2=0
cc_265 N_A_473_323#_c_210_n N_A_27_74#_c_639_n 0.00416942f $X=3.405 $Y=1.69
+ $X2=0 $Y2=0
cc_266 N_A_473_323#_c_213_n N_A_27_74#_c_639_n 0.0137368f $X=4.7 $Y=1.64 $X2=0
+ $Y2=0
cc_267 N_A_473_323#_c_214_n N_A_27_74#_c_639_n 0.00445757f $X=5.03 $Y=2.815
+ $X2=0 $Y2=0
cc_268 N_A_473_323#_c_212_n N_A_27_74#_c_640_n 0.0785503f $X=4.84 $Y=0.515 $X2=0
+ $Y2=0
cc_269 N_A_473_323#_c_206_n N_A_27_74#_c_642_n 0.0023366f $X=3.33 $Y=1.69 $X2=0
+ $Y2=0
cc_270 N_A_473_323#_c_212_n N_VGND_c_730_n 0.026158f $X=4.84 $Y=0.515 $X2=0
+ $Y2=0
cc_271 N_A_473_323#_c_212_n N_VGND_c_734_n 0.0172412f $X=4.84 $Y=0.515 $X2=0
+ $Y2=0
cc_272 N_A_473_323#_c_212_n N_VGND_c_736_n 0.0142144f $X=4.84 $Y=0.515 $X2=0
+ $Y2=0
cc_273 N_TE_c_319_n N_A_27_368#_c_423_n 6.07857e-19 $X=2.57 $Y=1.3 $X2=0 $Y2=0
cc_274 N_TE_c_321_n N_A_27_368#_c_426_n 6.73874e-19 $X=3.42 $Y=1.3 $X2=0 $Y2=0
cc_275 N_TE_c_323_n N_A_27_368#_c_426_n 2.50455e-19 $X=3.99 $Y=1.3 $X2=0 $Y2=0
cc_276 N_TE_c_327_n N_A_27_368#_c_467_n 2.51631e-19 $X=3.065 $Y=1.3 $X2=0 $Y2=0
cc_277 N_TE_c_333_n N_VPWR_c_573_n 0.00994907f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_278 N_TE_c_331_n N_VPWR_c_573_n 0.00595461f $X=5.255 $Y=1.495 $X2=0 $Y2=0
cc_279 N_TE_c_332_n N_VPWR_c_573_n 0.019603f $X=5.485 $Y=1.465 $X2=0 $Y2=0
cc_280 N_TE_c_333_n N_VPWR_c_576_n 0.00444469f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_281 N_TE_c_333_n N_VPWR_c_569_n 0.00862217f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_282 N_TE_c_317_n N_A_27_74#_c_634_n 0.00348233f $X=2.495 $Y=1.225 $X2=0 $Y2=0
cc_283 N_TE_c_317_n N_A_27_74#_c_635_n 0.011268f $X=2.495 $Y=1.225 $X2=0 $Y2=0
cc_284 N_TE_c_319_n N_A_27_74#_c_635_n 0.00315932f $X=2.57 $Y=1.3 $X2=0 $Y2=0
cc_285 N_TE_c_320_n N_A_27_74#_c_635_n 4.34235e-19 $X=3.065 $Y=1.225 $X2=0 $Y2=0
cc_286 N_TE_c_318_n N_A_27_74#_c_636_n 0.0118714f $X=2.99 $Y=1.3 $X2=0 $Y2=0
cc_287 N_TE_c_319_n N_A_27_74#_c_636_n 0.0069434f $X=2.57 $Y=1.3 $X2=0 $Y2=0
cc_288 N_TE_c_327_n N_A_27_74#_c_636_n 0.00696323f $X=3.065 $Y=1.3 $X2=0 $Y2=0
cc_289 N_TE_c_319_n N_A_27_74#_c_637_n 0.00120269f $X=2.57 $Y=1.3 $X2=0 $Y2=0
cc_290 N_TE_c_317_n N_A_27_74#_c_638_n 4.49351e-19 $X=2.495 $Y=1.225 $X2=0 $Y2=0
cc_291 N_TE_c_320_n N_A_27_74#_c_638_n 0.0125068f $X=3.065 $Y=1.225 $X2=0 $Y2=0
cc_292 N_TE_c_321_n N_A_27_74#_c_638_n 0.00434616f $X=3.42 $Y=1.3 $X2=0 $Y2=0
cc_293 N_TE_c_322_n N_A_27_74#_c_638_n 0.0125068f $X=3.495 $Y=1.225 $X2=0 $Y2=0
cc_294 N_TE_c_324_n N_A_27_74#_c_638_n 4.49351e-19 $X=4.065 $Y=1.225 $X2=0 $Y2=0
cc_295 N_TE_c_327_n N_A_27_74#_c_638_n 0.00227103f $X=3.065 $Y=1.3 $X2=0 $Y2=0
cc_296 N_TE_c_328_n N_A_27_74#_c_638_n 0.00227103f $X=3.495 $Y=1.3 $X2=0 $Y2=0
cc_297 N_TE_c_323_n N_A_27_74#_c_639_n 0.0118714f $X=3.99 $Y=1.3 $X2=0 $Y2=0
cc_298 N_TE_c_325_n N_A_27_74#_c_639_n 0.00473545f $X=4.98 $Y=1.3 $X2=0 $Y2=0
cc_299 N_TE_c_328_n N_A_27_74#_c_639_n 0.00696323f $X=3.495 $Y=1.3 $X2=0 $Y2=0
cc_300 N_TE_c_329_n N_A_27_74#_c_639_n 0.00726444f $X=4.065 $Y=1.3 $X2=0 $Y2=0
cc_301 N_TE_c_322_n N_A_27_74#_c_640_n 4.49351e-19 $X=3.495 $Y=1.225 $X2=0 $Y2=0
cc_302 N_TE_c_324_n N_A_27_74#_c_640_n 0.0140897f $X=4.065 $Y=1.225 $X2=0 $Y2=0
cc_303 N_TE_c_325_n N_A_27_74#_c_640_n 0.00830924f $X=4.98 $Y=1.3 $X2=0 $Y2=0
cc_304 N_TE_c_326_n N_A_27_74#_c_640_n 0.00123989f $X=5.055 $Y=1.225 $X2=0 $Y2=0
cc_305 N_TE_c_329_n N_A_27_74#_c_640_n 0.00227103f $X=4.065 $Y=1.3 $X2=0 $Y2=0
cc_306 N_TE_c_321_n N_A_27_74#_c_642_n 0.00334949f $X=3.42 $Y=1.3 $X2=0 $Y2=0
cc_307 N_TE_c_327_n N_A_27_74#_c_642_n 3.01213e-19 $X=3.065 $Y=1.3 $X2=0 $Y2=0
cc_308 N_TE_c_328_n N_A_27_74#_c_642_n 3.01213e-19 $X=3.495 $Y=1.3 $X2=0 $Y2=0
cc_309 N_TE_c_317_n N_VGND_c_727_n 0.00616282f $X=2.495 $Y=1.225 $X2=0 $Y2=0
cc_310 N_TE_c_318_n N_VGND_c_727_n 0.00525645f $X=2.99 $Y=1.3 $X2=0 $Y2=0
cc_311 N_TE_c_320_n N_VGND_c_727_n 0.00666821f $X=3.065 $Y=1.225 $X2=0 $Y2=0
cc_312 N_TE_c_322_n N_VGND_c_728_n 0.00666821f $X=3.495 $Y=1.225 $X2=0 $Y2=0
cc_313 N_TE_c_323_n N_VGND_c_728_n 0.00525645f $X=3.99 $Y=1.3 $X2=0 $Y2=0
cc_314 N_TE_c_324_n N_VGND_c_728_n 0.00805013f $X=4.065 $Y=1.225 $X2=0 $Y2=0
cc_315 N_TE_c_326_n N_VGND_c_730_n 0.0174858f $X=5.055 $Y=1.225 $X2=0 $Y2=0
cc_316 TE N_VGND_c_730_n 0.00881431f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_317 N_TE_c_331_n N_VGND_c_730_n 0.00676362f $X=5.255 $Y=1.495 $X2=0 $Y2=0
cc_318 N_TE_c_332_n N_VGND_c_730_n 0.0121897f $X=5.485 $Y=1.465 $X2=0 $Y2=0
cc_319 N_TE_c_320_n N_VGND_c_731_n 0.00434272f $X=3.065 $Y=1.225 $X2=0 $Y2=0
cc_320 N_TE_c_322_n N_VGND_c_731_n 0.00434272f $X=3.495 $Y=1.225 $X2=0 $Y2=0
cc_321 N_TE_c_317_n N_VGND_c_733_n 0.00430908f $X=2.495 $Y=1.225 $X2=0 $Y2=0
cc_322 N_TE_c_324_n N_VGND_c_734_n 0.00434272f $X=4.065 $Y=1.225 $X2=0 $Y2=0
cc_323 N_TE_c_326_n N_VGND_c_734_n 0.00434272f $X=5.055 $Y=1.225 $X2=0 $Y2=0
cc_324 N_TE_c_317_n N_VGND_c_736_n 0.00817403f $X=2.495 $Y=1.225 $X2=0 $Y2=0
cc_325 N_TE_c_320_n N_VGND_c_736_n 0.00821294f $X=3.065 $Y=1.225 $X2=0 $Y2=0
cc_326 N_TE_c_322_n N_VGND_c_736_n 0.00821294f $X=3.495 $Y=1.225 $X2=0 $Y2=0
cc_327 N_TE_c_324_n N_VGND_c_736_n 0.00826293f $X=4.065 $Y=1.225 $X2=0 $Y2=0
cc_328 N_TE_c_326_n N_VGND_c_736_n 0.0082925f $X=5.055 $Y=1.225 $X2=0 $Y2=0
cc_329 N_A_27_368#_c_419_n N_Z_M1000_s 0.00245557f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_330 N_A_27_368#_c_421_n N_Z_M1009_s 0.00197722f $X=2.065 $Y=2.99 $X2=0 $Y2=0
cc_331 N_A_27_368#_M1008_d N_Z_c_523_n 0.00480741f $X=1.08 $Y=1.84 $X2=0 $Y2=0
cc_332 N_A_27_368#_c_477_p N_Z_c_523_n 0.0184684f $X=1.28 $Y=2.455 $X2=0 $Y2=0
cc_333 N_A_27_368#_c_422_n N_Z_c_510_n 0.00625091f $X=2.23 $Y=1.985 $X2=0 $Y2=0
cc_334 N_A_27_368#_c_417_n N_Z_c_510_n 0.0141015f $X=2.395 $Y=1.725 $X2=0 $Y2=0
cc_335 N_A_27_368#_c_419_n N_Z_c_537_n 0.0185424f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_336 N_A_27_368#_c_477_p Z 0.0298377f $X=1.28 $Y=2.455 $X2=0 $Y2=0
cc_337 N_A_27_368#_c_421_n Z 0.0160777f $X=2.065 $Y=2.99 $X2=0 $Y2=0
cc_338 N_A_27_368#_c_421_n N_VPWR_c_570_n 0.0117278f $X=2.065 $Y=2.99 $X2=0
+ $Y2=0
cc_339 N_A_27_368#_c_423_n N_VPWR_c_570_n 0.0195643f $X=3.015 $Y=1.725 $X2=0
+ $Y2=0
cc_340 N_A_27_368#_c_425_n N_VPWR_c_570_n 0.0657084f $X=3.18 $Y=1.985 $X2=0
+ $Y2=0
cc_341 N_A_27_368#_c_425_n N_VPWR_c_571_n 0.0658989f $X=3.18 $Y=1.985 $X2=0
+ $Y2=0
cc_342 N_A_27_368#_c_426_n N_VPWR_c_571_n 0.0186422f $X=3.925 $Y=1.725 $X2=0
+ $Y2=0
cc_343 N_A_27_368#_c_427_n N_VPWR_c_571_n 0.0659091f $X=4.09 $Y=1.985 $X2=0
+ $Y2=0
cc_344 N_A_27_368#_c_419_n N_VPWR_c_574_n 0.0422607f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_345 N_A_27_368#_c_420_n N_VPWR_c_574_n 0.0236215f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_346 N_A_27_368#_c_421_n N_VPWR_c_574_n 0.0677651f $X=2.065 $Y=2.99 $X2=0
+ $Y2=0
cc_347 N_A_27_368#_c_428_n N_VPWR_c_574_n 0.0179217f $X=1.24 $Y=2.99 $X2=0 $Y2=0
cc_348 N_A_27_368#_c_425_n N_VPWR_c_575_n 0.0110241f $X=3.18 $Y=1.985 $X2=0
+ $Y2=0
cc_349 N_A_27_368#_c_427_n N_VPWR_c_576_n 0.0110241f $X=4.09 $Y=1.985 $X2=0
+ $Y2=0
cc_350 N_A_27_368#_c_419_n N_VPWR_c_569_n 0.0238634f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_351 N_A_27_368#_c_420_n N_VPWR_c_569_n 0.0127839f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_352 N_A_27_368#_c_421_n N_VPWR_c_569_n 0.0377062f $X=2.065 $Y=2.99 $X2=0
+ $Y2=0
cc_353 N_A_27_368#_c_425_n N_VPWR_c_569_n 0.00909194f $X=3.18 $Y=1.985 $X2=0
+ $Y2=0
cc_354 N_A_27_368#_c_427_n N_VPWR_c_569_n 0.00909194f $X=4.09 $Y=1.985 $X2=0
+ $Y2=0
cc_355 N_A_27_368#_c_428_n N_VPWR_c_569_n 0.00971942f $X=1.24 $Y=2.99 $X2=0
+ $Y2=0
cc_356 N_A_27_368#_c_423_n N_A_27_74#_c_636_n 0.0406282f $X=3.015 $Y=1.725 $X2=0
+ $Y2=0
cc_357 N_A_27_368#_c_467_n N_A_27_74#_c_636_n 0.00791142f $X=3.14 $Y=1.725 $X2=0
+ $Y2=0
cc_358 N_A_27_368#_c_423_n N_A_27_74#_c_637_n 0.00399999f $X=3.015 $Y=1.725
+ $X2=0 $Y2=0
cc_359 N_A_27_368#_c_417_n N_A_27_74#_c_637_n 0.0260989f $X=2.395 $Y=1.725 $X2=0
+ $Y2=0
cc_360 N_A_27_368#_c_426_n N_A_27_74#_c_639_n 0.0546439f $X=3.925 $Y=1.725 $X2=0
+ $Y2=0
cc_361 N_A_27_368#_c_426_n N_A_27_74#_c_642_n 0.0144544f $X=3.925 $Y=1.725 $X2=0
+ $Y2=0
cc_362 N_A_27_368#_c_467_n N_A_27_74#_c_642_n 0.0133727f $X=3.14 $Y=1.725 $X2=0
+ $Y2=0
cc_363 N_Z_c_508_n N_A_27_74#_M1005_d 0.00312259f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_364 N_Z_c_509_n N_A_27_74#_c_631_n 0.00540984f $X=0.945 $Y=1.095 $X2=0 $Y2=0
cc_365 N_Z_M1002_s N_A_27_74#_c_632_n 0.00289516f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_366 N_Z_c_513_n N_A_27_74#_c_632_n 0.0145454f $X=0.78 $Y=0.825 $X2=0 $Y2=0
cc_367 N_Z_c_508_n N_A_27_74#_c_632_n 0.00304353f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_368 N_Z_c_508_n N_A_27_74#_c_701_n 0.0178215f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_369 N_Z_M1014_s N_A_27_74#_c_634_n 0.00258847f $X=1.595 $Y=0.37 $X2=0 $Y2=0
cc_370 N_Z_c_508_n N_A_27_74#_c_634_n 0.00364245f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_371 N_Z_c_527_n N_A_27_74#_c_634_n 0.0133715f $X=1.78 $Y=0.825 $X2=0 $Y2=0
cc_372 N_Z_c_510_n N_A_27_74#_c_635_n 0.00816149f $X=1.755 $Y=1.95 $X2=0 $Y2=0
cc_373 N_Z_c_511_n N_A_27_74#_c_635_n 0.0100439f $X=1.78 $Y=1.095 $X2=0 $Y2=0
cc_374 N_Z_c_510_n N_A_27_74#_c_637_n 0.0118914f $X=1.755 $Y=1.95 $X2=0 $Y2=0
cc_375 N_A_27_74#_c_634_n N_VGND_c_727_n 0.011924f $X=2.115 $Y=0.34 $X2=0 $Y2=0
cc_376 N_A_27_74#_c_635_n N_VGND_c_727_n 0.0272062f $X=2.28 $Y=0.515 $X2=0 $Y2=0
cc_377 N_A_27_74#_c_636_n N_VGND_c_727_n 0.0264638f $X=3.115 $Y=1.385 $X2=0
+ $Y2=0
cc_378 N_A_27_74#_c_638_n N_VGND_c_727_n 0.0308484f $X=3.28 $Y=0.515 $X2=0 $Y2=0
cc_379 N_A_27_74#_c_638_n N_VGND_c_728_n 0.0308485f $X=3.28 $Y=0.515 $X2=0 $Y2=0
cc_380 N_A_27_74#_c_639_n N_VGND_c_728_n 0.0264638f $X=4.115 $Y=1.385 $X2=0
+ $Y2=0
cc_381 N_A_27_74#_c_640_n N_VGND_c_728_n 0.0308485f $X=4.28 $Y=0.515 $X2=0 $Y2=0
cc_382 N_A_27_74#_c_638_n N_VGND_c_731_n 0.0144922f $X=3.28 $Y=0.515 $X2=0 $Y2=0
cc_383 N_A_27_74#_c_632_n N_VGND_c_733_n 0.0423044f $X=1.115 $Y=0.34 $X2=0 $Y2=0
cc_384 N_A_27_74#_c_633_n N_VGND_c_733_n 0.0235688f $X=0.445 $Y=0.34 $X2=0 $Y2=0
cc_385 N_A_27_74#_c_634_n N_VGND_c_733_n 0.0658004f $X=2.115 $Y=0.34 $X2=0 $Y2=0
cc_386 N_A_27_74#_c_641_n N_VGND_c_733_n 0.023268f $X=1.28 $Y=0.34 $X2=0 $Y2=0
cc_387 N_A_27_74#_c_640_n N_VGND_c_734_n 0.0145639f $X=4.28 $Y=0.515 $X2=0 $Y2=0
cc_388 N_A_27_74#_c_632_n N_VGND_c_736_n 0.0239316f $X=1.115 $Y=0.34 $X2=0 $Y2=0
cc_389 N_A_27_74#_c_633_n N_VGND_c_736_n 0.0127152f $X=0.445 $Y=0.34 $X2=0 $Y2=0
cc_390 N_A_27_74#_c_634_n N_VGND_c_736_n 0.0365331f $X=2.115 $Y=0.34 $X2=0 $Y2=0
cc_391 N_A_27_74#_c_638_n N_VGND_c_736_n 0.0118826f $X=3.28 $Y=0.515 $X2=0 $Y2=0
cc_392 N_A_27_74#_c_640_n N_VGND_c_736_n 0.0119984f $X=4.28 $Y=0.515 $X2=0 $Y2=0
cc_393 N_A_27_74#_c_641_n N_VGND_c_736_n 0.0127566f $X=1.28 $Y=0.34 $X2=0 $Y2=0
