* File: sky130_fd_sc_ls__o31a_1.pex.spice
* Created: Wed Sep  2 11:21:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O31A_1%A_84_48# 1 2 9 11 13 15 16 17 20 24 28 31 36
+ 39 40
r74 33 36 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.59 $Y=1.485
+ $X2=0.71 $Y2=1.485
r75 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.485 $X2=0.59 $Y2=1.485
r76 31 40 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.17 $Y=1.95
+ $X2=3.17 $Y2=1.13
r77 26 40 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=3.085 $Y=0.96
+ $X2=3.085 $Y2=1.13
r78 26 28 11.6939 $w=3.38e-07 $l=3.45e-07 $layer=LI1_cond $X=3.085 $Y=0.96
+ $X2=3.085 $Y2=0.615
r79 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=2.035
+ $X2=2.36 $Y2=2.035
r80 24 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.085 $Y=2.035
+ $X2=3.17 $Y2=1.95
r81 24 25 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.085 $Y=2.035
+ $X2=2.525 $Y2=2.035
r82 20 22 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.36 $Y=2.375
+ $X2=2.36 $Y2=2.715
r83 18 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.12 $X2=2.36
+ $Y2=2.035
r84 18 20 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.36 $Y=2.12
+ $X2=2.36 $Y2=2.375
r85 16 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=2.035
+ $X2=2.36 $Y2=2.035
r86 16 17 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.195 $Y=2.035
+ $X2=0.795 $Y2=2.035
r87 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.71 $Y=1.95
+ $X2=0.795 $Y2=2.035
r88 14 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.71 $Y=1.65
+ $X2=0.71 $Y2=1.485
r89 14 15 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.71 $Y=1.65 $X2=0.71
+ $Y2=1.95
r90 11 34 57.4383 $w=2.94e-07 $l=3.13943e-07 $layer=POLY_cond $X=0.515 $Y=1.765
+ $X2=0.587 $Y2=1.485
r91 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.515 $Y=1.765
+ $X2=0.515 $Y2=2.4
r92 7 34 38.5845 $w=2.94e-07 $l=2.05925e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.587 $Y2=1.485
r93 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=0.74
r94 2 39 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.21
+ $Y=1.84 $X2=2.36 $Y2=2.035
r95 2 22 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=2.21
+ $Y=1.84 $X2=2.36 $Y2=2.715
r96 2 20 600 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=1 $X=2.21
+ $Y=1.84 $X2=2.36 $Y2=2.375
r97 1 28 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.87
+ $Y=0.47 $X2=3.08 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_1%A1 3 5 7 8 12
c33 5 0 1.19194e-19 $X=1.205 $Y=1.765
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.515 $X2=1.13 $Y2=1.515
r35 8 12 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=1.14 $Y=1.665
+ $X2=1.14 $Y2=1.515
r36 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.205 $Y=1.765
+ $X2=1.13 $Y2=1.515
r37 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.205 $Y=1.765
+ $X2=1.205 $Y2=2.34
r38 1 11 38.5562 $w=2.99e-07 $l=1.90526e-07 $layer=POLY_cond $X=1.075 $Y=1.35
+ $X2=1.13 $Y2=1.515
r39 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.075 $Y=1.35
+ $X2=1.075 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_1%A2 3 5 7 8 12
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.465 $X2=1.67 $Y2=1.465
r31 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.67 $Y=1.665 $X2=1.67
+ $Y2=1.465
r32 5 11 61.4066 $w=2.86e-07 $l=3.21714e-07 $layer=POLY_cond $X=1.625 $Y=1.765
+ $X2=1.67 $Y2=1.465
r33 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.625 $Y=1.765
+ $X2=1.625 $Y2=2.34
r34 1 11 38.6549 $w=2.86e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.58 $Y=1.3
+ $X2=1.67 $Y2=1.465
r35 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.58 $Y=1.3 $X2=1.58
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_1%A3 1 3 6 8 12
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.515 $X2=2.21 $Y2=1.515
r33 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.21 $Y=1.665
+ $X2=2.21 $Y2=1.515
r34 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.3 $Y=1.35
+ $X2=2.21 $Y2=1.515
r35 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.3 $Y=1.35 $X2=2.3
+ $Y2=0.79
r36 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.135 $Y=1.765
+ $X2=2.21 $Y2=1.515
r37 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.135 $Y=1.765
+ $X2=2.135 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_1%B1 1 3 6 8 12
r26 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.75
+ $Y=1.515 $X2=2.75 $Y2=1.515
r27 8 12 4.67207 $w=3.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.73 $Y=1.665
+ $X2=2.73 $Y2=1.515
r28 4 11 38.5562 $w=2.99e-07 $l=1.86145e-07 $layer=POLY_cond $X=2.795 $Y=1.35
+ $X2=2.75 $Y2=1.515
r29 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.795 $Y=1.35
+ $X2=2.795 $Y2=0.79
r30 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.675 $Y=1.765
+ $X2=2.75 $Y2=1.515
r31 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.675 $Y=1.765
+ $X2=2.675 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_1%X 1 2 9 13 14 15 16 23 32
c24 14 0 1.19194e-19 $X=0.155 $Y=1.95
r25 21 23 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=0.27 $Y=2.005
+ $X2=0.27 $Y2=2.035
r26 15 16 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=2.405
+ $X2=0.27 $Y2=2.775
r27 14 21 0.872119 $w=3.68e-07 $l=2.8e-08 $layer=LI1_cond $X=0.27 $Y=1.977
+ $X2=0.27 $Y2=2.005
r28 14 32 8.28963 $w=3.68e-07 $l=1.57e-07 $layer=LI1_cond $X=0.27 $Y=1.977
+ $X2=0.27 $Y2=1.82
r29 14 15 10.6835 $w=3.68e-07 $l=3.43e-07 $layer=LI1_cond $X=0.27 $Y=2.062
+ $X2=0.27 $Y2=2.405
r30 14 23 0.840972 $w=3.68e-07 $l=2.7e-08 $layer=LI1_cond $X=0.27 $Y=2.062
+ $X2=0.27 $Y2=2.035
r31 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.17 $Y=1.13 $X2=0.17
+ $Y2=1.82
r32 7 13 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=1.13
r33 7 9 13.9254 $w=3.58e-07 $l=4.35e-07 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=0.515
r34 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=1.985
r35 2 16 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=2.815
r36 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_1%VPWR 1 2 9 13 16 17 18 20 33 34 37
r37 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 31 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 25 37 10.8012 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=0.857 $Y2=3.33
r45 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.09 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 20 37 10.8012 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.857 $Y2=3.33
r49 20 22 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 18 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 18 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 16 30 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.735 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 16 17 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=2.735 $Y=3.33
+ $X2=2.892 $Y2=3.33
r54 15 33 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.05 $Y=3.33 $X2=3.12
+ $Y2=3.33
r55 15 17 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=3.05 $Y=3.33
+ $X2=2.892 $Y2=3.33
r56 11 17 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.892 $Y=3.245
+ $X2=2.892 $Y2=3.33
r57 11 13 28.9025 $w=3.13e-07 $l=7.9e-07 $layer=LI1_cond $X=2.892 $Y=3.245
+ $X2=2.892 $Y2=2.455
r58 7 37 1.88438 $w=4.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.857 $Y=3.245
+ $X2=0.857 $Y2=3.33
r59 7 9 21.478 $w=4.63e-07 $l=8.35e-07 $layer=LI1_cond $X=0.857 $Y=3.245
+ $X2=0.857 $Y2=2.41
r60 2 13 600 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=1 $X=2.75
+ $Y=1.84 $X2=2.9 $Y2=2.455
r61 1 9 300 $w=1.7e-07 $l=7.18227e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.84 $X2=0.925 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_1%VGND 1 2 9 15 18 19 20 22 35 36 39
r39 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r42 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r43 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r44 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r45 27 29 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.68
+ $Y2=0
r46 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r47 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r49 22 24 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r50 20 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r51 20 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r52 20 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r53 18 29 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.68
+ $Y2=0
r54 18 19 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.947
+ $Y2=0
r55 17 32 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.13 $Y=0 $X2=2.16
+ $Y2=0
r56 17 19 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=2.13 $Y=0 $X2=1.947
+ $Y2=0
r57 13 19 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.947 $Y=0.085
+ $X2=1.947 $Y2=0
r58 13 15 16.7341 $w=3.63e-07 $l=5.3e-07 $layer=LI1_cond $X=1.947 $Y=0.085
+ $X2=1.947 $Y2=0.615
r59 9 11 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.78 $Y=0.515
+ $X2=0.78 $Y2=0.965
r60 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r61 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0.515
r62 2 15 182 $w=1.7e-07 $l=3.55176e-07 $layer=licon1_NDIFF $count=1 $X=1.655
+ $Y=0.47 $X2=1.945 $Y2=0.615
r63 1 11 182 $w=1.7e-07 $l=6.9208e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.965
r64 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O31A_1%A_230_94# 1 2 9 11 12 15
r32 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.58 $Y=0.96
+ $X2=2.58 $Y2=0.615
r33 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.415 $Y=1.045
+ $X2=2.58 $Y2=0.96
r34 11 12 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=2.415 $Y=1.045
+ $X2=1.46 $Y2=1.045
r35 7 12 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=1.292 $Y=0.96
+ $X2=1.46 $Y2=1.045
r36 7 9 11.8684 $w=3.33e-07 $l=3.45e-07 $layer=LI1_cond $X=1.292 $Y=0.96
+ $X2=1.292 $Y2=0.615
r37 2 15 91 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=2 $X=2.375
+ $Y=0.47 $X2=2.58 $Y2=0.615
r38 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.15
+ $Y=0.47 $X2=1.29 $Y2=0.615
.ends

