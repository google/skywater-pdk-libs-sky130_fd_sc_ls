* File: sky130_fd_sc_ls__o211a_1.pex.spice
* Created: Fri Aug 28 13:43:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O211A_1%A_83_264# 1 2 3 12 14 16 18 21 22 23 24 27
+ 30 31 32 33 35 37 40 41 43 45
c110 43 0 1.43839e-19 $X=2.56 $Y=2.105
c111 22 0 1.605e-19 $X=1.01 $Y=1.97
c112 14 0 1.02493e-19 $X=0.505 $Y=1.765
r113 45 46 13.5953 $w=3.41e-07 $l=3.8e-07 $layer=LI1_cond $X=3.947 $Y=0.855
+ $X2=3.947 $Y2=1.235
r114 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.93
+ $Y=1.485 $X2=0.93 $Y2=1.485
r115 35 48 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=2.14 $X2=4.04
+ $Y2=2.055
r116 35 37 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.04 $Y=2.14
+ $X2=4.04 $Y2=2.815
r117 34 43 4.30018 $w=1.7e-07 $l=2.27376e-07 $layer=LI1_cond $X=2.835 $Y=2.055
+ $X2=2.615 $Y2=2.04
r118 33 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=2.055
+ $X2=4.04 $Y2=2.055
r119 33 34 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=3.875 $Y=2.055
+ $X2=2.835 $Y2=2.055
r120 31 46 4.81864 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=3.76 $Y=1.235
+ $X2=3.947 $Y2=1.235
r121 31 32 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=3.76 $Y=1.235
+ $X2=2.835 $Y2=1.235
r122 30 43 1.96316 $w=1.7e-07 $l=1.78115e-07 $layer=LI1_cond $X=2.75 $Y=1.94
+ $X2=2.615 $Y2=2.04
r123 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.75 $Y=1.32
+ $X2=2.835 $Y2=1.235
r124 29 30 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.75 $Y=1.32
+ $X2=2.75 $Y2=1.94
r125 25 43 1.96316 $w=3.3e-07 $l=1.24499e-07 $layer=LI1_cond $X=2.56 $Y=2.14
+ $X2=2.615 $Y2=2.04
r126 25 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.56 $Y=2.14
+ $X2=2.56 $Y2=2.815
r127 23 43 4.30018 $w=1.7e-07 $l=2.27376e-07 $layer=LI1_cond $X=2.395 $Y=2.055
+ $X2=2.615 $Y2=2.04
r128 23 24 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=2.395 $Y=2.055
+ $X2=1.095 $Y2=2.055
r129 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.01 $Y=1.97
+ $X2=1.095 $Y2=2.055
r130 21 40 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=1.65
+ $X2=1.01 $Y2=1.485
r131 21 22 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.01 $Y=1.65
+ $X2=1.01 $Y2=1.97
r132 17 41 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=0.595 $Y=1.485
+ $X2=0.93 $Y2=1.485
r133 17 18 5.03009 $w=3.3e-07 $l=1.15022e-07 $layer=POLY_cond $X=0.595 $Y=1.485
+ $X2=0.505 $Y2=1.542
r134 14 18 37.0704 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.542
r135 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r136 10 18 37.0704 $w=1.5e-07 $l=2.26945e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.505 $Y2=1.542
r137 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=0.74
r138 3 48 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.96 $X2=4.04 $Y2=2.135
r139 3 37 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.96 $X2=4.04 $Y2=2.815
r140 2 43 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=1.96 $X2=2.56 $Y2=2.105
r141 2 27 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=1.96 $X2=2.56 $Y2=2.815
r142 1 45 91 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_NDIFF $count=2 $X=3.785
+ $Y=0.68 $X2=3.97 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_1%A1 3 5 7 8 12 13
c38 5 0 1.43839e-19 $X=1.915 $Y=1.885
r39 12 14 10.2699 $w=3.52e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.677
+ $X2=1.915 $Y2=1.677
r40 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.84
+ $Y=1.635 $X2=1.84 $Y2=1.635
r41 10 12 20.5398 $w=3.52e-07 $l=1.5e-07 $layer=POLY_cond $X=1.69 $Y=1.677
+ $X2=1.84 $Y2=1.677
r42 8 13 0.535558 $w=6.68e-07 $l=3e-08 $layer=LI1_cond $X=1.67 $Y=1.665 $X2=1.67
+ $Y2=1.635
r43 5 14 22.7654 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.915 $Y=1.885
+ $X2=1.915 $Y2=1.677
r44 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.915 $Y=1.885
+ $X2=1.915 $Y2=2.46
r45 1 10 22.7654 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.69 $Y=1.47
+ $X2=1.69 $Y2=1.677
r46 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.69 $Y=1.47 $X2=1.69
+ $Y2=1
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_1%A2 1 2 3 5 9 11 12 13 20
r40 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.49
+ $Y=0.405 $X2=2.49 $Y2=0.405
r41 17 20 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=2.35 $Y=0.405
+ $X2=2.49 $Y2=0.405
r42 12 13 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=0.447
+ $X2=3.6 $Y2=0.447
r43 11 12 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=0.447
+ $X2=3.12 $Y2=0.447
r44 11 21 4.49004 $w=3.83e-07 $l=1.5e-07 $layer=LI1_cond $X=2.64 $Y=0.447
+ $X2=2.49 $Y2=0.447
r45 9 10 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.35 $Y=1 $X2=2.35
+ $Y2=1.41
r46 6 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=0.57
+ $X2=2.35 $Y2=0.405
r47 6 9 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.35 $Y=0.57 $X2=2.35
+ $Y2=1
r48 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.335 $Y=1.885
+ $X2=2.335 $Y2=2.46
r49 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.335 $Y=1.795 $X2=2.335
+ $Y2=1.885
r50 1 10 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.335 $Y=1.5 $X2=2.335
+ $Y2=1.41
r51 1 2 114.669 $w=1.8e-07 $l=2.95e-07 $layer=POLY_cond $X=2.335 $Y=1.5
+ $X2=2.335 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_1%B1 1 3 6 8 12
r36 12 14 8.87535 $w=3.53e-07 $l=6.5e-08 $layer=POLY_cond $X=3.17 $Y=1.677
+ $X2=3.235 $Y2=1.677
r37 10 12 52.5694 $w=3.53e-07 $l=3.85e-07 $layer=POLY_cond $X=2.785 $Y=1.677
+ $X2=3.17 $Y2=1.677
r38 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.635 $X2=3.17 $Y2=1.635
r39 4 14 22.8335 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.235 $Y=1.47
+ $X2=3.235 $Y2=1.677
r40 4 6 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.235 $Y=1.47 $X2=3.235
+ $Y2=1
r41 1 10 22.8335 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.785 $Y=1.885
+ $X2=2.785 $Y2=1.677
r42 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.785 $Y=1.885
+ $X2=2.785 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_1%C1 3 5 7 8
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.8
+ $Y=1.635 $X2=3.8 $Y2=1.635
r28 8 12 10.4092 $w=3.08e-07 $l=2.8e-07 $layer=LI1_cond $X=4.08 $Y=1.645 $X2=3.8
+ $Y2=1.645
r29 5 11 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=3.815 $Y=1.885
+ $X2=3.8 $Y2=1.635
r30 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.815 $Y=1.885
+ $X2=3.815 $Y2=2.46
r31 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.71 $Y=1.47
+ $X2=3.8 $Y2=1.635
r32 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.71 $Y=1.47 $X2=3.71
+ $Y2=1
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_1%X 1 2 9 13 14 15 16 23 32
c26 32 0 1.02493e-19 $X=0.265 $Y=1.82
r27 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=0.265 $Y=2 $X2=0.265
+ $Y2=2.035
r28 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.265 $Y=2.405
+ $X2=0.265 $Y2=2.775
r29 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.265 $Y=1.975
+ $X2=0.265 $Y2=2
r30 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=0.265 $Y=1.975
+ $X2=0.265 $Y2=1.82
r31 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=0.265 $Y=2.06
+ $X2=0.265 $Y2=2.405
r32 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.265 $Y=2.06
+ $X2=0.265 $Y2=2.035
r33 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.17 $Y=1.13 $X2=0.17
+ $Y2=1.82
r34 7 13 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=1.13
r35 7 9 13.9254 $w=3.58e-07 $l=4.35e-07 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=0.515
r36 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r37 2 16 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r38 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_1%VPWR 1 2 9 11 18 25 26 31 39 41
r42 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r43 38 39 13.4207 $w=1.103e-06 $l=1.65e-07 $layer=LI1_cond $X=1.69 $Y=2.862
+ $X2=1.855 $Y2=2.862
r44 35 38 0.110407 $w=1.103e-06 $l=1e-08 $layer=LI1_cond $X=1.68 $Y=2.862
+ $X2=1.69 $Y2=2.862
r45 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 33 35 9.93665 $w=1.103e-06 $l=9e-07 $layer=LI1_cond $X=0.78 $Y=2.862
+ $X2=1.68 $Y2=2.862
r47 30 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 29 33 0.662443 $w=1.103e-06 $l=6e-08 $layer=LI1_cond $X=0.72 $Y=2.862
+ $X2=0.78 $Y2=2.862
r49 29 31 12.7583 $w=1.103e-06 $l=1.05e-07 $layer=LI1_cond $X=0.72 $Y=2.862
+ $X2=0.615 $Y2=2.862
r50 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 26 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r53 23 41 14.7259 $w=1.7e-07 $l=4.05e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.3 $Y2=3.33
r54 23 25 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 22 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r56 21 39 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=1.855 $Y2=3.33
r57 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 18 41 14.7259 $w=1.7e-07 $l=4.05e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=3.3 $Y2=3.33
r59 18 21 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 16 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 15 31 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=0.615 $Y2=3.33
r62 15 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 11 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 11 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 7 41 3.15573 $w=8.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=3.245 $X2=3.3
+ $Y2=3.33
r66 7 9 12.5514 $w=8.08e-07 $l=8.5e-07 $layer=LI1_cond $X=3.3 $Y=3.245 $X2=3.3
+ $Y2=2.395
r67 2 9 150 $w=1.7e-07 $l=8.70747e-07 $layer=licon1_PDIFF $count=4 $X=2.86
+ $Y=1.96 $X2=3.54 $Y2=2.395
r68 1 38 200 $w=1.7e-07 $l=1.35947e-06 $layer=licon1_PDIFF $count=3 $X=0.58
+ $Y=1.84 $X2=1.69 $Y2=2.395
r69 1 33 200 $w=1.7e-07 $l=6.47321e-07 $layer=licon1_PDIFF $count=3 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r39 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r41 30 33 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r42 28 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r43 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r44 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r45 25 27 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.68
+ $Y2=0
r46 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r47 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r49 20 22 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r50 18 34 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r51 18 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r52 18 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r53 16 27 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.68
+ $Y2=0
r54 16 17 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.96
+ $Y2=0
r55 15 30 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.155 $Y=0 $X2=2.16
+ $Y2=0
r56 15 17 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.155 $Y=0 $X2=1.96
+ $Y2=0
r57 11 17 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0
r58 11 13 22.3101 $w=3.88e-07 $l=7.55e-07 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0.84
r59 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r60 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0.515
r61 2 13 182 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=1 $X=1.765
+ $Y=0.68 $X2=1.96 $Y2=0.84
r62 1 9 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O211A_1%A_257_136# 1 2 9 11 12 14 15 17
r38 15 17 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.495 $Y=0.895
+ $X2=3.02 $Y2=0.895
r39 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.41 $Y=0.98
+ $X2=2.495 $Y2=0.895
r40 13 14 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.41 $Y=0.98 $X2=2.41
+ $Y2=1.13
r41 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.325 $Y=1.215
+ $X2=2.41 $Y2=1.13
r42 11 12 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.325 $Y=1.215
+ $X2=1.595 $Y2=1.215
r43 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.43 $Y=1.13
+ $X2=1.595 $Y2=1.215
r44 7 9 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.43 $Y=1.13 $X2=1.43
+ $Y2=0.825
r45 2 17 91 $w=1.7e-07 $l=6.94226e-07 $layer=licon1_NDIFF $count=2 $X=2.425
+ $Y=0.68 $X2=3.02 $Y2=0.895
r46 1 9 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=1.285
+ $Y=0.68 $X2=1.475 $Y2=0.825
.ends

