* File: sky130_fd_sc_ls__a221o_2.spice
* Created: Fri Aug 28 12:52:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a221o_2.pex.spice"
.subckt sky130_fd_sc_ls__a221o_2  VNB VPB A2 A1 B1 B2 C1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C1	C1
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1012 N_X_M1012_d N_A_89_260#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1012_d N_A_89_260#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.17575 PD=1.02 PS=1.215 NRD=0 NRS=15.396 M=1 R=4.93333
+ SA=75000.6 SB=75003 A=0.111 P=1.78 MULT=1
MM1002 A_337_74# N_A2_M1002_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74 AD=0.0777
+ AS=0.17575 PD=0.95 PS=1.215 NRD=8.1 NRS=16.212 M=1 R=4.93333 SA=75001.2
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1011 N_A_89_260#_M1011_d N_A1_M1011_g A_337_74# VNB NSHORT L=0.15 W=0.74
+ AD=0.3034 AS=0.0777 PD=1.56 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75001.6
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1004 A_603_74# N_B1_M1004_g N_A_89_260#_M1011_d VNB NSHORT L=0.15 W=0.74
+ AD=0.0777 AS=0.3034 PD=0.95 PS=1.56 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_B2_M1006_g A_603_74# VNB NSHORT L=0.15 W=0.74 AD=0.1443
+ AS=0.0777 PD=1.13 PS=0.95 NRD=3.24 NRS=8.1 M=1 R=4.93333 SA=75002.9 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1009 N_A_89_260#_M1009_d N_C1_M1009_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1961 AS=0.1443 PD=2.01 PS=1.13 NRD=0 NRS=14.592 M=1 R=4.93333 SA=75003.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_X_M1007_d N_A_89_260#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1008 N_X_M1007_d N_A_89_260#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.210264 PD=1.42 PS=1.56906 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1010 N_A_316_392#_M1010_d N_A2_M1010_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.187736 PD=1.3 PS=1.40094 NRD=1.9503 NRS=14.775 M=1 R=6.66667
+ SA=75001.2 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g N_A_316_392#_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_316_392#_M1000_d N_B1_M1000_g N_A_515_392#_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1003 N_A_515_392#_M1003_d N_B2_M1003_g N_A_316_392#_M1000_d VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.6 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_A_89_260#_M1005_d N_C1_M1005_g N_A_515_392#_M1003_d VPB PHIGHVT L=0.15
+ W=1 AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__a221o_2.pxi.spice"
*
.ends
*
*
