* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 VGND B1 a_154_392# VNB nshort w=640000u l=150000u
+  ad=1.23862e+12p pd=1.191e+07u as=5.376e+11p ps=5.52e+06u
M1001 VGND a_154_392# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1002 a_154_392# C1 a_69_392# VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=8.5e+11p ps=7.7e+06u
M1003 a_334_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=1.2e+12p pd=1.04e+07u as=1.947e+12p ps=1.641e+07u
M1004 a_154_392# A1 a_1081_39# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=6.927e+11p ps=6.48e+06u
M1005 a_1081_39# A1 a_154_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_334_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_154_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1008 a_69_392# C1 a_154_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_154_392# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_888_105# A3 VGND VNB nshort w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=0p ps=0u
M1011 a_1081_39# A2 a_888_105# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_69_392# B1 a_334_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A2 a_334_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A3 a_888_105# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND C1 a_154_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A1 a_334_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_154_392# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_154_392# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_334_392# B1 a_69_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_888_105# A2 a_1081_39# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_154_392# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_154_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_154_392# B1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_154_392# C1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_154_392# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_334_392# A3 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR A3 a_334_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
