* File: sky130_fd_sc_ls__and4b_1.spice
* Created: Wed Sep  2 10:55:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__and4b_1.pex.spice"
.subckt sky130_fd_sc_ls__and4b_1  VNB VPB A_N B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_N_M1010_g N_A_27_74#_M1010_s VNB NSHORT L=0.15 W=0.55
+ AD=0.14575 AS=0.15675 PD=1.63 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1002 A_353_124# N_A_27_74#_M1002_g N_A_226_424#_M1002_s VNB NSHORT L=0.15
+ W=0.64 AD=0.110562 AS=0.1824 PD=1.04 PS=1.85 NRD=22.068 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002 A=0.096 P=1.58 MULT=1
MM1001 A_448_139# N_B_M1001_g A_353_124# VNB NSHORT L=0.15 W=0.64 AD=0.0768
+ AS=0.110562 PD=0.88 PS=1.04 NRD=12.18 NRS=22.068 M=1 R=4.26667 SA=75000.6
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1011 A_526_139# N_C_M1011_g A_448_139# VNB NSHORT L=0.15 W=0.64 AD=0.1709
+ AS=0.0768 PD=1.275 PS=0.88 NRD=39.744 NRS=12.18 M=1 R=4.26667 SA=75001
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1000_d N_D_M1000_g A_526_139# VNB NSHORT L=0.15 W=0.64
+ AD=0.144093 AS=0.1709 PD=1.08522 PS=1.275 NRD=14.988 NRS=39.744 M=1 R=4.26667
+ SA=75001.5 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1003 N_X_M1003_d N_A_226_424#_M1003_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.166607 PD=2.05 PS=1.25478 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VPWR_M1007_d N_A_N_M1007_g N_A_27_74#_M1007_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.168 AS=0.2478 PD=1.24 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75003.5 A=0.126 P=1.98 MULT=1
MM1005 N_A_226_424#_M1005_d N_A_27_74#_M1005_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1596 AS=0.168 PD=1.22 PS=1.24 NRD=5.8509 NRS=14.0658 M=1 R=5.6
+ SA=75000.8 SB=75003 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_B_M1004_g N_A_226_424#_M1005_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.3864 AS=0.1596 PD=1.76 PS=1.22 NRD=2.3443 NRS=17.5724 M=1 R=5.6
+ SA=75001.3 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1006 N_A_226_424#_M1006_d N_C_M1006_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.147 AS=0.3864 PD=1.19 PS=1.76 NRD=14.0658 NRS=2.3443 M=1 R=5.6 SA=75002.4
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_D_M1009_g N_A_226_424#_M1006_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2154 AS=0.147 PD=1.39714 PS=1.19 NRD=30.4759 NRS=2.3443 M=1 R=5.6
+ SA=75002.9 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1008 N_X_M1008_d N_A_226_424#_M1008_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.2872 PD=2.83 PS=1.86286 NRD=1.7533 NRS=17.5724 M=1 R=7.46667
+ SA=75002.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.224 P=13.68
*
.include "sky130_fd_sc_ls__and4b_1.pxi.spice"
*
.ends
*
*
