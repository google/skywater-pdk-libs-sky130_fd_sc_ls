# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__and3b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505000 1.180000 0.835000 1.510000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.755000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.350000 3.560000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.138200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.570000 1.800000 6.595000 1.970000 ;
        RECT 4.570000 1.970000 4.900000 2.980000 ;
        RECT 4.965000 0.350000 5.215000 0.960000 ;
        RECT 4.965000 0.960000 6.105000 1.130000 ;
        RECT 5.570000 1.970000 5.900000 2.980000 ;
        RECT 5.925000 0.350000 6.105000 0.960000 ;
        RECT 5.935000 1.130000 6.105000 1.800000 ;
        RECT 6.365000 1.550000 6.595000 1.800000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 0.285000 1.680000 ;
      RECT 0.115000  1.680000 1.305000 1.850000 ;
      RECT 0.475000  1.850000 0.805000 2.860000 ;
      RECT 0.615000  0.085000 0.875000 1.010000 ;
      RECT 0.975000  2.020000 1.305000 3.245000 ;
      RECT 1.135000  1.320000 1.525000 1.650000 ;
      RECT 1.135000  1.650000 1.305000 1.680000 ;
      RECT 1.175000  0.255000 2.365000 0.425000 ;
      RECT 1.175000  0.425000 1.505000 1.150000 ;
      RECT 1.475000  1.820000 1.865000 1.950000 ;
      RECT 1.475000  1.950000 3.900000 2.120000 ;
      RECT 1.475000  2.120000 1.805000 2.860000 ;
      RECT 1.685000  0.595000 1.865000 1.150000 ;
      RECT 1.695000  1.150000 1.865000 1.820000 ;
      RECT 1.975000  2.290000 2.305000 3.245000 ;
      RECT 2.035000  0.425000 2.365000 0.470000 ;
      RECT 2.035000  0.470000 3.295000 0.720000 ;
      RECT 2.035000  0.720000 2.365000 1.150000 ;
      RECT 2.475000  2.120000 2.805000 2.860000 ;
      RECT 2.535000  0.890000 2.865000 1.010000 ;
      RECT 2.535000  1.010000 4.285000 1.180000 ;
      RECT 2.975000  2.290000 3.305000 3.245000 ;
      RECT 3.525000  0.085000 3.855000 0.840000 ;
      RECT 3.535000  2.120000 3.900000 2.860000 ;
      RECT 3.730000  1.460000 5.765000 1.630000 ;
      RECT 3.730000  1.630000 3.900000 1.950000 ;
      RECT 4.035000  0.450000 4.285000 1.010000 ;
      RECT 4.070000  1.820000 4.400000 3.245000 ;
      RECT 4.465000  0.085000 4.795000 1.130000 ;
      RECT 4.755000  1.300000 5.765000 1.460000 ;
      RECT 5.070000  2.140000 5.400000 3.245000 ;
      RECT 5.395000  0.085000 5.725000 0.790000 ;
      RECT 6.070000  2.140000 6.400000 3.245000 ;
      RECT 6.275000  0.085000 6.605000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_ls__and3b_4
