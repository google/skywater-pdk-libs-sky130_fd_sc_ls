* NGSPICE file created from sky130_fd_sc_ls__a32o_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_244_368# B2 a_84_48# VPB phighvt w=1e+06u l=150000u
+  ad=8.95e+11p pd=7.79e+06u as=4e+11p ps=2.8e+06u
M1001 a_244_368# A3 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=1.1114e+12p ps=6.38e+06u
M1002 VPWR A2 a_244_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_84_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1004 a_601_94# B1 a_84_48# VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=4.032e+11p ps=2.54e+06u
M1005 a_259_94# A3 VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=6.004e+11p ps=4.48e+06u
M1006 a_337_94# A2 a_259_94# VNB nshort w=640000u l=150000u
+  ad=2.496e+11p pd=2.06e+06u as=0p ps=0u
M1007 a_244_368# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B2 a_601_94# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_84_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1010 a_84_48# B1 a_244_368# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_84_48# A1 a_337_94# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

