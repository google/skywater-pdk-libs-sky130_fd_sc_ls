* NGSPICE file created from sky130_fd_sc_ls__nand3_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nand3_2 A B C VGND VNB VPB VPWR Y
M1000 a_283_74# A Y VNB nshort w=740000u l=150000u
+  ad=7.123e+11p pd=5.5e+06u as=2.072e+11p ps=2.04e+06u
M1001 Y A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=1.0136e+12p pd=8.53e+06u as=1.4392e+12p ps=1.153e+07u
M1002 a_283_74# B a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=6.068e+11p ps=6.08e+06u
M1003 VPWR B Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_74# B a_283_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y C VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR C Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND C a_27_74# VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1008 Y B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A a_283_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_74# C VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

