* File: sky130_fd_sc_ls__decaphe_18.spice
* Created: Fri Aug 28 13:11:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__decaphe_18.pex.spice"
.subckt sky130_fd_sc_ls__decaphe_18  VNB VPB VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_s N_VPWR_M1000_g N_VGND_M1000_s VNB NSHORT L=7.85 W=0.775
+ AD=0.2015 AS=0.2015 PD=2.07 PS=2.07 NRD=0 NRS=0 M=1 R=0.0987261 SA=3.925e+06
+ SB=3.925e+06 A=6.08375 P=17.25 MULT=1
MM1001 N_VPWR_M1001_s N_VGND_M1001_g N_VPWR_M1001_s VPB PSHORT L=7.85 W=1.255
+ AD=0.3263 AS=0.3263 PD=3.03 PS=3.03 NRD=0 NRS=0 M=1 R=0.159873 SA=3.925e+06
+ SB=3.925e+06 A=9.85175 P=18.21 MULT=1
DX2_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_ls__decaphe_18.pxi.spice"
*
.ends
*
*
