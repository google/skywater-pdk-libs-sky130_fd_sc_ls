* File: sky130_fd_sc_ls__nor4bb_2.spice
* Created: Wed Sep  2 11:16:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nor4bb_2.pex.spice"
.subckt sky130_fd_sc_ls__nor4bb_2  VNB VPB C_N D_N B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* D_N	D_N
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_C_N_M1016_g N_A_27_392#_M1016_s VNB NSHORT L=0.15 W=0.64
+ AD=0.180725 AS=0.1824 PD=1.42 PS=1.85 NRD=15.936 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1004 N_A_311_124#_M1004_d N_D_N_M1004_g N_VGND_M1016_d VNB NSHORT L=0.15
+ W=0.64 AD=0.2496 AS=0.180725 PD=2.06 PS=1.42 NRD=17.808 NRS=42.624 M=1
+ R=4.26667 SA=75000.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1000 N_Y_M1000_d N_A_311_124#_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.4735 PD=1.02 PS=2.86 NRD=0 NRS=29.184 M=1 R=4.93333 SA=75000.5
+ SB=75004.1 A=0.111 P=1.78 MULT=1
MM1010 N_Y_M1000_d N_A_311_124#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2096 PD=1.02 PS=1.405 NRD=0 NRS=37.008 M=1 R=4.93333 SA=75000.9
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1010_s N_A_27_392#_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2096 AS=0.1036 PD=1.405 PS=1.02 NRD=37.008 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A_27_392#_M1011_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1011_d N_B_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.74 AD=0.1295
+ AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5 SB=75002.1
+ A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1019_d N_B_M1019_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.30155 AS=0.1036 PD=1.555 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.9
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VGND_M1019_d VNB NSHORT L=0.15 W=0.74
+ AD=0.12025 AS=0.30155 PD=1.065 PS=1.555 NRD=7.296 NRS=0 M=1 R=4.93333
+ SA=75003.9 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1017 N_Y_M1006_d N_A_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.74
+ AD=0.12025 AS=0.2109 PD=1.065 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.3
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_VPWR_M1014_d N_C_N_M1014_g N_A_27_392#_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.585 AS=0.295 PD=2.17 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1012 N_A_311_124#_M1012_d N_D_N_M1012_g N_VPWR_M1014_d VPB PHIGHVT L=0.15 W=1
+ AD=0.295 AS=0.585 PD=2.59 PS=2.17 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.5 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_A_493_368#_M1001_d N_A_311_124#_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1015 N_A_493_368#_M1015_d N_A_311_124#_M1015_g N_Y_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1005 N_A_772_368#_M1005_d N_A_27_392#_M1005_g N_A_493_368#_M1015_d VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=10.5395 NRS=1.7533 M=1
+ R=7.46667 SA=75001.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1008 N_A_772_368#_M1005_d N_A_27_392#_M1008_g N_A_493_368#_M1008_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.196 AS=0.3304 PD=1.47 PS=2.83 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75001.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1009 N_A_772_368#_M1009_d N_B_M1009_g N_A_985_368#_M1009_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1013 N_A_772_368#_M1009_d N_B_M1013_g N_A_985_368#_M1013_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1003 N_A_985_368#_M1013_s N_A_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1018 N_A_985_368#_M1018_d N_A_M1018_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=14.0988 P=18.88
*
.include "sky130_fd_sc_ls__nor4bb_2.pxi.spice"
*
.ends
*
*
