* File: sky130_fd_sc_ls__nor3b_4.spice
* Created: Wed Sep  2 11:15:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__nor3b_4.pex.spice"
.subckt sky130_fd_sc_ls__nor3b_4  VNB VPB B A C_N Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* C_N	C_N
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_B_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.74 AD=0.2442
+ AS=0.11285 PD=2.14 PS=1.045 NRD=7.296 NRS=4.044 M=1 R=4.93333 SA=75000.3
+ SB=75006.9 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_B_M1008_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.11285 PD=1.16 PS=1.045 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75006.4 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1008_d N_B_M1022_g N_Y_M1022_s VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.3 SB=75005.8
+ A=0.111 P=1.78 MULT=1
MM1025 N_VGND_M1025_d N_B_M1025_g N_Y_M1022_s VNB NSHORT L=0.15 W=0.74 AD=0.1295
+ AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.7 SB=75005.4
+ A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_A_468_264#_M1001_g N_VGND_M1025_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75004.9 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1001_d N_A_468_264#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75004.5 A=0.111 P=1.78 MULT=1
MM1011 N_Y_M1011_d N_A_468_264#_M1011_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.1
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1026 N_Y_M1011_d N_A_468_264#_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.6
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75004.1 SB=75003
+ A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1003_d N_A_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.2035 PD=1.02 PS=1.29 NRD=0 NRS=21.888 M=1 R=4.93333 SA=75004.6 SB=75002.5
+ A=0.111 P=1.78 MULT=1
MM1012 N_Y_M1012_d N_A_M1012_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74 AD=0.1295
+ AS=0.2035 PD=1.09 PS=1.29 NRD=0 NRS=21.888 M=1 R=4.93333 SA=75005.3 SB=75001.8
+ A=0.111 P=1.78 MULT=1
MM1020 N_Y_M1012_d N_A_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.74 AD=0.1295
+ AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75005.8 SB=75001.3
+ A=0.111 P=1.78 MULT=1
MM1007 N_A_468_264#_M1007_d N_C_N_M1007_g N_VGND_M1020_s VNB NSHORT L=0.15
+ W=0.74 AD=0.6771 AS=0.1295 PD=3.31 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75006.3 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1010 N_A_27_368#_M1010_d N_B_M1010_g N_A_126_368#_M1010_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.3 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1014 N_A_27_368#_M1014_d N_B_M1014_g N_A_126_368#_M1010_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75003 A=0.168 P=2.54 MULT=1
MM1016 N_A_27_368#_M1014_d N_B_M1016_g N_A_126_368#_M1016_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.21 PD=1.42 PS=1.495 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75001.2 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1021 N_A_27_368#_M1021_d N_B_M1021_g N_A_126_368#_M1016_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.21 PD=1.42 PS=1.495 NRD=1.7533 NRS=13.1793 M=1 R=7.46667
+ SA=75001.7 SB=75002 A=0.168 P=2.54 MULT=1
MM1002 N_Y_M1002_d N_A_468_264#_M1002_g N_A_27_368#_M1021_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1005 N_Y_M1002_d N_A_468_264#_M1005_g N_A_27_368#_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1017 N_Y_M1017_d N_A_468_264#_M1017_g N_A_27_368#_M1005_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1023 N_Y_M1017_d N_A_468_264#_M1023_g N_A_27_368#_M1023_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_126_368#_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g N_A_126_368#_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1018 N_VPWR_M1015_d N_A_M1018_g N_A_126_368#_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1024 N_VPWR_M1024_d N_A_M1024_g N_A_126_368#_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.264 AS=0.168 PD=1.77714 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75001 A=0.168 P=2.54 MULT=1
MM1013 N_A_468_264#_M1013_d N_C_N_M1013_g N_VPWR_M1024_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.126 AS=0.198 PD=1.14 PS=1.33286 NRD=2.3443 NRS=22.261 M=1 R=5.6
+ SA=75002.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1019 N_A_468_264#_M1013_d N_C_N_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.126 AS=0.2478 PD=1.14 PS=2.27 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75002.6 SB=75000.2 A=0.126 P=1.98 MULT=1
DX27_noxref VNB VPB NWDIODE A=14.9916 P=19.84
*
.include "sky130_fd_sc_ls__nor3b_4.pxi.spice"
*
.ends
*
*
