* NGSPICE file created from sky130_fd_sc_ls__dlrtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 VPWR RESET_B a_817_48# VPB phighvt w=1e+06u l=150000u
+  ad=1.5813e+12p pd=1.156e+07u as=3.5e+11p ps=2.7e+06u
M1001 a_643_74# a_216_424# a_568_392# VPB phighvt w=1e+06u l=150000u
+  ad=3.328e+11p pd=2.77e+06u as=2.7e+11p ps=2.54e+06u
M1002 a_216_424# GATE VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=9.349e+11p ps=8.16e+06u
M1003 VGND RESET_B a_1045_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1004 a_568_392# a_27_424# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_817_48# a_759_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.121e+11p ps=1.85e+06u
M1006 a_769_74# a_216_424# a_643_74# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.907e+11p ps=2.24e+06u
M1007 VGND a_817_48# a_769_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_216_424# GATE VPWR VPB phighvt w=840000u l=150000u
+  ad=4.3935e+11p pd=2.87e+06u as=0p ps=0u
M1009 a_759_508# a_363_74# a_643_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_216_424# a_363_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=3.2225e+11p ps=2.64e+06u
M1011 VPWR D a_27_424# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1012 Q a_817_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1013 Q a_817_48# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1014 a_1045_74# a_643_74# a_817_48# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1015 VPWR a_216_424# a_363_74# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1016 VGND D a_27_424# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1017 a_565_74# a_27_424# VGND VNB nshort w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1018 a_643_74# a_363_74# a_565_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_817_48# a_643_74# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

