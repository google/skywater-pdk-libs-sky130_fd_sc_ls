* File: sky130_fd_sc_ls__or4_4.pex.spice
* Created: Fri Aug 28 13:59:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__OR4_4%A_83_264# 1 2 3 10 12 15 17 19 22 24 26 29 31
+ 33 36 38 44 45 46 49 51 55 57 59 62 65 66 67 73
c159 57 0 6.34286e-20 $X=6.465 $Y=1.11
c160 24 0 2.58165e-20 $X=1.405 $Y=1.765
r161 80 81 49.5771 $w=3.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.495 $Y=1.542
+ $X2=1.855 $Y2=1.542
r162 77 78 56.4629 $w=3.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.995 $Y=1.542
+ $X2=1.405 $Y2=1.542
r163 76 77 5.50857 $w=3.5e-07 $l=4e-08 $layer=POLY_cond $X=0.955 $Y=1.542
+ $X2=0.995 $Y2=1.542
r164 75 76 53.7086 $w=3.5e-07 $l=3.9e-07 $layer=POLY_cond $X=0.565 $Y=1.542
+ $X2=0.955 $Y2=1.542
r165 74 75 8.26286 $w=3.5e-07 $l=6e-08 $layer=POLY_cond $X=0.505 $Y=1.542
+ $X2=0.565 $Y2=1.542
r166 71 73 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=5.46 $Y=2.07
+ $X2=5.625 $Y2=2.07
r167 67 68 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=4.935 $Y=0.875
+ $X2=4.935 $Y2=1.11
r168 65 83 12.3943 $w=3.5e-07 $l=9e-08 $layer=POLY_cond $X=2.16 $Y=1.542
+ $X2=2.25 $Y2=1.542
r169 65 81 42.0029 $w=3.5e-07 $l=3.05e-07 $layer=POLY_cond $X=2.16 $Y=1.542
+ $X2=1.855 $Y2=1.542
r170 64 65 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=1.485 $X2=2.16 $Y2=1.485
r171 61 62 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=6.55 $Y=1.195
+ $X2=6.55 $Y2=1.95
r172 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.465 $Y=2.035
+ $X2=6.55 $Y2=1.95
r173 59 73 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=6.465 $Y=2.035
+ $X2=5.625 $Y2=2.035
r174 58 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.1 $Y=1.11
+ $X2=4.935 $Y2=1.11
r175 57 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.465 $Y=1.11
+ $X2=6.55 $Y2=1.195
r176 57 58 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=6.465 $Y=1.11
+ $X2=5.1 $Y2=1.11
r177 53 67 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.935 $Y=0.79
+ $X2=4.935 $Y2=0.875
r178 53 55 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.935 $Y=0.79
+ $X2=4.935 $Y2=0.515
r179 52 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=0.875
+ $X2=3.085 $Y2=0.875
r180 51 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.77 $Y=0.875
+ $X2=4.935 $Y2=0.875
r181 51 52 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=4.77 $Y=0.875
+ $X2=3.25 $Y2=0.875
r182 47 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=0.79
+ $X2=3.085 $Y2=0.875
r183 47 49 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.085 $Y=0.79
+ $X2=3.085 $Y2=0.515
r184 45 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.92 $Y=0.875
+ $X2=3.085 $Y2=0.875
r185 45 46 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.92 $Y=0.875
+ $X2=2.325 $Y2=0.875
r186 44 64 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=1.32
+ $X2=2.24 $Y2=1.485
r187 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.24 $Y=0.96
+ $X2=2.325 $Y2=0.875
r188 43 44 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.24 $Y=0.96
+ $X2=2.24 $Y2=1.32
r189 41 80 2.06571 $w=3.5e-07 $l=1.5e-08 $layer=POLY_cond $X=1.48 $Y=1.542
+ $X2=1.495 $Y2=1.542
r190 41 78 10.3286 $w=3.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.48 $Y=1.542
+ $X2=1.405 $Y2=1.542
r191 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.48
+ $Y=1.485 $X2=1.48 $Y2=1.485
r192 38 64 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=1.485
+ $X2=2.24 $Y2=1.485
r193 38 40 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.155 $Y=1.485
+ $X2=1.48 $Y2=1.485
r194 34 83 22.6286 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.25 $Y=1.32
+ $X2=2.25 $Y2=1.542
r195 34 36 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.25 $Y=1.32
+ $X2=2.25 $Y2=0.74
r196 31 81 22.6286 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.542
r197 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r198 27 80 22.6286 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.495 $Y=1.32
+ $X2=1.495 $Y2=1.542
r199 27 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.495 $Y=1.32
+ $X2=1.495 $Y2=0.74
r200 24 78 22.6286 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.542
r201 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r202 20 77 22.6286 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.995 $Y=1.32
+ $X2=0.995 $Y2=1.542
r203 20 22 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.995 $Y=1.32
+ $X2=0.995 $Y2=0.74
r204 17 76 22.6286 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.542
r205 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r206 13 75 22.6286 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.565 $Y=1.32
+ $X2=0.565 $Y2=1.542
r207 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.565 $Y=1.32
+ $X2=0.565 $Y2=0.74
r208 10 74 22.6286 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.542
r209 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r210 3 71 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.31
+ $Y=1.96 $X2=5.46 $Y2=2.105
r211 2 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.795
+ $Y=0.37 $X2=4.935 $Y2=0.515
r212 1 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.37 $X2=3.085 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_4%B 1 2 3 5 6 8 10 11 13 14 15 16 20 22 23
c87 16 0 1.3894e-19 $X=4.23 $Y=1.215
r88 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.78
+ $Y=1.385 $X2=2.78 $Y2=1.385
r89 23 28 10.3184 $w=4.02e-07 $l=3.4e-07 $layer=LI1_cond $X=3.12 $Y=1.34
+ $X2=2.78 $Y2=1.34
r90 22 28 4.24876 $w=4.02e-07 $l=1.4e-07 $layer=LI1_cond $X=2.64 $Y=1.34
+ $X2=2.78 $Y2=1.34
r91 20 31 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=1.385
+ $X2=4.23 $Y2=1.55
r92 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.23
+ $Y=1.385 $X2=4.23 $Y2=1.385
r93 16 19 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.23 $Y=1.215
+ $X2=4.23 $Y2=1.385
r94 15 23 7.646 $w=4.02e-07 $l=1.73205e-07 $layer=LI1_cond $X=3.235 $Y=1.215
+ $X2=3.12 $Y2=1.34
r95 14 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.065 $Y=1.215
+ $X2=4.23 $Y2=1.215
r96 14 15 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.065 $Y=1.215
+ $X2=3.235 $Y2=1.215
r97 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.235 $Y=1.885
+ $X2=4.235 $Y2=2.46
r98 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.235 $Y=1.795
+ $X2=4.235 $Y2=1.885
r99 10 31 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=4.235 $Y=1.795
+ $X2=4.235 $Y2=1.55
r100 6 27 38.5662 $w=2.97e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.87 $Y=1.22
+ $X2=2.785 $Y2=1.385
r101 6 8 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.87 $Y=1.22 $X2=2.87
+ $Y2=0.74
r102 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.865 $Y=1.885
+ $X2=2.865 $Y2=2.46
r103 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.865 $Y=1.795
+ $X2=2.865 $Y2=1.885
r104 1 27 48.8089 $w=2.97e-07 $l=2.92276e-07 $layer=POLY_cond $X=2.865 $Y=1.64
+ $X2=2.785 $Y2=1.385
r105 1 2 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=2.865 $Y=1.64
+ $X2=2.865 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_4%A 3 5 7 8 10 11 16
c48 5 0 1.55009e-19 $X=3.315 $Y=1.885
r49 16 18 24.8651 $w=3.78e-07 $l=1.95e-07 $layer=POLY_cond $X=3.57 $Y=1.677
+ $X2=3.765 $Y2=1.677
r50 14 16 32.5159 $w=3.78e-07 $l=2.55e-07 $layer=POLY_cond $X=3.315 $Y=1.677
+ $X2=3.57 $Y2=1.677
r51 13 14 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=3.3 $Y=1.677
+ $X2=3.315 $Y2=1.677
r52 11 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.635 $X2=3.57 $Y2=1.635
r53 8 18 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.765 $Y=1.885
+ $X2=3.765 $Y2=1.677
r54 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.765 $Y=1.885
+ $X2=3.765 $Y2=2.46
r55 5 14 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.885
+ $X2=3.315 $Y2=1.677
r56 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.885
+ $X2=3.315 $Y2=2.46
r57 1 13 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.3 $Y=1.47 $X2=3.3
+ $Y2=1.677
r58 1 3 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=3.3 $Y=1.47 $X2=3.3
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_4%C 3 5 7 8 10 11 12 13 22 23
c64 5 0 2.44757e-19 $X=4.735 $Y=1.885
c65 3 0 6.34286e-20 $X=4.72 $Y=0.74
r66 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.15
+ $Y=1.53 $X2=6.15 $Y2=1.53
r67 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.77
+ $Y=1.605 $X2=4.77 $Y2=1.605
r68 13 22 4.16546 $w=4.13e-07 $l=1.5e-07 $layer=LI1_cond $X=6 $Y=1.572 $X2=6.15
+ $Y2=1.572
r69 12 13 13.3295 $w=4.13e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.572 $X2=6
+ $Y2=1.572
r70 12 23 4.99855 $w=4.13e-07 $l=1.8e-07 $layer=LI1_cond $X=5.52 $Y=1.572
+ $X2=5.34 $Y2=1.572
r71 11 23 8.81928 $w=4.15e-07 $l=3e-07 $layer=LI1_cond $X=5.04 $Y=1.572 $X2=5.34
+ $Y2=1.572
r72 11 19 8.03415 $w=4.1e-07 $l=2.7e-07 $layer=LI1_cond $X=5.04 $Y=1.572
+ $X2=4.77 $Y2=1.572
r73 8 21 69.185 $w=2.99e-07 $l=3.62422e-07 $layer=POLY_cond $X=6.135 $Y=1.885
+ $X2=6.15 $Y2=1.53
r74 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.135 $Y=1.885
+ $X2=6.135 $Y2=2.46
r75 5 18 57.6553 $w=2.91e-07 $l=2.96985e-07 $layer=POLY_cond $X=4.735 $Y=1.885
+ $X2=4.77 $Y2=1.605
r76 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.735 $Y=1.885
+ $X2=4.735 $Y2=2.46
r77 1 18 38.6072 $w=2.91e-07 $l=1.88348e-07 $layer=POLY_cond $X=4.72 $Y=1.44
+ $X2=4.77 $Y2=1.605
r78 1 3 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=4.72 $Y=1.44 $X2=4.72
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_4%D 1 3 5 6 8 10 11 13 15 16 17 22 25 28 29
c60 28 0 7.13014e-20 $X=6.45 $Y=0.42
r61 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.45
+ $Y=0.42 $X2=6.45 $Y2=0.42
r62 25 29 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.45 $Y=0.555
+ $X2=6.45 $Y2=0.42
r63 24 28 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=6.45 $Y=0.775
+ $X2=6.45 $Y2=0.42
r64 21 22 2.99935 $w=3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.685 $Y=1.335 $X2=5.7
+ $Y2=1.335
r65 20 21 89.9803 $w=3e-07 $l=4.5e-07 $layer=POLY_cond $X=5.235 $Y=1.335
+ $X2=5.685 $Y2=1.335
r66 18 20 2.99935 $w=3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.22 $Y=1.335
+ $X2=5.235 $Y2=1.335
r67 16 24 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.285 $Y=0.85
+ $X2=6.45 $Y2=0.775
r68 16 17 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=6.285 $Y=0.85
+ $X2=5.775 $Y2=0.85
r69 15 22 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.7 $Y=1.185 $X2=5.7
+ $Y2=1.335
r70 14 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.7 $Y=0.925
+ $X2=5.775 $Y2=0.85
r71 14 15 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=5.7 $Y=0.925 $X2=5.7
+ $Y2=1.185
r72 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.685 $Y=1.885
+ $X2=5.685 $Y2=2.46
r73 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.685 $Y=1.795
+ $X2=5.685 $Y2=1.885
r74 9 21 14.7197 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.685 $Y=1.485
+ $X2=5.685 $Y2=1.335
r75 9 10 120.5 $w=1.8e-07 $l=3.1e-07 $layer=POLY_cond $X=5.685 $Y=1.485
+ $X2=5.685 $Y2=1.795
r76 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.235 $Y=1.885
+ $X2=5.235 $Y2=2.46
r77 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.235 $Y=1.795 $X2=5.235
+ $Y2=1.885
r78 4 20 14.7197 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.235 $Y=1.485
+ $X2=5.235 $Y2=1.335
r79 4 5 120.5 $w=1.8e-07 $l=3.1e-07 $layer=POLY_cond $X=5.235 $Y=1.485 $X2=5.235
+ $Y2=1.795
r80 1 18 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.22 $Y=1.185
+ $X2=5.22 $Y2=1.335
r81 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.22 $Y=1.185
+ $X2=5.22 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_4%VPWR 1 2 3 4 13 15 19 23 27 29 31 36 41 51 52
+ 58 61 64
r86 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r87 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r88 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r89 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r90 51 52 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r91 49 52 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6.48 $Y2=3.33
r92 49 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r93 48 51 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=6.48 $Y2=3.33
r94 48 49 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r95 46 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.54 $Y2=3.33
r96 46 48 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r97 45 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r98 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r99 42 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.08 $Y2=3.33
r100 42 44 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=3.12 $Y2=3.33
r101 41 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.54 $Y2=3.33
r102 41 44 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.12 $Y2=3.33
r103 40 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 40 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r105 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r106 37 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r107 37 39 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r108 36 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=2.08 $Y2=3.33
r109 36 39 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=1.68 $Y2=3.33
r110 35 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 35 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r112 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 32 55 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r114 32 34 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r115 31 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r116 31 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r117 29 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.6 $Y2=3.33
r118 29 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r119 25 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=3.245
+ $X2=3.54 $Y2=3.33
r120 25 27 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.54 $Y=3.245
+ $X2=3.54 $Y2=2.815
r121 21 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.08 $Y2=3.33
r122 21 23 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.08 $Y2=2.405
r123 17 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r124 17 19 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.405
r125 13 55 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r126 13 15 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.405
r127 4 27 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.39
+ $Y=1.96 $X2=3.54 $Y2=2.815
r128 3 23 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.405
r129 2 19 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.405
r130 1 15 300 $w=1.7e-07 $l=6.33364e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.405
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_4%X 1 2 3 4 15 17 19 21 25 29 31 33 34 35 42
c69 17 0 2.58165e-20 $X=0.73 $Y=2.15
r70 43 53 5.02295 $w=3.3e-07 $l=4.1e-07 $layer=LI1_cond $X=0.945 $Y=1.985
+ $X2=0.535 $Y2=1.985
r71 34 42 3.78902 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=1.63 $Y=1.985
+ $X2=1.515 $Y2=1.985
r72 34 46 3.78902 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=1.63 $Y=1.985
+ $X2=1.745 $Y2=1.985
r73 34 35 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.755 $Y=1.985
+ $X2=2.16 $Y2=1.985
r74 34 46 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=1.755 $Y=1.985
+ $X2=1.745 $Y2=1.985
r75 33 42 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.2 $Y=1.985
+ $X2=1.515 $Y2=1.985
r76 33 43 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.2 $Y=1.985
+ $X2=0.945 $Y2=1.985
r77 31 53 0.890511 $w=6.85e-07 $l=5e-08 $layer=LI1_cond $X=0.535 $Y=2.035
+ $X2=0.535 $Y2=1.985
r78 27 29 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.78 $Y=0.98
+ $X2=1.78 $Y2=0.515
r79 23 34 2.66947 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.63 $Y=2.15
+ $X2=1.63 $Y2=1.985
r80 23 25 11.775 $w=2.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.63 $Y=2.15
+ $X2=1.63 $Y2=2.385
r81 22 53 16.3854 $w=6.85e-07 $l=1.10616e-06 $layer=LI1_cond $X=0.945 $Y=1.065
+ $X2=0.535 $Y2=1.985
r82 21 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.615 $Y=1.065
+ $X2=1.78 $Y2=0.98
r83 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=1.065
+ $X2=0.945 $Y2=1.065
r84 17 31 7.81937 $w=6.85e-07 $l=2.45866e-07 $layer=LI1_cond $X=0.73 $Y=2.15
+ $X2=0.535 $Y2=2.035
r85 17 19 11.775 $w=2.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.73 $Y=2.15
+ $X2=0.73 $Y2=2.385
r86 13 22 4.8017 $w=6.85e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=0.98
+ $X2=0.945 $Y2=1.065
r87 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.78 $Y=0.98
+ $X2=0.78 $Y2=0.515
r88 4 34 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=1.985
r89 4 25 300 $w=1.7e-07 $l=6.15447e-07 $layer=licon1_PDIFF $count=2 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.385
r90 3 53 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r91 3 19 300 $w=1.7e-07 $l=6.15447e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.385
r92 2 29 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.57
+ $Y=0.37 $X2=1.78 $Y2=0.515
r93 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_4%A_499_392# 1 2 3 10 12 14 16 17 20 22 30 32
r69 23 30 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.675 $Y=2.445
+ $X2=4.51 $Y2=2.445
r70 22 32 4.85386 $w=1.7e-07 $l=1.81659e-07 $layer=LI1_cond $X=6.245 $Y=2.445
+ $X2=6.41 $Y2=2.41
r71 22 23 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=6.245 $Y=2.445
+ $X2=4.675 $Y2=2.445
r72 18 30 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.51 $Y=2.53 $X2=4.51
+ $Y2=2.445
r73 18 20 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=4.51 $Y=2.53
+ $X2=4.51 $Y2=2.815
r74 17 30 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.51 $Y=2.36 $X2=4.51
+ $Y2=2.445
r75 16 29 2.77363 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=4.51 $Y=2.14 $X2=4.51
+ $Y2=2.04
r76 16 17 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=4.51 $Y=2.14
+ $X2=4.51 $Y2=2.36
r77 15 27 3.96311 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=2.805 $Y=2.055
+ $X2=2.64 $Y2=2.065
r78 14 29 4.99254 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.345 $Y=2.055
+ $X2=4.51 $Y2=2.04
r79 14 15 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=4.345 $Y=2.055
+ $X2=2.805 $Y2=2.055
r80 10 27 3.39695 $w=2.8e-07 $l=1.36931e-07 $layer=LI1_cond $X=2.615 $Y=2.19
+ $X2=2.64 $Y2=2.065
r81 10 12 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=2.615 $Y=2.19
+ $X2=2.615 $Y2=2.445
r82 3 32 300 $w=1.7e-07 $l=5.86536e-07 $layer=licon1_PDIFF $count=2 $X=6.21
+ $Y=1.96 $X2=6.41 $Y2=2.455
r83 2 29 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=4.31
+ $Y=1.96 $X2=4.51 $Y2=2.105
r84 2 20 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=4.31
+ $Y=1.96 $X2=4.51 $Y2=2.815
r85 1 27 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.96 $X2=2.64 $Y2=2.105
r86 1 12 300 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=1.96 $X2=2.64 $Y2=2.445
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_4%A_588_392# 1 2 7 9 11 13 15
c28 15 0 1.05817e-19 $X=4 $Y=2.815
c29 9 0 1.55009e-19 $X=3.09 $Y=2.815
r30 13 20 3.14031 $w=2.8e-07 $l=1.41421e-07 $layer=LI1_cond $X=4.035 $Y=2.56
+ $X2=4 $Y2=2.435
r31 13 15 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=4.035 $Y=2.56
+ $X2=4.035 $Y2=2.815
r32 12 18 4.12165 $w=2e-07 $l=1.4e-07 $layer=LI1_cond $X=3.205 $Y=2.46 $X2=3.065
+ $Y2=2.46
r33 11 20 3.92538 $w=2e-07 $l=1.87083e-07 $layer=LI1_cond $X=3.825 $Y=2.46 $X2=4
+ $Y2=2.435
r34 11 12 34.3818 $w=1.98e-07 $l=6.2e-07 $layer=LI1_cond $X=3.825 $Y=2.46
+ $X2=3.205 $Y2=2.46
r35 7 18 2.94404 $w=2.8e-07 $l=1e-07 $layer=LI1_cond $X=3.065 $Y=2.56 $X2=3.065
+ $Y2=2.46
r36 7 9 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=3.065 $Y=2.56
+ $X2=3.065 $Y2=2.815
r37 2 20 600 $w=1.7e-07 $l=5.08748e-07 $layer=licon1_PDIFF $count=1 $X=3.84
+ $Y=1.96 $X2=4 $Y2=2.395
r38 2 15 600 $w=1.7e-07 $l=9.31571e-07 $layer=licon1_PDIFF $count=1 $X=3.84
+ $Y=1.96 $X2=4 $Y2=2.815
r39 1 18 600 $w=1.7e-07 $l=5.70088e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.96 $X2=3.09 $Y2=2.46
r40 1 9 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.96 $X2=3.09 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_4%A_962_392# 1 2 11
r14 8 11 37.0428 $w=2.78e-07 $l=9e-07 $layer=LI1_cond $X=5.01 $Y=2.84 $X2=5.91
+ $Y2=2.84
r15 2 11 600 $w=1.7e-07 $l=9.11921e-07 $layer=licon1_PDIFF $count=1 $X=5.76
+ $Y=1.96 $X2=5.91 $Y2=2.8
r16 1 8 600 $w=1.7e-07 $l=9.34666e-07 $layer=licon1_PDIFF $count=1 $X=4.81
+ $Y=1.96 $X2=5.01 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_LS__OR4_4%VGND 1 2 3 4 5 16 18 22 26 28 30 35 52 53 59
+ 62 66 75 78 84
c77 53 0 7.13014e-20 $X=6.48 $Y=0
r78 82 84 10.4353 $w=7.63e-07 $l=1.15e-07 $layer=LI1_cond $X=6 $Y=0.297
+ $X2=6.115 $Y2=0.297
r79 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r80 80 82 0.781751 $w=7.63e-07 $l=5e-08 $layer=LI1_cond $X=5.95 $Y=0.297 $X2=6
+ $Y2=0.297
r81 77 80 8.05203 $w=7.63e-07 $l=5.15e-07 $layer=LI1_cond $X=5.435 $Y=0.297
+ $X2=5.95 $Y2=0.297
r82 77 78 11.2171 $w=7.63e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=0.297
+ $X2=5.27 $Y2=0.297
r83 74 75 10.8372 $w=7.03e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=0.267
+ $X2=4.59 $Y2=0.267
r84 71 74 5.85315 $w=7.03e-07 $l=3.45e-07 $layer=LI1_cond $X=4.08 $Y=0.267
+ $X2=4.425 $Y2=0.267
r85 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r86 69 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r87 68 71 8.14351 $w=7.03e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=0.267
+ $X2=4.08 $Y2=0.267
r88 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r89 65 68 0.0848283 $w=7.03e-07 $l=5e-09 $layer=LI1_cond $X=3.595 $Y=0.267
+ $X2=3.6 $Y2=0.267
r90 65 66 10.8372 $w=7.03e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=0.267
+ $X2=3.43 $Y2=0.267
r91 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r92 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r93 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r94 53 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r95 52 84 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=6.115
+ $Y2=0
r96 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r97 49 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r98 49 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.08
+ $Y2=0
r99 48 78 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=5.27
+ $Y2=0
r100 48 75 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=4.59
+ $Y2=0
r101 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r102 44 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r103 43 66 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=3.43
+ $Y2=0
r104 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r105 41 62 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=2.56
+ $Y2=0
r106 41 43 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=3.12
+ $Y2=0
r107 39 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r108 39 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r109 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r110 36 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.28
+ $Y2=0
r111 36 38 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.445 $Y=0
+ $X2=2.16 $Y2=0
r112 35 62 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.38 $Y=0 $X2=2.56
+ $Y2=0
r113 35 38 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.38 $Y=0 $X2=2.16
+ $Y2=0
r114 34 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r115 34 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r116 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r117 31 56 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r118 31 33 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r119 30 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.28
+ $Y2=0
r120 30 33 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=0.72 $Y2=0
r121 28 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r122 28 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r123 24 62 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0
r124 24 26 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0.455
r125 20 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0
r126 20 22 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0.58
r127 16 56 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r128 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.515
r129 5 80 182 $w=1.7e-07 $l=7.23878e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.37 $X2=5.95 $Y2=0.515
r130 5 77 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.37 $X2=5.435 $Y2=0.515
r131 4 74 121.333 $w=1.7e-07 $l=1.09167e-06 $layer=licon1_NDIFF $count=1
+ $X=3.375 $Y=0.37 $X2=4.425 $Y2=0.455
r132 4 65 121.333 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1
+ $X=3.375 $Y=0.37 $X2=3.595 $Y2=0.455
r133 3 26 182 $w=1.7e-07 $l=2.74226e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.37 $X2=2.56 $Y2=0.455
r134 2 22 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.58
r135 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

