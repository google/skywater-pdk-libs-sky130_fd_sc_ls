* NGSPICE file created from sky130_fd_sc_ls__o21ba_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 X a_193_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=2.2288e+12p ps=1.517e+07u
M1001 VPWR a_27_368# a_193_48# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=5.52e+11p ps=4.88e+06u
M1002 VPWR A1 a_892_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=6e+11p ps=5.2e+06u
M1003 VGND a_193_48# X VNB nshort w=740000u l=150000u
+  ad=1.0914e+12p pd=1.012e+07u as=4.218e+11p ps=4.1e+06u
M1004 VGND A2 a_618_94# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=7.9445e+11p ps=7.84e+06u
M1005 VGND a_193_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_618_94# A1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_193_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_193_48# a_27_368# a_618_94# VNB nshort w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1009 a_618_94# A2 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1 a_618_94# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_193_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_193_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_892_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_618_94# a_27_368# a_193_48# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR B1_N a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1016 a_193_48# a_27_368# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_193_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND B1_N a_27_368# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1019 X a_193_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_193_48# A2 a_892_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_892_392# A2 a_193_48# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

