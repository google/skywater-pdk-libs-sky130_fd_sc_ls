* File: sky130_fd_sc_ls__dfxbp_1.spice
* Created: Fri Aug 28 13:16:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dfxbp_1.pex.spice"
.subckt sky130_fd_sc_ls__dfxbp_1  VNB VPB CLK D VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1023 N_VGND_M1023_d N_CLK_M1023_g N_A_27_74#_M1023_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2017 AS=0.2109 PD=1.35 PS=2.05 NRD=17.832 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1016 N_A_205_368#_M1016_d N_A_27_74#_M1016_g N_VGND_M1023_d VNB NSHORT L=0.15
+ W=0.74 AD=0.3252 AS=0.2017 PD=2.59 PS=1.35 NRD=62.34 NRS=4.452 M=1 R=4.93333
+ SA=75000.8 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1008 N_A_420_503#_M1008_d N_D_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.368725 PD=0.7 PS=2.64 NRD=0 NRS=235.116 M=1 R=2.8 SA=75000.6
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_543_447#_M1002_d N_A_27_74#_M1002_g N_A_420_503#_M1008_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0756875 AS=0.0588 PD=0.83 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1011 A_713_102# N_A_205_368#_M1011_g N_A_543_447#_M1002_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0756875 PD=0.63 PS=0.83 NRD=14.28 NRS=12.852 M=1 R=2.8
+ SA=75001.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_701_463#_M1003_g A_713_102# VNB NSHORT L=0.15 W=0.42
+ AD=0.125675 AS=0.0441 PD=1.03052 PS=0.63 NRD=69.768 NRS=14.28 M=1 R=2.8
+ SA=75001.6 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1006 N_A_701_463#_M1006_d N_A_543_447#_M1006_g N_VGND_M1003_d VNB NSHORT
+ L=0.15 W=0.55 AD=0.11825 AS=0.164575 PD=1.13 PS=1.34948 NRD=34.908 NRS=3.264
+ M=1 R=3.66667 SA=75001.7 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1010 N_A_1005_120#_M1010_d N_A_205_368#_M1010_g N_A_701_463#_M1006_d VNB
+ NSHORT L=0.15 W=0.55 AD=0.147026 AS=0.11825 PD=1.23608 PS=1.13 NRD=27.264
+ NRS=0 M=1 R=3.66667 SA=75001.8 SB=75001 A=0.0825 P=1.4 MULT=1
MM1019 A_1143_146# N_A_27_74#_M1019_g N_A_1005_120#_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.112274 PD=0.66 PS=0.943918 NRD=18.564 NRS=38.568 M=1
+ R=2.8 SA=75002.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_1191_120#_M1012_g A_1143_146# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_1005_120#_M1018_g N_A_1191_120#_M1018_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.11874 AS=0.15675 PD=0.989147 PS=1.67 NRD=15.264 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1004 N_Q_M1004_d N_A_1191_120#_M1004_g N_VGND_M1018_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.15976 PD=2.05 PS=1.33085 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1022_d N_A_1191_120#_M1022_g N_A_1644_112#_M1022_s VNB NSHORT
+ L=0.15 W=0.55 AD=0.107506 AS=0.15675 PD=0.937984 PS=1.67 NRD=18 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1026 N_Q_N_M1026_d N_A_1644_112#_M1026_g N_VGND_M1022_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.144644 PD=2.05 PS=1.26202 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_VPWR_M1020_d N_CLK_M1020_g N_A_27_74#_M1020_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3248 PD=1.42 PS=2.82 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1021 N_A_205_368#_M1021_d N_A_27_74#_M1021_g N_VPWR_M1020_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3192 AS=0.168 PD=2.81 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1015 N_A_420_503#_M1015_d N_D_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.146375 AS=0.2282 PD=1.335 PS=2.1 NRD=137.664 NRS=229.032 M=1 R=2.8
+ SA=75000.3 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1024 N_A_543_447#_M1024_d N_A_205_368#_M1024_g N_A_420_503#_M1015_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.107537 AS=0.146375 PD=1.11 PS=1.335 NRD=0
+ NRS=137.664 M=1 R=2.8 SA=75000.5 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1007 A_650_508# N_A_27_74#_M1007_g N_A_543_447#_M1024_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.107537 PD=0.69 PS=1.11 NRD=37.5088 NRS=94.2842 M=1 R=2.8
+ SA=75000.5 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_701_463#_M1001_g A_650_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.15505 AS=0.0567 PD=1.14333 PS=0.69 NRD=60.9715 NRS=37.5088 M=1 R=2.8
+ SA=75001 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1017 N_A_701_463#_M1017_d N_A_543_447#_M1017_g N_VPWR_M1001_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2541 AS=0.3101 PD=1.445 PS=2.28667 NRD=3.5066 NRS=73.678
+ M=1 R=5.6 SA=75001 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1025 N_A_1005_120#_M1025_d N_A_27_74#_M1025_g N_A_701_463#_M1017_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1878 AS=0.2541 PD=1.63333 PS=1.445 NRD=2.3443 NRS=56.2829
+ M=1 R=5.6 SA=75001.7 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1014 A_1158_482# N_A_205_368#_M1014_g N_A_1005_120#_M1025_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0939 PD=0.66 PS=0.816667 NRD=30.4759 NRS=44.5417 M=1
+ R=2.8 SA=75002.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1027 N_VPWR_M1027_d N_A_1191_120#_M1027_g A_1158_482# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.8
+ SA=75003.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_1005_120#_M1009_g N_A_1191_120#_M1009_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.182453 AS=0.29 PD=1.39151 PS=2.58 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1013 N_Q_M1013_d N_A_1191_120#_M1013_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3192 AS=0.204347 PD=2.81 PS=1.55849 NRD=1.7533 NRS=11.426 M=1
+ R=7.46667 SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_VPWR_M1000_d N_A_1191_120#_M1000_g N_A_1644_112#_M1000_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1596 AS=0.2394 PD=1.26429 PS=2.25 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1005 N_Q_N_M1005_d N_A_1644_112#_M1005_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3248 AS=0.2128 PD=2.82 PS=1.68571 NRD=1.7533 NRS=11.426 M=1
+ R=7.46667 SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX28_noxref VNB VPB NWDIODE A=18.5628 P=23.68
c_203 VPB 0 8.5492e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__dfxbp_1.pxi.spice"
*
.ends
*
*
