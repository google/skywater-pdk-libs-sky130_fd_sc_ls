* File: sky130_fd_sc_ls__sdfrtn_1.pxi.spice
* Created: Wed Sep  2 11:27:08 2020
* 
x_PM_SKY130_FD_SC_LS__SDFRTN_1%SCE N_SCE_M1037_g N_SCE_c_280_n N_SCE_c_289_n
+ N_SCE_M1030_g N_SCE_M1031_g N_SCE_M1003_g N_SCE_c_282_n N_SCE_c_283_n
+ N_SCE_c_284_n N_SCE_c_285_n SCE N_SCE_c_286_n N_SCE_c_287_n
+ PM_SKY130_FD_SC_LS__SDFRTN_1%SCE
x_PM_SKY130_FD_SC_LS__SDFRTN_1%A_27_88# N_A_27_88#_M1037_s N_A_27_88#_M1030_s
+ N_A_27_88#_M1019_g N_A_27_88#_c_355_n N_A_27_88#_c_356_n N_A_27_88#_M1035_g
+ N_A_27_88#_c_347_n N_A_27_88#_c_348_n N_A_27_88#_c_358_n N_A_27_88#_c_359_n
+ N_A_27_88#_c_360_n N_A_27_88#_c_349_n N_A_27_88#_c_350_n N_A_27_88#_c_362_n
+ N_A_27_88#_c_351_n N_A_27_88#_c_352_n N_A_27_88#_c_353_n N_A_27_88#_c_354_n
+ PM_SKY130_FD_SC_LS__SDFRTN_1%A_27_88#
x_PM_SKY130_FD_SC_LS__SDFRTN_1%D N_D_c_440_n N_D_M1002_g N_D_c_441_n N_D_M1022_g
+ N_D_c_443_n D D N_D_c_444_n N_D_c_445_n PM_SKY130_FD_SC_LS__SDFRTN_1%D
x_PM_SKY130_FD_SC_LS__SDFRTN_1%SCD N_SCD_c_482_n N_SCD_M1016_g N_SCD_c_483_n
+ N_SCD_M1034_g N_SCD_c_484_n SCD SCD N_SCD_c_481_n
+ PM_SKY130_FD_SC_LS__SDFRTN_1%SCD
x_PM_SKY130_FD_SC_LS__SDFRTN_1%CLK_N N_CLK_N_c_530_n N_CLK_N_M1012_g
+ N_CLK_N_M1024_g N_CLK_N_c_531_n N_CLK_N_c_532_n CLK_N
+ PM_SKY130_FD_SC_LS__SDFRTN_1%CLK_N
x_PM_SKY130_FD_SC_LS__SDFRTN_1%A_1049_347# N_A_1049_347#_M1010_d
+ N_A_1049_347#_M1028_d N_A_1049_347#_c_569_n N_A_1049_347#_M1023_g
+ N_A_1049_347#_M1018_g N_A_1049_347#_c_570_n N_A_1049_347#_c_589_n
+ N_A_1049_347#_M1009_g N_A_1049_347#_c_571_n N_A_1049_347#_c_572_n
+ N_A_1049_347#_M1032_g N_A_1049_347#_c_573_n N_A_1049_347#_c_574_n
+ N_A_1049_347#_c_575_n N_A_1049_347#_c_725_p N_A_1049_347#_c_576_n
+ N_A_1049_347#_c_577_n N_A_1049_347#_c_578_n N_A_1049_347#_c_579_n
+ N_A_1049_347#_c_599_p N_A_1049_347#_c_580_n N_A_1049_347#_c_581_n
+ N_A_1049_347#_c_582_n N_A_1049_347#_c_609_p N_A_1049_347#_c_583_n
+ N_A_1049_347#_c_584_n N_A_1049_347#_c_585_n N_A_1049_347#_c_586_n
+ PM_SKY130_FD_SC_LS__SDFRTN_1%A_1049_347#
x_PM_SKY130_FD_SC_LS__SDFRTN_1%A_1402_308# N_A_1402_308#_M1036_d
+ N_A_1402_308#_M1020_d N_A_1402_308#_M1025_g N_A_1402_308#_M1029_g
+ N_A_1402_308#_c_753_n N_A_1402_308#_c_754_n N_A_1402_308#_c_755_n
+ N_A_1402_308#_c_771_n N_A_1402_308#_c_760_n N_A_1402_308#_c_776_n
+ N_A_1402_308#_c_756_n N_A_1402_308#_c_757_n
+ PM_SKY130_FD_SC_LS__SDFRTN_1%A_1402_308#
x_PM_SKY130_FD_SC_LS__SDFRTN_1%RESET_B N_RESET_B_M1039_g N_RESET_B_c_865_n
+ N_RESET_B_c_866_n N_RESET_B_M1026_g N_RESET_B_c_849_n N_RESET_B_M1013_g
+ N_RESET_B_M1011_g N_RESET_B_c_869_n N_RESET_B_M1007_g N_RESET_B_c_852_n
+ N_RESET_B_c_871_n N_RESET_B_M1005_g N_RESET_B_c_872_n N_RESET_B_c_873_n
+ N_RESET_B_c_853_n N_RESET_B_c_854_n N_RESET_B_c_855_n N_RESET_B_c_856_n
+ N_RESET_B_c_857_n RESET_B N_RESET_B_c_858_n N_RESET_B_c_859_n
+ N_RESET_B_c_860_n N_RESET_B_c_861_n N_RESET_B_c_862_n N_RESET_B_c_863_n
+ PM_SKY130_FD_SC_LS__SDFRTN_1%RESET_B
x_PM_SKY130_FD_SC_LS__SDFRTN_1%A_1251_463# N_A_1251_463#_M1023_d
+ N_A_1251_463#_M1004_d N_A_1251_463#_M1013_d N_A_1251_463#_c_1091_n
+ N_A_1251_463#_M1036_g N_A_1251_463#_c_1096_n N_A_1251_463#_M1020_g
+ N_A_1251_463#_c_1097_n N_A_1251_463#_c_1098_n N_A_1251_463#_c_1099_n
+ N_A_1251_463#_c_1092_n N_A_1251_463#_c_1101_n N_A_1251_463#_c_1102_n
+ N_A_1251_463#_c_1103_n N_A_1251_463#_c_1093_n N_A_1251_463#_c_1094_n
+ N_A_1251_463#_c_1095_n N_A_1251_463#_c_1106_n N_A_1251_463#_c_1107_n
+ PM_SKY130_FD_SC_LS__SDFRTN_1%A_1251_463#
x_PM_SKY130_FD_SC_LS__SDFRTN_1%A_854_74# N_A_854_74#_M1012_d N_A_854_74#_M1024_s
+ N_A_854_74#_c_1219_n N_A_854_74#_M1028_g N_A_854_74#_c_1220_n
+ N_A_854_74#_M1010_g N_A_854_74#_c_1221_n N_A_854_74#_M1004_g
+ N_A_854_74#_c_1223_n N_A_854_74#_c_1224_n N_A_854_74#_M1014_g
+ N_A_854_74#_c_1226_n N_A_854_74#_c_1227_n N_A_854_74#_M1038_g
+ N_A_854_74#_c_1229_n N_A_854_74#_c_1244_n N_A_854_74#_M1021_g
+ N_A_854_74#_c_1230_n N_A_854_74#_c_1231_n N_A_854_74#_c_1232_n
+ N_A_854_74#_c_1257_n N_A_854_74#_c_1245_n N_A_854_74#_c_1246_n
+ N_A_854_74#_c_1233_n N_A_854_74#_c_1234_n N_A_854_74#_c_1235_n
+ N_A_854_74#_c_1236_n N_A_854_74#_c_1237_n N_A_854_74#_c_1238_n
+ N_A_854_74#_c_1239_n PM_SKY130_FD_SC_LS__SDFRTN_1%A_854_74#
x_PM_SKY130_FD_SC_LS__SDFRTN_1%A_2087_410# N_A_2087_410#_M1008_d
+ N_A_2087_410#_M1005_d N_A_2087_410#_c_1429_n N_A_2087_410#_M1000_g
+ N_A_2087_410#_M1001_g N_A_2087_410#_c_1431_n N_A_2087_410#_c_1432_n
+ N_A_2087_410#_c_1427_n N_A_2087_410#_c_1433_n N_A_2087_410#_c_1428_n
+ N_A_2087_410#_c_1435_n N_A_2087_410#_c_1436_n
+ PM_SKY130_FD_SC_LS__SDFRTN_1%A_2087_410#
x_PM_SKY130_FD_SC_LS__SDFRTN_1%A_1827_144# N_A_1827_144#_M1038_d
+ N_A_1827_144#_M1009_d N_A_1827_144#_c_1517_n N_A_1827_144#_M1008_g
+ N_A_1827_144#_c_1518_n N_A_1827_144#_c_1519_n N_A_1827_144#_c_1531_n
+ N_A_1827_144#_c_1532_n N_A_1827_144#_M1017_g N_A_1827_144#_c_1533_n
+ N_A_1827_144#_c_1520_n N_A_1827_144#_c_1534_n N_A_1827_144#_M1027_g
+ N_A_1827_144#_c_1521_n N_A_1827_144#_M1033_g N_A_1827_144#_c_1522_n
+ N_A_1827_144#_c_1535_n N_A_1827_144#_c_1536_n N_A_1827_144#_c_1523_n
+ N_A_1827_144#_c_1524_n N_A_1827_144#_c_1537_n N_A_1827_144#_c_1538_n
+ N_A_1827_144#_c_1525_n N_A_1827_144#_c_1526_n N_A_1827_144#_c_1539_n
+ N_A_1827_144#_c_1527_n N_A_1827_144#_c_1528_n N_A_1827_144#_c_1529_n
+ N_A_1827_144#_c_1541_n PM_SKY130_FD_SC_LS__SDFRTN_1%A_1827_144#
x_PM_SKY130_FD_SC_LS__SDFRTN_1%A_2492_424# N_A_2492_424#_M1033_s
+ N_A_2492_424#_M1027_s N_A_2492_424#_c_1681_n N_A_2492_424#_M1006_g
+ N_A_2492_424#_M1015_g N_A_2492_424#_c_1677_n N_A_2492_424#_c_1678_n
+ N_A_2492_424#_c_1679_n N_A_2492_424#_c_1684_n N_A_2492_424#_c_1680_n
+ PM_SKY130_FD_SC_LS__SDFRTN_1%A_2492_424#
x_PM_SKY130_FD_SC_LS__SDFRTN_1%VPWR N_VPWR_M1030_d N_VPWR_M1016_d N_VPWR_M1024_d
+ N_VPWR_M1025_d N_VPWR_M1020_s N_VPWR_M1000_d N_VPWR_M1017_d N_VPWR_M1027_d
+ N_VPWR_c_1722_n N_VPWR_c_1723_n N_VPWR_c_1724_n N_VPWR_c_1725_n
+ N_VPWR_c_1726_n N_VPWR_c_1727_n N_VPWR_c_1728_n N_VPWR_c_1729_n
+ N_VPWR_c_1730_n N_VPWR_c_1731_n VPWR N_VPWR_c_1732_n N_VPWR_c_1733_n
+ N_VPWR_c_1734_n N_VPWR_c_1735_n N_VPWR_c_1736_n N_VPWR_c_1737_n
+ N_VPWR_c_1738_n N_VPWR_c_1721_n N_VPWR_c_1740_n N_VPWR_c_1741_n
+ N_VPWR_c_1742_n N_VPWR_c_1743_n N_VPWR_c_1744_n N_VPWR_c_1745_n
+ PM_SKY130_FD_SC_LS__SDFRTN_1%VPWR
x_PM_SKY130_FD_SC_LS__SDFRTN_1%A_284_464# N_A_284_464#_M1022_d
+ N_A_284_464#_M1023_s N_A_284_464#_M1002_d N_A_284_464#_M1039_d
+ N_A_284_464#_M1004_s N_A_284_464#_c_1877_n N_A_284_464#_c_1887_n
+ N_A_284_464#_c_1861_n N_A_284_464#_c_1862_n N_A_284_464#_c_1863_n
+ N_A_284_464#_c_1868_n N_A_284_464#_c_1869_n N_A_284_464#_c_1870_n
+ N_A_284_464#_c_1871_n N_A_284_464#_c_1946_n N_A_284_464#_c_1864_n
+ N_A_284_464#_c_1865_n N_A_284_464#_c_1953_n N_A_284_464#_c_1873_n
+ N_A_284_464#_c_1874_n N_A_284_464#_c_1875_n N_A_284_464#_c_1866_n
+ N_A_284_464#_c_1884_n N_A_284_464#_c_1889_n N_A_284_464#_c_1867_n
+ N_A_284_464#_c_1876_n PM_SKY130_FD_SC_LS__SDFRTN_1%A_284_464#
x_PM_SKY130_FD_SC_LS__SDFRTN_1%Q N_Q_M1015_d N_Q_M1006_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LS__SDFRTN_1%Q
x_PM_SKY130_FD_SC_LS__SDFRTN_1%VGND N_VGND_M1037_d N_VGND_M1026_d N_VGND_M1010_s
+ N_VGND_M1011_d N_VGND_M1001_d N_VGND_M1033_d N_VGND_c_2036_n N_VGND_c_2037_n
+ N_VGND_c_2038_n N_VGND_c_2039_n VGND N_VGND_c_2040_n N_VGND_c_2041_n
+ N_VGND_c_2042_n N_VGND_c_2043_n N_VGND_c_2044_n N_VGND_c_2045_n
+ N_VGND_c_2046_n N_VGND_c_2047_n N_VGND_c_2048_n N_VGND_c_2049_n
+ N_VGND_c_2050_n N_VGND_c_2051_n N_VGND_c_2052_n N_VGND_c_2053_n
+ PM_SKY130_FD_SC_LS__SDFRTN_1%VGND
x_PM_SKY130_FD_SC_LS__SDFRTN_1%noxref_24 N_noxref_24_M1019_s N_noxref_24_M1034_d
+ N_noxref_24_c_2153_n N_noxref_24_c_2154_n N_noxref_24_c_2155_n
+ N_noxref_24_c_2156_n PM_SKY130_FD_SC_LS__SDFRTN_1%noxref_24
cc_1 VNB N_SCE_M1037_g 0.05663f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_2 VNB N_SCE_c_280_n 0.00333779f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.93
cc_3 VNB N_SCE_M1003_g 0.0185275f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=0.615
cc_4 VNB N_SCE_c_282_n 0.00276011f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.575
cc_5 VNB N_SCE_c_283_n 0.0317758f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.575
cc_6 VNB N_SCE_c_284_n 0.0256442f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=1.267
cc_7 VNB N_SCE_c_285_n 0.00942789f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.267
cc_8 VNB N_SCE_c_286_n 0.0114065f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.12
cc_9 VNB N_SCE_c_287_n 0.046047f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=1.12
cc_10 VNB N_A_27_88#_c_347_n 0.0276281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_88#_c_348_n 0.0210999f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.495
cc_12 VNB N_A_27_88#_c_349_n 0.0146462f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.12
cc_13 VNB N_A_27_88#_c_350_n 0.0108567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_88#_c_351_n 0.00647888f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.182
cc_15 VNB N_A_27_88#_c_352_n 0.03765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_88#_c_353_n 0.0215459f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.182
cc_17 VNB N_A_27_88#_c_354_n 0.0189579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_D_M1022_g 0.0631098f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_19 VNB N_SCD_M1034_g 0.0488825f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_20 VNB SCD 0.00419665f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=0.615
cc_21 VNB N_SCD_c_481_n 0.0148775f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=1.495
cc_22 VNB N_CLK_N_c_530_n 0.0224902f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.41
cc_23 VNB N_CLK_N_c_531_n 0.0189312f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_24 VNB N_CLK_N_c_532_n 0.0482629f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_25 VNB CLK_N 0.0038408f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.245
cc_26 VNB N_A_1049_347#_c_569_n 0.0171643f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.245
cc_27 VNB N_A_1049_347#_c_570_n 0.0292221f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=0.615
cc_28 VNB N_A_1049_347#_c_571_n 0.0299484f $X=-0.19 $Y=-0.245 $X2=1.875
+ $Y2=1.495
cc_29 VNB N_A_1049_347#_c_572_n 0.0175454f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.495
cc_30 VNB N_A_1049_347#_c_573_n 0.00346036f $X=-0.19 $Y=-0.245 $X2=1.875
+ $Y2=1.267
cc_31 VNB N_A_1049_347#_c_574_n 5.54636e-19 $X=-0.19 $Y=-0.245 $X2=2.075
+ $Y2=1.21
cc_32 VNB N_A_1049_347#_c_575_n 0.0097397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_1049_347#_c_576_n 0.00409104f $X=-0.19 $Y=-0.245 $X2=2.385
+ $Y2=1.12
cc_34 VNB N_A_1049_347#_c_577_n 0.0185358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_1049_347#_c_578_n 6.38447e-19 $X=-0.19 $Y=-0.245 $X2=2.16
+ $Y2=1.182
cc_36 VNB N_A_1049_347#_c_579_n 0.00260945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_1049_347#_c_580_n 0.00208056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_1049_347#_c_581_n 6.5087e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1049_347#_c_582_n 0.0598631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1049_347#_c_583_n 0.0067212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1049_347#_c_584_n 0.00134446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1049_347#_c_585_n 6.71187e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1049_347#_c_586_n 0.0435569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1402_308#_M1029_g 0.0306319f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=0.955
cc_45 VNB N_A_1402_308#_c_753_n 0.00394955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1402_308#_c_754_n 0.00749325f $X=-0.19 $Y=-0.245 $X2=0.865
+ $Y2=1.495
cc_47 VNB N_A_1402_308#_c_755_n 0.00266045f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.495
cc_48 VNB N_A_1402_308#_c_756_n 0.00342912f $X=-0.19 $Y=-0.245 $X2=2.385
+ $Y2=1.12
cc_49 VNB N_A_1402_308#_c_757_n 0.0335457f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.182
cc_50 VNB N_RESET_B_M1026_g 0.0431367f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_51 VNB N_RESET_B_c_849_n 0.0102324f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_52 VNB N_RESET_B_M1011_g 0.0318942f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=1.495
cc_53 VNB N_RESET_B_M1007_g 0.0335346f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=1.267
cc_54 VNB N_RESET_B_c_852_n 0.0059249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_RESET_B_c_853_n 0.014478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_RESET_B_c_854_n 4.19263e-19 $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.182
cc_57 VNB N_RESET_B_c_855_n 0.0163609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_RESET_B_c_856_n 8.92608e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_RESET_B_c_857_n 0.00211188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_RESET_B_c_858_n 0.0193532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_RESET_B_c_859_n 0.00168181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_RESET_B_c_860_n 0.0215933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_RESET_B_c_861_n 0.00325463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_RESET_B_c_862_n 0.0293012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_RESET_B_c_863_n 0.00974625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1251_463#_c_1091_n 0.0195095f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.245
cc_67 VNB N_A_1251_463#_c_1092_n 0.00700528f $X=-0.19 $Y=-0.245 $X2=0.7
+ $Y2=1.575
cc_68 VNB N_A_1251_463#_c_1093_n 0.0013425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1251_463#_c_1094_n 0.0363897f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=1.12
cc_70 VNB N_A_1251_463#_c_1095_n 0.00235971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_854_74#_c_1219_n 0.0258783f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_72 VNB N_A_854_74#_c_1220_n 0.0221872f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_73 VNB N_A_854_74#_c_1221_n 0.0484145f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=0.615
cc_74 VNB N_A_854_74#_M1004_g 0.0191872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_854_74#_c_1223_n 0.0180995f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.495
cc_76 VNB N_A_854_74#_c_1224_n 0.019091f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.575
cc_77 VNB N_A_854_74#_M1014_g 0.0246129f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_78 VNB N_A_854_74#_c_1226_n 0.151323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_854_74#_c_1227_n 0.0102922f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.575
cc_80 VNB N_A_854_74#_M1038_g 0.0450814f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.12
cc_81 VNB N_A_854_74#_c_1229_n 0.00591217f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=1.12
cc_82 VNB N_A_854_74#_c_1230_n 0.0058413f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.182
cc_83 VNB N_A_854_74#_c_1231_n 0.0238216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_854_74#_c_1232_n 0.00590081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_854_74#_c_1233_n 0.00273923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_854_74#_c_1234_n 0.00193318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_854_74#_c_1235_n 0.006264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_854_74#_c_1236_n 0.0237946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_854_74#_c_1237_n 0.00312043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_854_74#_c_1238_n 0.0320997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_854_74#_c_1239_n 0.00932697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2087_410#_M1001_g 0.0627011f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_93 VNB N_A_2087_410#_c_1427_n 0.00234211f $X=-0.19 $Y=-0.245 $X2=0.865
+ $Y2=1.495
cc_94 VNB N_A_2087_410#_c_1428_n 0.0133151f $X=-0.19 $Y=-0.245 $X2=2.075
+ $Y2=1.21
cc_95 VNB N_A_1827_144#_c_1517_n 0.0218114f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.245
cc_96 VNB N_A_1827_144#_c_1518_n 0.0200739f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.64
cc_97 VNB N_A_1827_144#_c_1519_n 0.00490842f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=0.955
cc_98 VNB N_A_1827_144#_c_1520_n 0.0770594f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.495
cc_99 VNB N_A_1827_144#_c_1521_n 0.0208776f $X=-0.19 $Y=-0.245 $X2=2.045
+ $Y2=1.267
cc_100 VNB N_A_1827_144#_c_1522_n 0.0175897f $X=-0.19 $Y=-0.245 $X2=0.642
+ $Y2=1.575
cc_101 VNB N_A_1827_144#_c_1523_n 0.00222143f $X=-0.19 $Y=-0.245 $X2=2.385
+ $Y2=1.182
cc_102 VNB N_A_1827_144#_c_1524_n 0.00135104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1827_144#_c_1525_n 0.0381536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1827_144#_c_1526_n 0.00146089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1827_144#_c_1527_n 0.00113131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1827_144#_c_1528_n 0.0199884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1827_144#_c_1529_n 0.0106578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_2492_424#_M1015_g 0.0336704f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.64
cc_109 VNB N_A_2492_424#_c_1677_n 0.0509652f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=0.615
cc_110 VNB N_A_2492_424#_c_1678_n 0.0161427f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=0.615
cc_111 VNB N_A_2492_424#_c_1679_n 0.0173592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2492_424#_c_1680_n 0.00257436f $X=-0.19 $Y=-0.245 $X2=1.875
+ $Y2=1.267
cc_113 VNB N_VPWR_c_1721_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_284_464#_c_1861_n 0.00320002f $X=-0.19 $Y=-0.245 $X2=1.875
+ $Y2=1.267
cc_115 VNB N_A_284_464#_c_1862_n 0.0213865f $X=-0.19 $Y=-0.245 $X2=2.045
+ $Y2=1.267
cc_116 VNB N_A_284_464#_c_1863_n 0.00512961f $X=-0.19 $Y=-0.245 $X2=2.075
+ $Y2=1.21
cc_117 VNB N_A_284_464#_c_1864_n 0.00764057f $X=-0.19 $Y=-0.245 $X2=2.16
+ $Y2=1.182
cc_118 VNB N_A_284_464#_c_1865_n 0.0180549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_284_464#_c_1866_n 0.00676717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_284_464#_c_1867_n 0.00123517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB Q 0.0545639f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_122 VNB N_VGND_c_2036_n 0.0212574f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.495
cc_123 VNB N_VGND_c_2037_n 0.0160815f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=1.267
cc_124 VNB N_VGND_c_2038_n 0.00450109f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.575
cc_125 VNB N_VGND_c_2039_n 0.015381f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.12
cc_126 VNB N_VGND_c_2040_n 0.0194805f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.182
cc_127 VNB N_VGND_c_2041_n 0.0194733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2042_n 0.0667461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2043_n 0.0701843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2044_n 0.0500113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2045_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2046_n 0.73935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2047_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2048_n 0.0627249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2049_n 0.0175441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2050_n 0.0157128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2051_n 0.00461401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2052_n 0.00865198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2053_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_noxref_24_c_2153_n 0.00347762f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.64
cc_141 VNB N_noxref_24_c_2154_n 0.0148058f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_142 VNB N_noxref_24_c_2155_n 0.00461646f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.64
cc_143 VNB N_noxref_24_c_2156_n 0.0026427f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=0.615
cc_144 VPB N_SCE_c_280_n 0.0785994f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.93
cc_145 VPB N_SCE_c_289_n 0.0331559f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_146 VPB N_SCE_c_282_n 0.00272259f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.575
cc_147 VPB N_A_27_88#_c_355_n 0.0150795f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_148 VPB N_A_27_88#_c_356_n 0.0281089f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_149 VPB N_A_27_88#_c_348_n 0.0319763f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.495
cc_150 VPB N_A_27_88#_c_358_n 0.0214794f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.575
cc_151 VPB N_A_27_88#_c_359_n 0.0184521f $X=-0.19 $Y=1.66 $X2=1.875 $Y2=1.267
cc_152 VPB N_A_27_88#_c_360_n 0.00325282f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.12
cc_153 VPB N_A_27_88#_c_349_n 0.021371f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.12
cc_154 VPB N_A_27_88#_c_362_n 0.00717703f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=1.12
cc_155 VPB N_D_c_440_n 0.0206307f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.41
cc_156 VPB N_D_c_441_n 0.0146877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_D_M1022_g 0.00943149f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_158 VPB N_D_c_443_n 0.0205457f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.245
cc_159 VPB N_D_c_444_n 0.0336862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_D_c_445_n 0.0162449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_SCD_c_482_n 0.0169752f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.41
cc_162 VPB N_SCD_c_483_n 0.0136324f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.632
cc_163 VPB N_SCD_c_484_n 0.0287642f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_164 VPB SCD 0.00642005f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=0.615
cc_165 VPB N_SCD_c_481_n 0.0178291f $X=-0.19 $Y=1.66 $X2=1.875 $Y2=1.495
cc_166 VPB N_CLK_N_M1024_g 0.0239999f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.93
cc_167 VPB N_A_1049_347#_M1018_g 0.0227189f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_168 VPB N_A_1049_347#_c_570_n 7.86941e-19 $X=-0.19 $Y=1.66 $X2=2.615
+ $Y2=0.615
cc_169 VPB N_A_1049_347#_c_589_n 0.028997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_1049_347#_c_574_n 0.00547365f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.21
cc_171 VPB N_A_1049_347#_c_583_n 0.0224997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_1049_347#_c_584_n 0.0106238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_1402_308#_M1025_g 0.0317208f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_174 VPB N_A_1402_308#_c_753_n 0.00228499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_1402_308#_c_760_n 0.00695194f $X=-0.19 $Y=1.66 $X2=2.045
+ $Y2=1.267
cc_176 VPB N_A_1402_308#_c_756_n 0.00190176f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.12
cc_177 VPB N_A_1402_308#_c_757_n 0.0153161f $X=-0.19 $Y=1.66 $X2=2.16 $Y2=1.182
cc_178 VPB N_RESET_B_M1039_g 0.0141325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_RESET_B_c_865_n 0.329154f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.632
cc_180 VPB N_RESET_B_c_866_n 0.0124423f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.93
cc_181 VPB N_RESET_B_c_849_n 0.0672676f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_182 VPB N_RESET_B_M1013_g 0.0277424f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_RESET_B_c_869_n 0.0180429f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.575
cc_184 VPB N_RESET_B_c_852_n 0.0349147f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_RESET_B_c_871_n 0.017636f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.575
cc_186 VPB N_RESET_B_c_872_n 0.0258265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_RESET_B_c_873_n 0.0150132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_RESET_B_c_853_n 0.0193653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_RESET_B_c_854_n 4.25177e-19 $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.182
cc_190 VPB N_RESET_B_c_855_n 0.00114121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_RESET_B_c_856_n 2.20672e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_RESET_B_c_857_n 0.00221319f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_RESET_B_c_859_n 0.00266259f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_RESET_B_c_860_n 0.00543554f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_RESET_B_c_861_n 4.3193e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_RESET_B_c_863_n 6.46864e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1251_463#_c_1096_n 0.0211423f $X=-0.19 $Y=1.66 $X2=2.615
+ $Y2=0.955
cc_198 VPB N_A_1251_463#_c_1097_n 0.00155811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1251_463#_c_1098_n 0.00202538f $X=-0.19 $Y=1.66 $X2=0.865
+ $Y2=1.495
cc_200 VPB N_A_1251_463#_c_1099_n 0.00296853f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.495
cc_201 VPB N_A_1251_463#_c_1092_n 0.00150835f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.575
cc_202 VPB N_A_1251_463#_c_1101_n 0.0088739f $X=-0.19 $Y=1.66 $X2=2.045
+ $Y2=1.182
cc_203 VPB N_A_1251_463#_c_1102_n 0.00993973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_1251_463#_c_1103_n 0.0171747f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.41
cc_205 VPB N_A_1251_463#_c_1093_n 0.00303633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_1251_463#_c_1094_n 0.0191822f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=1.12
cc_207 VPB N_A_1251_463#_c_1106_n 0.00194613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_1251_463#_c_1107_n 0.00407506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_854_74#_c_1219_n 0.00635671f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_210 VPB N_A_854_74#_M1028_g 0.0225247f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_211 VPB N_A_854_74#_M1004_g 0.0485335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_854_74#_c_1229_n 0.0379367f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=1.12
cc_213 VPB N_A_854_74#_c_1244_n 0.0217507f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_854_74#_c_1245_n 0.00251318f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_854_74#_c_1246_n 0.0024675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_854_74#_c_1233_n 0.00133445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_854_74#_c_1235_n 0.00313142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_854_74#_c_1236_n 0.0107083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_2087_410#_c_1429_n 0.0562969f $X=-0.19 $Y=1.66 $X2=0.505
+ $Y2=2.245
cc_220 VPB N_A_2087_410#_M1001_g 0.0217533f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_221 VPB N_A_2087_410#_c_1431_n 0.010007f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=0.615
cc_222 VPB N_A_2087_410#_c_1432_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_2087_410#_c_1433_n 0.010671f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=1.182
cc_224 VPB N_A_2087_410#_c_1428_n 0.00836152f $X=-0.19 $Y=1.66 $X2=2.075
+ $Y2=1.21
cc_225 VPB N_A_2087_410#_c_1435_n 0.00347726f $X=-0.19 $Y=1.66 $X2=0.642
+ $Y2=1.575
cc_226 VPB N_A_2087_410#_c_1436_n 0.00251499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1827_144#_c_1519_n 0.0140687f $X=-0.19 $Y=1.66 $X2=2.615
+ $Y2=0.955
cc_228 VPB N_A_1827_144#_c_1531_n 0.0206982f $X=-0.19 $Y=1.66 $X2=2.615
+ $Y2=0.615
cc_229 VPB N_A_1827_144#_c_1532_n 0.0233137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_1827_144#_c_1533_n 0.0748364f $X=-0.19 $Y=1.66 $X2=1.875
+ $Y2=1.495
cc_231 VPB N_A_1827_144#_c_1534_n 0.0189909f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.575
cc_232 VPB N_A_1827_144#_c_1535_n 0.00569915f $X=-0.19 $Y=1.66 $X2=0.642
+ $Y2=1.41
cc_233 VPB N_A_1827_144#_c_1536_n 0.00407057f $X=-0.19 $Y=1.66 $X2=2.615
+ $Y2=1.12
cc_234 VPB N_A_1827_144#_c_1537_n 0.013426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_1827_144#_c_1538_n 0.00333305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_1827_144#_c_1539_n 0.01246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_1827_144#_c_1527_n 0.0041497f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_1827_144#_c_1541_n 0.0081065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_2492_424#_c_1681_n 0.0211258f $X=-0.19 $Y=1.66 $X2=0.505
+ $Y2=2.245
cc_240 VPB N_A_2492_424#_c_1677_n 0.0194078f $X=-0.19 $Y=1.66 $X2=2.615
+ $Y2=0.615
cc_241 VPB N_A_2492_424#_c_1678_n 0.0085619f $X=-0.19 $Y=1.66 $X2=2.615
+ $Y2=0.615
cc_242 VPB N_A_2492_424#_c_1684_n 0.0163308f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.575
cc_243 VPB N_A_2492_424#_c_1680_n 3.52822e-19 $X=-0.19 $Y=1.66 $X2=1.875
+ $Y2=1.267
cc_244 VPB N_VPWR_c_1722_n 0.00396467f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.21
cc_245 VPB N_VPWR_c_1723_n 0.0161419f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.12
cc_246 VPB N_VPWR_c_1724_n 0.0129753f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=1.12
cc_247 VPB N_VPWR_c_1725_n 0.0163398f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.182
cc_248 VPB N_VPWR_c_1726_n 0.012683f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1727_n 0.0160012f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1728_n 0.0625388f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1729_n 0.00223798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1730_n 0.0187266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1731_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1732_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1733_n 0.0518169f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1734_n 0.0477117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1735_n 0.0257316f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1736_n 0.054077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1737_n 0.0215226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1738_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1721_n 0.133324f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1740_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1741_n 0.0139505f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1742_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1743_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1744_n 0.0201883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1745_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_A_284_464#_c_1868_n 0.0153439f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.575
cc_269 VPB N_A_284_464#_c_1869_n 0.00853637f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.12
cc_270 VPB N_A_284_464#_c_1870_n 0.00772972f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.12
cc_271 VPB N_A_284_464#_c_1871_n 0.00169858f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.12
cc_272 VPB N_A_284_464#_c_1864_n 0.0147324f $X=-0.19 $Y=1.66 $X2=2.16 $Y2=1.182
cc_273 VPB N_A_284_464#_c_1873_n 0.0074538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_284_464#_c_1874_n 0.0152378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_A_284_464#_c_1875_n 0.00161322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_284_464#_c_1876_n 0.00471545f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB Q 0.0536464f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_278 N_SCE_M1037_g N_A_27_88#_c_347_n 0.0173492f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_279 N_SCE_M1037_g N_A_27_88#_c_348_n 0.0255944f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_280 N_SCE_c_280_n N_A_27_88#_c_348_n 0.00687726f $X=0.642 $Y=1.93 $X2=0 $Y2=0
cc_281 N_SCE_c_289_n N_A_27_88#_c_348_n 0.00176852f $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_282 N_SCE_c_282_n N_A_27_88#_c_348_n 0.0525665f $X=0.7 $Y=1.575 $X2=0 $Y2=0
cc_283 N_SCE_c_289_n N_A_27_88#_c_358_n 0.00517645f $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_284 N_SCE_c_280_n N_A_27_88#_c_359_n 0.00421788f $X=0.642 $Y=1.93 $X2=0 $Y2=0
cc_285 N_SCE_c_289_n N_A_27_88#_c_359_n 0.0346587f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_286 N_SCE_c_282_n N_A_27_88#_c_359_n 0.0221414f $X=0.7 $Y=1.575 $X2=0 $Y2=0
cc_287 N_SCE_c_286_n N_A_27_88#_c_360_n 0.0282051f $X=2.385 $Y=1.12 $X2=0 $Y2=0
cc_288 N_SCE_c_287_n N_A_27_88#_c_360_n 3.15902e-19 $X=2.615 $Y=1.12 $X2=0 $Y2=0
cc_289 N_SCE_c_285_n N_A_27_88#_c_349_n 6.75701e-19 $X=2.045 $Y=1.267 $X2=0
+ $Y2=0
cc_290 N_SCE_c_286_n N_A_27_88#_c_349_n 0.00372722f $X=2.385 $Y=1.12 $X2=0 $Y2=0
cc_291 N_SCE_c_287_n N_A_27_88#_c_349_n 0.0150169f $X=2.615 $Y=1.12 $X2=0 $Y2=0
cc_292 N_SCE_M1037_g N_A_27_88#_c_350_n 0.00558381f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_293 N_SCE_c_285_n N_A_27_88#_c_351_n 0.016963f $X=2.045 $Y=1.267 $X2=0 $Y2=0
cc_294 N_SCE_M1037_g N_A_27_88#_c_352_n 0.00404033f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_295 N_SCE_c_284_n N_A_27_88#_c_352_n 0.00396344f $X=1.875 $Y=1.267 $X2=0
+ $Y2=0
cc_296 N_SCE_c_285_n N_A_27_88#_c_352_n 4.95772e-19 $X=2.045 $Y=1.267 $X2=0
+ $Y2=0
cc_297 N_SCE_M1037_g N_A_27_88#_c_353_n 0.0161451f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_298 N_SCE_c_282_n N_A_27_88#_c_353_n 0.0264209f $X=0.7 $Y=1.575 $X2=0 $Y2=0
cc_299 N_SCE_c_283_n N_A_27_88#_c_353_n 0.00207087f $X=0.7 $Y=1.575 $X2=0 $Y2=0
cc_300 N_SCE_c_284_n N_A_27_88#_c_353_n 0.0568522f $X=1.875 $Y=1.267 $X2=0 $Y2=0
cc_301 N_SCE_c_289_n N_D_c_440_n 0.044837f $X=0.505 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_302 N_SCE_M1003_g N_D_M1022_g 0.0146952f $X=2.615 $Y=0.615 $X2=0 $Y2=0
cc_303 N_SCE_c_284_n N_D_M1022_g 0.00734487f $X=1.875 $Y=1.267 $X2=0 $Y2=0
cc_304 N_SCE_c_285_n N_D_M1022_g 0.027662f $X=2.045 $Y=1.267 $X2=0 $Y2=0
cc_305 N_SCE_c_287_n N_D_M1022_g 0.0181201f $X=2.615 $Y=1.12 $X2=0 $Y2=0
cc_306 N_SCE_c_280_n N_D_c_443_n 0.0186437f $X=0.642 $Y=1.93 $X2=0 $Y2=0
cc_307 N_SCE_c_284_n N_D_c_443_n 0.00120387f $X=1.875 $Y=1.267 $X2=0 $Y2=0
cc_308 N_SCE_c_280_n N_D_c_444_n 3.94848e-19 $X=0.642 $Y=1.93 $X2=0 $Y2=0
cc_309 N_SCE_c_284_n N_D_c_444_n 0.00395715f $X=1.875 $Y=1.267 $X2=0 $Y2=0
cc_310 N_SCE_c_280_n N_D_c_445_n 0.00644204f $X=0.642 $Y=1.93 $X2=0 $Y2=0
cc_311 N_SCE_c_282_n N_D_c_445_n 0.0207563f $X=0.7 $Y=1.575 $X2=0 $Y2=0
cc_312 N_SCE_c_284_n N_D_c_445_n 0.0621482f $X=1.875 $Y=1.267 $X2=0 $Y2=0
cc_313 N_SCE_M1003_g N_SCD_M1034_g 0.0515549f $X=2.615 $Y=0.615 $X2=0 $Y2=0
cc_314 N_SCE_c_286_n N_SCD_M1034_g 0.00466427f $X=2.385 $Y=1.12 $X2=0 $Y2=0
cc_315 N_SCE_c_289_n N_VPWR_c_1722_n 0.0201296f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_316 N_SCE_c_289_n N_VPWR_c_1732_n 0.00413917f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_317 N_SCE_c_289_n N_VPWR_c_1733_n 0.00413917f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_318 N_SCE_c_289_n N_VPWR_c_1721_n 0.0163846f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_319 N_SCE_M1003_g N_A_284_464#_c_1877_n 0.0148189f $X=2.615 $Y=0.615 $X2=0
+ $Y2=0
cc_320 N_SCE_c_285_n N_A_284_464#_c_1877_n 0.0386304f $X=2.045 $Y=1.267 $X2=0
+ $Y2=0
cc_321 N_SCE_c_287_n N_A_284_464#_c_1877_n 0.00694878f $X=2.615 $Y=1.12 $X2=0
+ $Y2=0
cc_322 N_SCE_M1003_g N_A_284_464#_c_1861_n 0.00382794f $X=2.615 $Y=0.615 $X2=0
+ $Y2=0
cc_323 N_SCE_c_286_n N_A_284_464#_c_1861_n 0.0046738f $X=2.385 $Y=1.12 $X2=0
+ $Y2=0
cc_324 N_SCE_c_286_n N_A_284_464#_c_1863_n 0.0151459f $X=2.385 $Y=1.12 $X2=0
+ $Y2=0
cc_325 N_SCE_c_287_n N_A_284_464#_c_1863_n 0.00154341f $X=2.615 $Y=1.12 $X2=0
+ $Y2=0
cc_326 N_SCE_c_289_n N_A_284_464#_c_1884_n 9.1451e-19 $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_327 N_SCE_M1037_g N_VGND_c_2036_n 0.0137116f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_328 N_SCE_M1037_g N_VGND_c_2040_n 0.00504315f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_329 N_SCE_M1037_g N_VGND_c_2046_n 0.00523671f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_330 N_SCE_M1003_g N_VGND_c_2048_n 9.15902e-19 $X=2.615 $Y=0.615 $X2=0 $Y2=0
cc_331 N_SCE_M1003_g N_noxref_24_c_2154_n 0.0105907f $X=2.615 $Y=0.615 $X2=0
+ $Y2=0
cc_332 N_SCE_c_285_n N_noxref_24_c_2154_n 0.00237332f $X=2.045 $Y=1.267 $X2=0
+ $Y2=0
cc_333 N_SCE_M1003_g N_noxref_24_c_2156_n 9.86067e-19 $X=2.615 $Y=0.615 $X2=0
+ $Y2=0
cc_334 N_A_27_88#_c_359_n N_D_c_440_n 0.0161468f $X=2.215 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_335 N_A_27_88#_c_359_n N_D_c_441_n 0.00373424f $X=2.215 $Y=2.375 $X2=0 $Y2=0
cc_336 N_A_27_88#_c_360_n N_D_M1022_g 0.00125677f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_337 N_A_27_88#_c_349_n N_D_M1022_g 0.0173599f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_338 N_A_27_88#_c_351_n N_D_M1022_g 0.00101912f $X=1.455 $Y=1.1 $X2=0 $Y2=0
cc_339 N_A_27_88#_c_354_n N_D_M1022_g 0.0606403f $X=1.455 $Y=0.935 $X2=0 $Y2=0
cc_340 N_A_27_88#_c_359_n N_D_c_443_n 7.57779e-19 $X=2.215 $Y=2.375 $X2=0 $Y2=0
cc_341 N_A_27_88#_c_352_n N_D_c_443_n 0.0032894f $X=1.455 $Y=1.1 $X2=0 $Y2=0
cc_342 N_A_27_88#_c_355_n N_D_c_444_n 0.0173599f $X=2.28 $Y=2.155 $X2=0 $Y2=0
cc_343 N_A_27_88#_c_360_n N_D_c_444_n 3.97221e-19 $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_344 N_A_27_88#_c_359_n N_D_c_445_n 0.0698127f $X=2.215 $Y=2.375 $X2=0 $Y2=0
cc_345 N_A_27_88#_c_360_n N_D_c_445_n 0.0208146f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_346 N_A_27_88#_c_349_n N_D_c_445_n 0.00108531f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_347 N_A_27_88#_c_356_n N_SCD_c_482_n 0.0453956f $X=2.28 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_348 N_A_27_88#_c_359_n N_SCD_c_482_n 0.00143143f $X=2.215 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_349 N_A_27_88#_c_360_n N_SCD_c_482_n 0.00117622f $X=2.38 $Y=1.72 $X2=-0.19
+ $Y2=-0.245
cc_350 N_A_27_88#_c_355_n N_SCD_c_483_n 0.00468854f $X=2.28 $Y=2.155 $X2=0 $Y2=0
cc_351 N_A_27_88#_c_360_n N_SCD_c_483_n 0.0015238f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_352 N_A_27_88#_c_355_n N_SCD_c_484_n 0.00926518f $X=2.28 $Y=2.155 $X2=0 $Y2=0
cc_353 N_A_27_88#_c_360_n N_SCD_c_484_n 0.0031165f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_354 N_A_27_88#_c_355_n SCD 2.48643e-19 $X=2.28 $Y=2.155 $X2=0 $Y2=0
cc_355 N_A_27_88#_c_360_n SCD 0.0326702f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_356 N_A_27_88#_c_349_n SCD 0.00133605f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_357 N_A_27_88#_c_360_n N_SCD_c_481_n 0.00113065f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_358 N_A_27_88#_c_349_n N_SCD_c_481_n 0.0160213f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_359 N_A_27_88#_c_359_n N_VPWR_M1030_d 0.00197722f $X=2.215 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_360 N_A_27_88#_c_358_n N_VPWR_c_1722_n 0.0234974f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_361 N_A_27_88#_c_359_n N_VPWR_c_1722_n 0.0171813f $X=2.215 $Y=2.375 $X2=0
+ $Y2=0
cc_362 N_A_27_88#_c_358_n N_VPWR_c_1732_n 0.011066f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_363 N_A_27_88#_c_356_n N_VPWR_c_1733_n 0.00361401f $X=2.28 $Y=2.245 $X2=0
+ $Y2=0
cc_364 N_A_27_88#_c_356_n N_VPWR_c_1721_n 0.00564686f $X=2.28 $Y=2.245 $X2=0
+ $Y2=0
cc_365 N_A_27_88#_c_358_n N_VPWR_c_1721_n 0.00915947f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_366 N_A_27_88#_c_359_n A_206_464# 0.0048076f $X=2.215 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_367 N_A_27_88#_c_359_n N_A_284_464#_M1002_d 0.0104201f $X=2.215 $Y=2.375
+ $X2=0 $Y2=0
cc_368 N_A_27_88#_c_354_n N_A_284_464#_c_1877_n 4.55233e-19 $X=1.455 $Y=0.935
+ $X2=0 $Y2=0
cc_369 N_A_27_88#_c_356_n N_A_284_464#_c_1887_n 0.00720935f $X=2.28 $Y=2.245
+ $X2=0 $Y2=0
cc_370 N_A_27_88#_c_359_n N_A_284_464#_c_1884_n 0.0529153f $X=2.215 $Y=2.375
+ $X2=0 $Y2=0
cc_371 N_A_27_88#_c_356_n N_A_284_464#_c_1889_n 0.00338647f $X=2.28 $Y=2.245
+ $X2=0 $Y2=0
cc_372 N_A_27_88#_c_359_n N_A_284_464#_c_1889_n 0.0212534f $X=2.215 $Y=2.375
+ $X2=0 $Y2=0
cc_373 N_A_27_88#_c_359_n A_471_464# 0.00139778f $X=2.215 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_374 N_A_27_88#_c_347_n N_VGND_c_2036_n 0.0188413f $X=0.28 $Y=0.65 $X2=0 $Y2=0
cc_375 N_A_27_88#_c_353_n N_VGND_c_2036_n 0.0279144f $X=1.29 $Y=1.087 $X2=0
+ $Y2=0
cc_376 N_A_27_88#_c_354_n N_VGND_c_2036_n 0.00400291f $X=1.455 $Y=0.935 $X2=0
+ $Y2=0
cc_377 N_A_27_88#_c_347_n N_VGND_c_2040_n 0.0113438f $X=0.28 $Y=0.65 $X2=0 $Y2=0
cc_378 N_A_27_88#_c_347_n N_VGND_c_2046_n 0.011567f $X=0.28 $Y=0.65 $X2=0 $Y2=0
cc_379 N_A_27_88#_c_354_n N_VGND_c_2048_n 9.34861e-19 $X=1.455 $Y=0.935 $X2=0
+ $Y2=0
cc_380 N_A_27_88#_c_351_n N_noxref_24_c_2153_n 0.0138157f $X=1.455 $Y=1.1 $X2=0
+ $Y2=0
cc_381 N_A_27_88#_c_352_n N_noxref_24_c_2153_n 0.00399118f $X=1.455 $Y=1.1 $X2=0
+ $Y2=0
cc_382 N_A_27_88#_c_353_n N_noxref_24_c_2153_n 0.00699077f $X=1.29 $Y=1.087
+ $X2=0 $Y2=0
cc_383 N_A_27_88#_c_354_n N_noxref_24_c_2153_n 0.0059422f $X=1.455 $Y=0.935
+ $X2=0 $Y2=0
cc_384 N_A_27_88#_c_351_n N_noxref_24_c_2154_n 0.00360351f $X=1.455 $Y=1.1 $X2=0
+ $Y2=0
cc_385 N_A_27_88#_c_354_n N_noxref_24_c_2154_n 0.00794258f $X=1.455 $Y=0.935
+ $X2=0 $Y2=0
cc_386 N_A_27_88#_c_354_n N_noxref_24_c_2155_n 0.00331383f $X=1.455 $Y=0.935
+ $X2=0 $Y2=0
cc_387 N_D_c_440_n N_VPWR_c_1722_n 0.00157508f $X=1.345 $Y=2.245 $X2=0 $Y2=0
cc_388 N_D_c_440_n N_VPWR_c_1733_n 0.00444752f $X=1.345 $Y=2.245 $X2=0 $Y2=0
cc_389 N_D_c_440_n N_VPWR_c_1721_n 0.00859236f $X=1.345 $Y=2.245 $X2=0 $Y2=0
cc_390 N_D_M1022_g N_A_284_464#_c_1877_n 0.00653506f $X=1.905 $Y=0.615 $X2=0
+ $Y2=0
cc_391 N_D_c_440_n N_A_284_464#_c_1884_n 0.00569115f $X=1.345 $Y=2.245 $X2=0
+ $Y2=0
cc_392 N_D_M1022_g N_VGND_c_2048_n 9.15902e-19 $X=1.905 $Y=0.615 $X2=0 $Y2=0
cc_393 N_D_M1022_g N_noxref_24_c_2153_n 0.00131656f $X=1.905 $Y=0.615 $X2=0
+ $Y2=0
cc_394 N_D_M1022_g N_noxref_24_c_2154_n 0.0127325f $X=1.905 $Y=0.615 $X2=0 $Y2=0
cc_395 N_SCD_c_482_n N_RESET_B_M1039_g 0.0198603f $X=2.67 $Y=2.245 $X2=0 $Y2=0
cc_396 N_SCD_M1034_g N_RESET_B_M1026_g 0.0389277f $X=3.005 $Y=0.615 $X2=0 $Y2=0
cc_397 N_SCD_c_483_n N_RESET_B_c_849_n 0.00563201f $X=2.875 $Y=2.095 $X2=0 $Y2=0
cc_398 N_SCD_c_484_n N_RESET_B_c_849_n 0.0084254f $X=2.875 $Y=2.17 $X2=0 $Y2=0
cc_399 SCD N_RESET_B_c_849_n 0.00354804f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_400 SCD N_RESET_B_c_854_n 0.00160474f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_401 SCD N_RESET_B_c_858_n 0.00478487f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_402 N_SCD_c_481_n N_RESET_B_c_858_n 0.0173672f $X=2.965 $Y=1.69 $X2=0 $Y2=0
cc_403 N_SCD_M1034_g N_RESET_B_c_859_n 9.76155e-19 $X=3.005 $Y=0.615 $X2=0 $Y2=0
cc_404 SCD N_RESET_B_c_859_n 0.0388123f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_405 N_SCD_c_481_n N_RESET_B_c_859_n 3.23745e-19 $X=2.965 $Y=1.69 $X2=0 $Y2=0
cc_406 N_SCD_c_482_n N_VPWR_c_1733_n 0.00314375f $X=2.67 $Y=2.245 $X2=0 $Y2=0
cc_407 N_SCD_c_482_n N_VPWR_c_1721_n 0.00390183f $X=2.67 $Y=2.245 $X2=0 $Y2=0
cc_408 N_SCD_c_482_n N_VPWR_c_1741_n 0.00343384f $X=2.67 $Y=2.245 $X2=0 $Y2=0
cc_409 N_SCD_c_482_n N_A_284_464#_c_1887_n 0.0158977f $X=2.67 $Y=2.245 $X2=0
+ $Y2=0
cc_410 N_SCD_c_484_n N_A_284_464#_c_1887_n 0.00417458f $X=2.875 $Y=2.17 $X2=0
+ $Y2=0
cc_411 SCD N_A_284_464#_c_1887_n 0.0151519f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_412 N_SCD_M1034_g N_A_284_464#_c_1861_n 0.00437851f $X=3.005 $Y=0.615 $X2=0
+ $Y2=0
cc_413 N_SCD_M1034_g N_A_284_464#_c_1862_n 0.0124676f $X=3.005 $Y=0.615 $X2=0
+ $Y2=0
cc_414 SCD N_A_284_464#_c_1862_n 0.0161025f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_415 N_SCD_c_481_n N_A_284_464#_c_1862_n 5.41371e-19 $X=2.965 $Y=1.69 $X2=0
+ $Y2=0
cc_416 SCD N_A_284_464#_c_1863_n 0.00463754f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_417 N_SCD_c_481_n N_A_284_464#_c_1863_n 6.23418e-19 $X=2.965 $Y=1.69 $X2=0
+ $Y2=0
cc_418 N_SCD_c_484_n N_A_284_464#_c_1871_n 2.21134e-19 $X=2.875 $Y=2.17 $X2=0
+ $Y2=0
cc_419 SCD N_A_284_464#_c_1864_n 0.00365391f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_420 N_SCD_c_482_n N_A_284_464#_c_1889_n 7.6548e-19 $X=2.67 $Y=2.245 $X2=0
+ $Y2=0
cc_421 N_SCD_M1034_g N_VGND_c_2048_n 9.34905e-19 $X=3.005 $Y=0.615 $X2=0 $Y2=0
cc_422 N_SCD_M1034_g N_noxref_24_c_2154_n 0.0109613f $X=3.005 $Y=0.615 $X2=0
+ $Y2=0
cc_423 N_SCD_M1034_g N_noxref_24_c_2156_n 0.00602784f $X=3.005 $Y=0.615 $X2=0
+ $Y2=0
cc_424 N_CLK_N_M1024_g N_RESET_B_c_865_n 0.0103562f $X=4.72 $Y=2.235 $X2=0 $Y2=0
cc_425 N_CLK_N_c_530_n N_RESET_B_M1026_g 0.0154061f $X=4.195 $Y=1.22 $X2=0 $Y2=0
cc_426 N_CLK_N_M1024_g N_RESET_B_c_853_n 0.00680016f $X=4.72 $Y=2.235 $X2=0
+ $Y2=0
cc_427 N_CLK_N_c_531_n N_RESET_B_c_853_n 0.0142169f $X=4.27 $Y=1.385 $X2=0 $Y2=0
cc_428 CLK_N N_RESET_B_c_853_n 0.012286f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_429 N_CLK_N_c_531_n N_RESET_B_c_858_n 0.00553134f $X=4.27 $Y=1.385 $X2=0
+ $Y2=0
cc_430 N_CLK_N_c_532_n N_A_854_74#_c_1219_n 0.0213223f $X=4.645 $Y=1.385 $X2=0
+ $Y2=0
cc_431 CLK_N N_A_854_74#_c_1219_n 2.32931e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_432 N_CLK_N_M1024_g N_A_854_74#_M1028_g 0.039099f $X=4.72 $Y=2.235 $X2=0
+ $Y2=0
cc_433 N_CLK_N_c_532_n N_A_854_74#_c_1220_n 5.45517e-19 $X=4.645 $Y=1.385 $X2=0
+ $Y2=0
cc_434 N_CLK_N_c_530_n N_A_854_74#_c_1232_n 0.00265264f $X=4.195 $Y=1.22 $X2=0
+ $Y2=0
cc_435 N_CLK_N_c_532_n N_A_854_74#_c_1232_n 0.00755098f $X=4.645 $Y=1.385 $X2=0
+ $Y2=0
cc_436 CLK_N N_A_854_74#_c_1232_n 0.0287856f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_437 N_CLK_N_M1024_g N_A_854_74#_c_1257_n 0.00819326f $X=4.72 $Y=2.235 $X2=0
+ $Y2=0
cc_438 N_CLK_N_c_531_n N_A_854_74#_c_1246_n 0.0082943f $X=4.27 $Y=1.385 $X2=0
+ $Y2=0
cc_439 CLK_N N_A_854_74#_c_1246_n 0.0118859f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_440 N_CLK_N_M1024_g N_A_854_74#_c_1233_n 0.00366752f $X=4.72 $Y=2.235 $X2=0
+ $Y2=0
cc_441 N_CLK_N_c_530_n N_A_854_74#_c_1234_n 0.00336749f $X=4.195 $Y=1.22 $X2=0
+ $Y2=0
cc_442 N_CLK_N_c_532_n N_A_854_74#_c_1234_n 0.00366752f $X=4.645 $Y=1.385 $X2=0
+ $Y2=0
cc_443 CLK_N N_A_854_74#_c_1234_n 0.0276846f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_444 N_CLK_N_M1024_g N_VPWR_c_1723_n 0.0174456f $X=4.72 $Y=2.235 $X2=0 $Y2=0
cc_445 N_CLK_N_M1024_g N_VPWR_c_1721_n 8.51577e-19 $X=4.72 $Y=2.235 $X2=0 $Y2=0
cc_446 N_CLK_N_c_530_n N_A_284_464#_c_1864_n 0.00498249f $X=4.195 $Y=1.22 $X2=0
+ $Y2=0
cc_447 N_CLK_N_M1024_g N_A_284_464#_c_1864_n 0.00652376f $X=4.72 $Y=2.235 $X2=0
+ $Y2=0
cc_448 CLK_N N_A_284_464#_c_1864_n 0.0229434f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_449 N_CLK_N_c_530_n N_A_284_464#_c_1865_n 0.0173623f $X=4.195 $Y=1.22 $X2=0
+ $Y2=0
cc_450 N_CLK_N_M1024_g N_A_284_464#_c_1873_n 0.012568f $X=4.72 $Y=2.235 $X2=0
+ $Y2=0
cc_451 N_CLK_N_c_531_n N_A_284_464#_c_1873_n 0.00390191f $X=4.27 $Y=1.385 $X2=0
+ $Y2=0
cc_452 N_CLK_N_M1024_g N_A_284_464#_c_1874_n 0.0069622f $X=4.72 $Y=2.235 $X2=0
+ $Y2=0
cc_453 N_CLK_N_c_530_n N_A_284_464#_c_1867_n 0.00342374f $X=4.195 $Y=1.22 $X2=0
+ $Y2=0
cc_454 N_CLK_N_c_530_n N_VGND_c_2041_n 0.00314375f $X=4.195 $Y=1.22 $X2=0 $Y2=0
cc_455 N_CLK_N_c_530_n N_VGND_c_2046_n 0.00398514f $X=4.195 $Y=1.22 $X2=0 $Y2=0
cc_456 N_CLK_N_c_530_n N_VGND_c_2049_n 0.00428186f $X=4.195 $Y=1.22 $X2=0 $Y2=0
cc_457 N_CLK_N_c_530_n N_VGND_c_2050_n 0.00302001f $X=4.195 $Y=1.22 $X2=0 $Y2=0
cc_458 N_A_1049_347#_c_579_n N_A_1402_308#_M1036_d 0.0101435f $X=9.495 $Y=0.875
+ $X2=-0.19 $Y2=-0.245
cc_459 N_A_1049_347#_M1018_g N_A_1402_308#_M1025_g 0.0310025f $X=6.63 $Y=2.525
+ $X2=0 $Y2=0
cc_460 N_A_1049_347#_c_577_n N_A_1402_308#_M1029_g 0.00754889f $X=7.495 $Y=0.4
+ $X2=0 $Y2=0
cc_461 N_A_1049_347#_c_578_n N_A_1402_308#_M1029_g 0.00234219f $X=7.607 $Y=0.79
+ $X2=0 $Y2=0
cc_462 N_A_1049_347#_c_577_n N_A_1402_308#_c_754_n 6.3199e-19 $X=7.495 $Y=0.4
+ $X2=0 $Y2=0
cc_463 N_A_1049_347#_c_579_n N_A_1402_308#_c_754_n 0.0585797f $X=9.495 $Y=0.875
+ $X2=0 $Y2=0
cc_464 N_A_1049_347#_c_599_p N_A_1402_308#_c_754_n 0.0155432f $X=7.72 $Y=0.875
+ $X2=0 $Y2=0
cc_465 N_A_1049_347#_c_577_n N_A_1402_308#_c_755_n 0.00796913f $X=7.495 $Y=0.4
+ $X2=0 $Y2=0
cc_466 N_A_1049_347#_c_570_n N_A_1402_308#_c_771_n 3.25791e-19 $X=9.62 $Y=1.795
+ $X2=0 $Y2=0
cc_467 N_A_1049_347#_c_579_n N_A_1402_308#_c_771_n 0.0205002f $X=9.495 $Y=0.875
+ $X2=0 $Y2=0
cc_468 N_A_1049_347#_c_585_n N_A_1402_308#_c_771_n 0.00237334f $X=9.66 $Y=0.875
+ $X2=0 $Y2=0
cc_469 N_A_1049_347#_c_586_n N_A_1402_308#_c_771_n 3.9309e-19 $X=9.66 $Y=0.94
+ $X2=0 $Y2=0
cc_470 N_A_1049_347#_c_589_n N_A_1402_308#_c_760_n 0.00894366f $X=9.62 $Y=1.885
+ $X2=0 $Y2=0
cc_471 N_A_1049_347#_c_589_n N_A_1402_308#_c_776_n 0.00208707f $X=9.62 $Y=1.885
+ $X2=0 $Y2=0
cc_472 N_A_1049_347#_c_570_n N_A_1402_308#_c_756_n 0.00177595f $X=9.62 $Y=1.795
+ $X2=0 $Y2=0
cc_473 N_A_1049_347#_c_589_n N_A_1402_308#_c_756_n 6.95486e-19 $X=9.62 $Y=1.885
+ $X2=0 $Y2=0
cc_474 N_A_1049_347#_c_609_p N_A_1402_308#_c_757_n 2.86365e-19 $X=6.63 $Y=1.9
+ $X2=0 $Y2=0
cc_475 N_A_1049_347#_c_583_n N_A_1402_308#_c_757_n 0.019749f $X=6.63 $Y=1.9
+ $X2=0 $Y2=0
cc_476 N_A_1049_347#_M1018_g N_RESET_B_c_865_n 0.0100627f $X=6.63 $Y=2.525 $X2=0
+ $Y2=0
cc_477 N_A_1049_347#_c_577_n N_RESET_B_M1011_g 0.00162035f $X=7.495 $Y=0.4 $X2=0
+ $Y2=0
cc_478 N_A_1049_347#_c_578_n N_RESET_B_M1011_g 0.00611692f $X=7.607 $Y=0.79
+ $X2=0 $Y2=0
cc_479 N_A_1049_347#_c_579_n N_RESET_B_M1011_g 0.00712239f $X=9.495 $Y=0.875
+ $X2=0 $Y2=0
cc_480 N_A_1049_347#_c_599_p N_RESET_B_M1011_g 0.00232086f $X=7.72 $Y=0.875
+ $X2=0 $Y2=0
cc_481 N_A_1049_347#_M1028_d N_RESET_B_c_853_n 0.00128576f $X=5.245 $Y=1.735
+ $X2=0 $Y2=0
cc_482 N_A_1049_347#_c_574_n N_RESET_B_c_853_n 0.0311989f $X=5.55 $Y=1.735 $X2=0
+ $Y2=0
cc_483 N_A_1049_347#_c_575_n N_RESET_B_c_853_n 0.022138f $X=6.325 $Y=1.365 $X2=0
+ $Y2=0
cc_484 N_A_1049_347#_c_580_n N_RESET_B_c_853_n 0.0025432f $X=5.51 $Y=0.99 $X2=0
+ $Y2=0
cc_485 N_A_1049_347#_c_583_n N_RESET_B_c_853_n 0.00493928f $X=6.63 $Y=1.9 $X2=0
+ $Y2=0
cc_486 N_A_1049_347#_c_584_n N_RESET_B_c_853_n 0.0367773f $X=6.495 $Y=1.9 $X2=0
+ $Y2=0
cc_487 N_A_1049_347#_c_570_n N_RESET_B_c_855_n 0.0101256f $X=9.62 $Y=1.795 $X2=0
+ $Y2=0
cc_488 N_A_1049_347#_c_576_n N_A_1251_463#_M1023_d 0.00440809f $X=6.41 $Y=1.265
+ $X2=-0.19 $Y2=-0.245
cc_489 N_A_1049_347#_c_578_n N_A_1251_463#_c_1091_n 7.87457e-19 $X=7.607 $Y=0.79
+ $X2=0 $Y2=0
cc_490 N_A_1049_347#_c_579_n N_A_1251_463#_c_1091_n 0.0116106f $X=9.495 $Y=0.875
+ $X2=0 $Y2=0
cc_491 N_A_1049_347#_M1018_g N_A_1251_463#_c_1097_n 0.00561939f $X=6.63 $Y=2.525
+ $X2=0 $Y2=0
cc_492 N_A_1049_347#_M1018_g N_A_1251_463#_c_1098_n 0.00894477f $X=6.63 $Y=2.525
+ $X2=0 $Y2=0
cc_493 N_A_1049_347#_c_609_p N_A_1251_463#_c_1098_n 0.0101611f $X=6.63 $Y=1.9
+ $X2=0 $Y2=0
cc_494 N_A_1049_347#_c_583_n N_A_1251_463#_c_1098_n 0.00329986f $X=6.63 $Y=1.9
+ $X2=0 $Y2=0
cc_495 N_A_1049_347#_M1018_g N_A_1251_463#_c_1099_n 0.00167907f $X=6.63 $Y=2.525
+ $X2=0 $Y2=0
cc_496 N_A_1049_347#_c_609_p N_A_1251_463#_c_1099_n 0.00587482f $X=6.63 $Y=1.9
+ $X2=0 $Y2=0
cc_497 N_A_1049_347#_c_583_n N_A_1251_463#_c_1099_n 0.00210819f $X=6.63 $Y=1.9
+ $X2=0 $Y2=0
cc_498 N_A_1049_347#_c_584_n N_A_1251_463#_c_1099_n 0.0124877f $X=6.495 $Y=1.9
+ $X2=0 $Y2=0
cc_499 N_A_1049_347#_c_575_n N_A_1251_463#_c_1092_n 0.00890944f $X=6.325
+ $Y=1.365 $X2=0 $Y2=0
cc_500 N_A_1049_347#_c_576_n N_A_1251_463#_c_1092_n 0.00673678f $X=6.41 $Y=1.265
+ $X2=0 $Y2=0
cc_501 N_A_1049_347#_c_609_p N_A_1251_463#_c_1092_n 0.0256803f $X=6.63 $Y=1.9
+ $X2=0 $Y2=0
cc_502 N_A_1049_347#_c_583_n N_A_1251_463#_c_1092_n 0.00209786f $X=6.63 $Y=1.9
+ $X2=0 $Y2=0
cc_503 N_A_1049_347#_c_579_n N_A_1251_463#_c_1094_n 5.01488e-19 $X=9.495
+ $Y=0.875 $X2=0 $Y2=0
cc_504 N_A_1049_347#_c_569_n N_A_1251_463#_c_1095_n 0.00114937f $X=6.285
+ $Y=0.505 $X2=0 $Y2=0
cc_505 N_A_1049_347#_c_576_n N_A_1251_463#_c_1095_n 0.028804f $X=6.41 $Y=1.265
+ $X2=0 $Y2=0
cc_506 N_A_1049_347#_c_577_n N_A_1251_463#_c_1095_n 0.0261693f $X=7.495 $Y=0.4
+ $X2=0 $Y2=0
cc_507 N_A_1049_347#_c_609_p N_A_1251_463#_c_1095_n 6.22678e-19 $X=6.63 $Y=1.9
+ $X2=0 $Y2=0
cc_508 N_A_1049_347#_M1018_g N_A_1251_463#_c_1106_n 0.003748f $X=6.63 $Y=2.525
+ $X2=0 $Y2=0
cc_509 N_A_1049_347#_c_574_n N_A_854_74#_c_1219_n 0.00722098f $X=5.55 $Y=1.735
+ $X2=0 $Y2=0
cc_510 N_A_1049_347#_c_581_n N_A_854_74#_c_1219_n 0.00300836f $X=5.55 $Y=1.365
+ $X2=0 $Y2=0
cc_511 N_A_1049_347#_c_574_n N_A_854_74#_M1028_g 0.00495049f $X=5.55 $Y=1.735
+ $X2=0 $Y2=0
cc_512 N_A_1049_347#_c_573_n N_A_854_74#_c_1220_n 0.00308584f $X=5.55 $Y=1.265
+ $X2=0 $Y2=0
cc_513 N_A_1049_347#_c_580_n N_A_854_74#_c_1220_n 0.00315086f $X=5.51 $Y=0.99
+ $X2=0 $Y2=0
cc_514 N_A_1049_347#_c_574_n N_A_854_74#_c_1221_n 0.0104084f $X=5.55 $Y=1.735
+ $X2=0 $Y2=0
cc_515 N_A_1049_347#_c_575_n N_A_854_74#_c_1221_n 0.0143536f $X=6.325 $Y=1.365
+ $X2=0 $Y2=0
cc_516 N_A_1049_347#_c_581_n N_A_854_74#_c_1221_n 0.00821424f $X=5.55 $Y=1.365
+ $X2=0 $Y2=0
cc_517 N_A_1049_347#_c_584_n N_A_854_74#_c_1221_n 0.00839874f $X=6.495 $Y=1.9
+ $X2=0 $Y2=0
cc_518 N_A_1049_347#_M1018_g N_A_854_74#_M1004_g 0.0174741f $X=6.63 $Y=2.525
+ $X2=0 $Y2=0
cc_519 N_A_1049_347#_c_574_n N_A_854_74#_M1004_g 0.00434404f $X=5.55 $Y=1.735
+ $X2=0 $Y2=0
cc_520 N_A_1049_347#_c_609_p N_A_854_74#_M1004_g 4.61832e-19 $X=6.63 $Y=1.9
+ $X2=0 $Y2=0
cc_521 N_A_1049_347#_c_583_n N_A_854_74#_M1004_g 0.0213253f $X=6.63 $Y=1.9 $X2=0
+ $Y2=0
cc_522 N_A_1049_347#_c_584_n N_A_854_74#_M1004_g 0.0207517f $X=6.495 $Y=1.9
+ $X2=0 $Y2=0
cc_523 N_A_1049_347#_c_575_n N_A_854_74#_c_1223_n 0.00944798f $X=6.325 $Y=1.365
+ $X2=0 $Y2=0
cc_524 N_A_1049_347#_c_583_n N_A_854_74#_c_1223_n 0.019343f $X=6.63 $Y=1.9 $X2=0
+ $Y2=0
cc_525 N_A_1049_347#_c_584_n N_A_854_74#_c_1223_n 0.00488434f $X=6.495 $Y=1.9
+ $X2=0 $Y2=0
cc_526 N_A_1049_347#_c_583_n N_A_854_74#_c_1224_n 0.00129223f $X=6.63 $Y=1.9
+ $X2=0 $Y2=0
cc_527 N_A_1049_347#_c_569_n N_A_854_74#_M1014_g 0.00772147f $X=6.285 $Y=0.505
+ $X2=0 $Y2=0
cc_528 N_A_1049_347#_c_576_n N_A_854_74#_M1014_g 0.00376358f $X=6.41 $Y=1.265
+ $X2=0 $Y2=0
cc_529 N_A_1049_347#_c_577_n N_A_854_74#_M1014_g 0.014613f $X=7.495 $Y=0.4 $X2=0
+ $Y2=0
cc_530 N_A_1049_347#_c_577_n N_A_854_74#_c_1226_n 0.0169588f $X=7.495 $Y=0.4
+ $X2=0 $Y2=0
cc_531 N_A_1049_347#_c_579_n N_A_854_74#_c_1226_n 0.012696f $X=9.495 $Y=0.875
+ $X2=0 $Y2=0
cc_532 N_A_1049_347#_c_577_n N_A_854_74#_c_1227_n 0.00169598f $X=7.495 $Y=0.4
+ $X2=0 $Y2=0
cc_533 N_A_1049_347#_c_582_n N_A_854_74#_c_1227_n 0.0184785f $X=6.49 $Y=0.34
+ $X2=0 $Y2=0
cc_534 N_A_1049_347#_c_570_n N_A_854_74#_M1038_g 0.0072592f $X=9.62 $Y=1.795
+ $X2=0 $Y2=0
cc_535 N_A_1049_347#_c_579_n N_A_854_74#_M1038_g 0.0155998f $X=9.495 $Y=0.875
+ $X2=0 $Y2=0
cc_536 N_A_1049_347#_c_585_n N_A_854_74#_M1038_g 0.00155872f $X=9.66 $Y=0.875
+ $X2=0 $Y2=0
cc_537 N_A_1049_347#_c_586_n N_A_854_74#_M1038_g 0.0127811f $X=9.66 $Y=0.94
+ $X2=0 $Y2=0
cc_538 N_A_1049_347#_c_589_n N_A_854_74#_c_1229_n 0.022891f $X=9.62 $Y=1.885
+ $X2=0 $Y2=0
cc_539 N_A_1049_347#_c_589_n N_A_854_74#_c_1244_n 0.0107863f $X=9.62 $Y=1.885
+ $X2=0 $Y2=0
cc_540 N_A_1049_347#_c_569_n N_A_854_74#_c_1230_n 0.00978913f $X=6.285 $Y=0.505
+ $X2=0 $Y2=0
cc_541 N_A_1049_347#_c_575_n N_A_854_74#_c_1230_n 0.00545608f $X=6.325 $Y=1.365
+ $X2=0 $Y2=0
cc_542 N_A_1049_347#_c_569_n N_A_854_74#_c_1231_n 7.97985e-19 $X=6.285 $Y=0.505
+ $X2=0 $Y2=0
cc_543 N_A_1049_347#_c_575_n N_A_854_74#_c_1231_n 0.00297996f $X=6.325 $Y=1.365
+ $X2=0 $Y2=0
cc_544 N_A_1049_347#_c_576_n N_A_854_74#_c_1231_n 0.00299468f $X=6.41 $Y=1.265
+ $X2=0 $Y2=0
cc_545 N_A_1049_347#_c_577_n N_A_854_74#_c_1231_n 0.00142638f $X=7.495 $Y=0.4
+ $X2=0 $Y2=0
cc_546 N_A_1049_347#_c_582_n N_A_854_74#_c_1231_n 7.52532e-19 $X=6.49 $Y=0.34
+ $X2=0 $Y2=0
cc_547 N_A_1049_347#_c_609_p N_A_854_74#_c_1231_n 7.90828e-19 $X=6.63 $Y=1.9
+ $X2=0 $Y2=0
cc_548 N_A_1049_347#_c_574_n N_A_854_74#_c_1257_n 0.013092f $X=5.55 $Y=1.735
+ $X2=0 $Y2=0
cc_549 N_A_1049_347#_c_574_n N_A_854_74#_c_1245_n 0.00875048f $X=5.55 $Y=1.735
+ $X2=0 $Y2=0
cc_550 N_A_1049_347#_c_573_n N_A_854_74#_c_1233_n 0.0022818f $X=5.55 $Y=1.265
+ $X2=0 $Y2=0
cc_551 N_A_1049_347#_c_574_n N_A_854_74#_c_1233_n 0.0119751f $X=5.55 $Y=1.735
+ $X2=0 $Y2=0
cc_552 N_A_1049_347#_c_581_n N_A_854_74#_c_1233_n 0.0167142f $X=5.55 $Y=1.365
+ $X2=0 $Y2=0
cc_553 N_A_1049_347#_c_573_n N_A_854_74#_c_1234_n 0.005951f $X=5.55 $Y=1.265
+ $X2=0 $Y2=0
cc_554 N_A_1049_347#_c_570_n N_A_854_74#_c_1235_n 0.00379509f $X=9.62 $Y=1.795
+ $X2=0 $Y2=0
cc_555 N_A_1049_347#_c_579_n N_A_854_74#_c_1235_n 0.010781f $X=9.495 $Y=0.875
+ $X2=0 $Y2=0
cc_556 N_A_1049_347#_c_570_n N_A_854_74#_c_1236_n 0.0211113f $X=9.62 $Y=1.795
+ $X2=0 $Y2=0
cc_557 N_A_1049_347#_c_579_n N_A_854_74#_c_1236_n 6.48422e-19 $X=9.495 $Y=0.875
+ $X2=0 $Y2=0
cc_558 N_A_1049_347#_c_570_n N_A_854_74#_c_1237_n 8.24492e-19 $X=9.62 $Y=1.795
+ $X2=0 $Y2=0
cc_559 N_A_1049_347#_c_571_n N_A_854_74#_c_1237_n 3.59891e-19 $X=10.215 $Y=0.94
+ $X2=0 $Y2=0
cc_560 N_A_1049_347#_c_570_n N_A_854_74#_c_1238_n 0.0122344f $X=9.62 $Y=1.795
+ $X2=0 $Y2=0
cc_561 N_A_1049_347#_c_571_n N_A_854_74#_c_1238_n 0.0206875f $X=10.215 $Y=0.94
+ $X2=0 $Y2=0
cc_562 N_A_1049_347#_c_586_n N_A_854_74#_c_1238_n 3.57698e-19 $X=9.66 $Y=0.94
+ $X2=0 $Y2=0
cc_563 N_A_1049_347#_c_570_n N_A_854_74#_c_1239_n 0.0122704f $X=9.62 $Y=1.795
+ $X2=0 $Y2=0
cc_564 N_A_1049_347#_c_571_n N_A_854_74#_c_1239_n 0.00508082f $X=10.215 $Y=0.94
+ $X2=0 $Y2=0
cc_565 N_A_1049_347#_c_579_n N_A_854_74#_c_1239_n 0.00587076f $X=9.495 $Y=0.875
+ $X2=0 $Y2=0
cc_566 N_A_1049_347#_c_585_n N_A_854_74#_c_1239_n 0.023223f $X=9.66 $Y=0.875
+ $X2=0 $Y2=0
cc_567 N_A_1049_347#_c_586_n N_A_854_74#_c_1239_n 0.00358594f $X=9.66 $Y=0.94
+ $X2=0 $Y2=0
cc_568 N_A_1049_347#_c_572_n N_A_2087_410#_M1001_g 0.0383232f $X=10.29 $Y=0.865
+ $X2=0 $Y2=0
cc_569 N_A_1049_347#_c_579_n N_A_1827_144#_M1038_d 0.00486106f $X=9.495 $Y=0.875
+ $X2=-0.19 $Y2=-0.245
cc_570 N_A_1049_347#_c_585_n N_A_1827_144#_M1038_d 0.00351901f $X=9.66 $Y=0.875
+ $X2=-0.19 $Y2=-0.245
cc_571 N_A_1049_347#_c_589_n N_A_1827_144#_c_1536_n 0.00398969f $X=9.62 $Y=1.885
+ $X2=0 $Y2=0
cc_572 N_A_1049_347#_c_572_n N_A_1827_144#_c_1523_n 0.00722667f $X=10.29
+ $Y=0.865 $X2=0 $Y2=0
cc_573 N_A_1049_347#_c_571_n N_A_1827_144#_c_1524_n 0.00394505f $X=10.215
+ $Y=0.94 $X2=0 $Y2=0
cc_574 N_A_1049_347#_c_572_n N_A_1827_144#_c_1524_n 0.00616225f $X=10.29
+ $Y=0.865 $X2=0 $Y2=0
cc_575 N_A_1049_347#_c_585_n N_A_1827_144#_c_1524_n 0.0062694f $X=9.66 $Y=0.875
+ $X2=0 $Y2=0
cc_576 N_A_1049_347#_c_570_n N_A_1827_144#_c_1538_n 0.0038782f $X=9.62 $Y=1.795
+ $X2=0 $Y2=0
cc_577 N_A_1049_347#_c_571_n N_A_1827_144#_c_1525_n 0.0127777f $X=10.215 $Y=0.94
+ $X2=0 $Y2=0
cc_578 N_A_1049_347#_c_571_n N_A_1827_144#_c_1526_n 0.00537903f $X=10.215
+ $Y=0.94 $X2=0 $Y2=0
cc_579 N_A_1049_347#_c_585_n N_A_1827_144#_c_1526_n 0.0136829f $X=9.66 $Y=0.875
+ $X2=0 $Y2=0
cc_580 N_A_1049_347#_c_586_n N_A_1827_144#_c_1526_n 5.82391e-19 $X=9.66 $Y=0.94
+ $X2=0 $Y2=0
cc_581 N_A_1049_347#_c_579_n N_A_1827_144#_c_1529_n 0.0227442f $X=9.495 $Y=0.875
+ $X2=0 $Y2=0
cc_582 N_A_1049_347#_c_585_n N_A_1827_144#_c_1529_n 0.02606f $X=9.66 $Y=0.875
+ $X2=0 $Y2=0
cc_583 N_A_1049_347#_c_586_n N_A_1827_144#_c_1529_n 0.00780225f $X=9.66 $Y=0.94
+ $X2=0 $Y2=0
cc_584 N_A_1049_347#_c_589_n N_VPWR_c_1736_n 0.00439937f $X=9.62 $Y=1.885 $X2=0
+ $Y2=0
cc_585 N_A_1049_347#_M1018_g N_VPWR_c_1721_n 9.39239e-19 $X=6.63 $Y=2.525 $X2=0
+ $Y2=0
cc_586 N_A_1049_347#_c_589_n N_VPWR_c_1721_n 0.00845445f $X=9.62 $Y=1.885 $X2=0
+ $Y2=0
cc_587 N_A_1049_347#_M1010_d N_A_284_464#_c_1865_n 0.00672786f $X=5.37 $Y=0.395
+ $X2=0 $Y2=0
cc_588 N_A_1049_347#_c_569_n N_A_284_464#_c_1865_n 0.00300858f $X=6.285 $Y=0.505
+ $X2=0 $Y2=0
cc_589 N_A_1049_347#_c_575_n N_A_284_464#_c_1865_n 0.00758662f $X=6.325 $Y=1.365
+ $X2=0 $Y2=0
cc_590 N_A_1049_347#_c_725_p N_A_284_464#_c_1865_n 0.00133713f $X=6.41 $Y=0.545
+ $X2=0 $Y2=0
cc_591 N_A_1049_347#_c_576_n N_A_284_464#_c_1865_n 0.00846067f $X=6.41 $Y=1.265
+ $X2=0 $Y2=0
cc_592 N_A_1049_347#_c_580_n N_A_284_464#_c_1865_n 0.0217849f $X=5.51 $Y=0.99
+ $X2=0 $Y2=0
cc_593 N_A_1049_347#_M1028_d N_A_284_464#_c_1874_n 0.012782f $X=5.245 $Y=1.735
+ $X2=0 $Y2=0
cc_594 N_A_1049_347#_M1018_g N_A_284_464#_c_1874_n 4.15589e-19 $X=6.63 $Y=2.525
+ $X2=0 $Y2=0
cc_595 N_A_1049_347#_c_574_n N_A_284_464#_c_1874_n 0.0294456f $X=5.55 $Y=1.735
+ $X2=0 $Y2=0
cc_596 N_A_1049_347#_c_584_n N_A_284_464#_c_1874_n 0.0344103f $X=6.495 $Y=1.9
+ $X2=0 $Y2=0
cc_597 N_A_1049_347#_c_569_n N_A_284_464#_c_1866_n 0.00132847f $X=6.285 $Y=0.505
+ $X2=0 $Y2=0
cc_598 N_A_1049_347#_c_575_n N_A_284_464#_c_1866_n 0.0200739f $X=6.325 $Y=1.365
+ $X2=0 $Y2=0
cc_599 N_A_1049_347#_c_576_n N_A_284_464#_c_1866_n 0.0157403f $X=6.41 $Y=1.265
+ $X2=0 $Y2=0
cc_600 N_A_1049_347#_c_580_n N_A_284_464#_c_1866_n 0.0148107f $X=5.51 $Y=0.99
+ $X2=0 $Y2=0
cc_601 N_A_1049_347#_c_579_n N_VGND_M1011_d 0.00709166f $X=9.495 $Y=0.875 $X2=0
+ $Y2=0
cc_602 N_A_1049_347#_c_577_n N_VGND_c_2037_n 0.0252077f $X=7.495 $Y=0.4 $X2=0
+ $Y2=0
cc_603 N_A_1049_347#_c_578_n N_VGND_c_2037_n 0.00548912f $X=7.607 $Y=0.79 $X2=0
+ $Y2=0
cc_604 N_A_1049_347#_c_579_n N_VGND_c_2037_n 0.0259785f $X=9.495 $Y=0.875 $X2=0
+ $Y2=0
cc_605 N_A_1049_347#_c_572_n N_VGND_c_2038_n 0.00143784f $X=10.29 $Y=0.865 $X2=0
+ $Y2=0
cc_606 N_A_1049_347#_c_725_p N_VGND_c_2042_n 0.0115893f $X=6.41 $Y=0.545 $X2=0
+ $Y2=0
cc_607 N_A_1049_347#_c_577_n N_VGND_c_2042_n 0.079826f $X=7.495 $Y=0.4 $X2=0
+ $Y2=0
cc_608 N_A_1049_347#_c_582_n N_VGND_c_2042_n 0.0105761f $X=6.49 $Y=0.34 $X2=0
+ $Y2=0
cc_609 N_A_1049_347#_c_572_n N_VGND_c_2043_n 0.00461464f $X=10.29 $Y=0.865 $X2=0
+ $Y2=0
cc_610 N_A_1049_347#_c_572_n N_VGND_c_2046_n 0.00914127f $X=10.29 $Y=0.865 $X2=0
+ $Y2=0
cc_611 N_A_1049_347#_c_725_p N_VGND_c_2046_n 0.00583135f $X=6.41 $Y=0.545 $X2=0
+ $Y2=0
cc_612 N_A_1049_347#_c_577_n N_VGND_c_2046_n 0.0423052f $X=7.495 $Y=0.4 $X2=0
+ $Y2=0
cc_613 N_A_1049_347#_c_579_n N_VGND_c_2046_n 0.0372313f $X=9.495 $Y=0.875 $X2=0
+ $Y2=0
cc_614 N_A_1049_347#_c_582_n N_VGND_c_2046_n 0.0169086f $X=6.49 $Y=0.34 $X2=0
+ $Y2=0
cc_615 N_A_1049_347#_c_586_n N_VGND_c_2046_n 0.00102356f $X=9.66 $Y=0.94 $X2=0
+ $Y2=0
cc_616 N_A_1049_347#_c_599_p A_1489_123# 0.00142589f $X=7.72 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_617 N_A_1402_308#_M1025_g N_RESET_B_c_865_n 0.0103219f $X=7.085 $Y=2.525
+ $X2=0 $Y2=0
cc_618 N_A_1402_308#_M1029_g N_RESET_B_M1011_g 0.054628f $X=7.37 $Y=0.825 $X2=0
+ $Y2=0
cc_619 N_A_1402_308#_c_753_n N_RESET_B_M1011_g 0.00354335f $X=7.31 $Y=1.705
+ $X2=0 $Y2=0
cc_620 N_A_1402_308#_c_754_n N_RESET_B_M1011_g 0.0108751f $X=8.69 $Y=1.215 $X2=0
+ $Y2=0
cc_621 N_A_1402_308#_M1025_g N_RESET_B_c_869_n 0.0042902f $X=7.085 $Y=2.525
+ $X2=0 $Y2=0
cc_622 N_A_1402_308#_M1025_g N_RESET_B_c_872_n 0.0147496f $X=7.085 $Y=2.525
+ $X2=0 $Y2=0
cc_623 N_A_1402_308#_c_757_n N_RESET_B_c_872_n 9.81926e-19 $X=7.37 $Y=1.705
+ $X2=0 $Y2=0
cc_624 N_A_1402_308#_c_753_n N_RESET_B_c_853_n 0.0220824f $X=7.31 $Y=1.705 $X2=0
+ $Y2=0
cc_625 N_A_1402_308#_c_754_n N_RESET_B_c_853_n 0.00836974f $X=8.69 $Y=1.215
+ $X2=0 $Y2=0
cc_626 N_A_1402_308#_c_757_n N_RESET_B_c_853_n 0.00847455f $X=7.37 $Y=1.705
+ $X2=0 $Y2=0
cc_627 N_A_1402_308#_c_754_n N_RESET_B_c_855_n 0.0122156f $X=8.69 $Y=1.215 $X2=0
+ $Y2=0
cc_628 N_A_1402_308#_c_771_n N_RESET_B_c_855_n 0.0039881f $X=8.775 $Y=1.3 $X2=0
+ $Y2=0
cc_629 N_A_1402_308#_c_776_n N_RESET_B_c_855_n 0.0139612f $X=8.96 $Y=2.135 $X2=0
+ $Y2=0
cc_630 N_A_1402_308#_c_756_n N_RESET_B_c_855_n 0.0219481f $X=9.127 $Y=1.97 $X2=0
+ $Y2=0
cc_631 N_A_1402_308#_c_753_n N_RESET_B_c_856_n 5.09359e-19 $X=7.31 $Y=1.705
+ $X2=0 $Y2=0
cc_632 N_A_1402_308#_c_754_n N_RESET_B_c_856_n 0.00251018f $X=8.69 $Y=1.215
+ $X2=0 $Y2=0
cc_633 N_A_1402_308#_c_753_n N_RESET_B_c_860_n 0.00112909f $X=7.31 $Y=1.705
+ $X2=0 $Y2=0
cc_634 N_A_1402_308#_c_754_n N_RESET_B_c_860_n 0.0040357f $X=8.69 $Y=1.215 $X2=0
+ $Y2=0
cc_635 N_A_1402_308#_c_757_n N_RESET_B_c_860_n 0.021912f $X=7.37 $Y=1.705 $X2=0
+ $Y2=0
cc_636 N_A_1402_308#_c_753_n N_RESET_B_c_861_n 0.0187627f $X=7.31 $Y=1.705 $X2=0
+ $Y2=0
cc_637 N_A_1402_308#_c_754_n N_RESET_B_c_861_n 0.0238842f $X=8.69 $Y=1.215 $X2=0
+ $Y2=0
cc_638 N_A_1402_308#_c_757_n N_RESET_B_c_861_n 9.28438e-19 $X=7.37 $Y=1.705
+ $X2=0 $Y2=0
cc_639 N_A_1402_308#_c_754_n N_A_1251_463#_c_1091_n 0.0123021f $X=8.69 $Y=1.215
+ $X2=0 $Y2=0
cc_640 N_A_1402_308#_c_756_n N_A_1251_463#_c_1091_n 0.00380436f $X=9.127 $Y=1.97
+ $X2=0 $Y2=0
cc_641 N_A_1402_308#_c_760_n N_A_1251_463#_c_1096_n 0.0165257f $X=8.96 $Y=2.815
+ $X2=0 $Y2=0
cc_642 N_A_1402_308#_c_776_n N_A_1251_463#_c_1096_n 0.010014f $X=8.96 $Y=2.135
+ $X2=0 $Y2=0
cc_643 N_A_1402_308#_c_756_n N_A_1251_463#_c_1096_n 0.0028748f $X=9.127 $Y=1.97
+ $X2=0 $Y2=0
cc_644 N_A_1402_308#_M1025_g N_A_1251_463#_c_1097_n 8.84448e-19 $X=7.085
+ $Y=2.525 $X2=0 $Y2=0
cc_645 N_A_1402_308#_M1025_g N_A_1251_463#_c_1098_n 2.77965e-19 $X=7.085
+ $Y=2.525 $X2=0 $Y2=0
cc_646 N_A_1402_308#_M1025_g N_A_1251_463#_c_1092_n 0.00449197f $X=7.085
+ $Y=2.525 $X2=0 $Y2=0
cc_647 N_A_1402_308#_M1029_g N_A_1251_463#_c_1092_n 0.00123795f $X=7.37 $Y=0.825
+ $X2=0 $Y2=0
cc_648 N_A_1402_308#_c_753_n N_A_1251_463#_c_1092_n 0.0409458f $X=7.31 $Y=1.705
+ $X2=0 $Y2=0
cc_649 N_A_1402_308#_c_755_n N_A_1251_463#_c_1092_n 0.0136822f $X=7.475 $Y=1.215
+ $X2=0 $Y2=0
cc_650 N_A_1402_308#_c_757_n N_A_1251_463#_c_1092_n 0.0093719f $X=7.37 $Y=1.705
+ $X2=0 $Y2=0
cc_651 N_A_1402_308#_M1025_g N_A_1251_463#_c_1101_n 0.0107384f $X=7.085 $Y=2.525
+ $X2=0 $Y2=0
cc_652 N_A_1402_308#_c_753_n N_A_1251_463#_c_1101_n 0.0185663f $X=7.31 $Y=1.705
+ $X2=0 $Y2=0
cc_653 N_A_1402_308#_c_757_n N_A_1251_463#_c_1101_n 0.00415575f $X=7.37 $Y=1.705
+ $X2=0 $Y2=0
cc_654 N_A_1402_308#_M1025_g N_A_1251_463#_c_1102_n 5.45053e-19 $X=7.085
+ $Y=2.525 $X2=0 $Y2=0
cc_655 N_A_1402_308#_c_754_n N_A_1251_463#_c_1103_n 0.00193481f $X=8.69 $Y=1.215
+ $X2=0 $Y2=0
cc_656 N_A_1402_308#_c_776_n N_A_1251_463#_c_1103_n 0.0147905f $X=8.96 $Y=2.135
+ $X2=0 $Y2=0
cc_657 N_A_1402_308#_c_754_n N_A_1251_463#_c_1093_n 0.0178831f $X=8.69 $Y=1.215
+ $X2=0 $Y2=0
cc_658 N_A_1402_308#_c_756_n N_A_1251_463#_c_1093_n 0.0355404f $X=9.127 $Y=1.97
+ $X2=0 $Y2=0
cc_659 N_A_1402_308#_c_754_n N_A_1251_463#_c_1094_n 0.00727625f $X=8.69 $Y=1.215
+ $X2=0 $Y2=0
cc_660 N_A_1402_308#_c_756_n N_A_1251_463#_c_1094_n 0.0121655f $X=9.127 $Y=1.97
+ $X2=0 $Y2=0
cc_661 N_A_1402_308#_M1029_g N_A_1251_463#_c_1095_n 0.0017182f $X=7.37 $Y=0.825
+ $X2=0 $Y2=0
cc_662 N_A_1402_308#_M1025_g N_A_1251_463#_c_1106_n 0.00906899f $X=7.085
+ $Y=2.525 $X2=0 $Y2=0
cc_663 N_A_1402_308#_M1025_g N_A_1251_463#_c_1107_n 5.94501e-19 $X=7.085
+ $Y=2.525 $X2=0 $Y2=0
cc_664 N_A_1402_308#_c_754_n N_A_1251_463#_c_1107_n 4.94171e-19 $X=8.69 $Y=1.215
+ $X2=0 $Y2=0
cc_665 N_A_1402_308#_c_757_n N_A_854_74#_c_1224_n 0.00251163f $X=7.37 $Y=1.705
+ $X2=0 $Y2=0
cc_666 N_A_1402_308#_M1029_g N_A_854_74#_M1014_g 0.0424842f $X=7.37 $Y=0.825
+ $X2=0 $Y2=0
cc_667 N_A_1402_308#_c_755_n N_A_854_74#_M1014_g 0.001136f $X=7.475 $Y=1.215
+ $X2=0 $Y2=0
cc_668 N_A_1402_308#_M1029_g N_A_854_74#_c_1226_n 0.00973286f $X=7.37 $Y=0.825
+ $X2=0 $Y2=0
cc_669 N_A_1402_308#_c_771_n N_A_854_74#_M1038_g 0.00746547f $X=8.775 $Y=1.3
+ $X2=0 $Y2=0
cc_670 N_A_1402_308#_c_756_n N_A_854_74#_M1038_g 0.00329096f $X=9.127 $Y=1.97
+ $X2=0 $Y2=0
cc_671 N_A_1402_308#_c_760_n N_A_854_74#_c_1244_n 3.62308e-19 $X=8.96 $Y=2.815
+ $X2=0 $Y2=0
cc_672 N_A_1402_308#_M1029_g N_A_854_74#_c_1231_n 0.00354086f $X=7.37 $Y=0.825
+ $X2=0 $Y2=0
cc_673 N_A_1402_308#_c_776_n N_A_854_74#_c_1235_n 0.0246346f $X=8.96 $Y=2.135
+ $X2=0 $Y2=0
cc_674 N_A_1402_308#_c_756_n N_A_854_74#_c_1235_n 0.0296228f $X=9.127 $Y=1.97
+ $X2=0 $Y2=0
cc_675 N_A_1402_308#_c_776_n N_A_854_74#_c_1236_n 0.00410579f $X=8.96 $Y=2.135
+ $X2=0 $Y2=0
cc_676 N_A_1402_308#_c_776_n N_A_854_74#_c_1239_n 0.00363905f $X=8.96 $Y=2.135
+ $X2=0 $Y2=0
cc_677 N_A_1402_308#_c_776_n N_A_1827_144#_c_1536_n 0.0430929f $X=8.96 $Y=2.135
+ $X2=0 $Y2=0
cc_678 N_A_1402_308#_M1025_g N_VPWR_c_1724_n 0.00574172f $X=7.085 $Y=2.525 $X2=0
+ $Y2=0
cc_679 N_A_1402_308#_c_760_n N_VPWR_c_1725_n 0.0260221f $X=8.96 $Y=2.815 $X2=0
+ $Y2=0
cc_680 N_A_1402_308#_c_760_n N_VPWR_c_1736_n 0.0342121f $X=8.96 $Y=2.815 $X2=0
+ $Y2=0
cc_681 N_A_1402_308#_M1025_g N_VPWR_c_1721_n 9.39239e-19 $X=7.085 $Y=2.525 $X2=0
+ $Y2=0
cc_682 N_A_1402_308#_c_760_n N_VPWR_c_1721_n 0.0282732f $X=8.96 $Y=2.815 $X2=0
+ $Y2=0
cc_683 N_A_1402_308#_c_754_n N_VGND_M1011_d 0.00610455f $X=8.69 $Y=1.215 $X2=0
+ $Y2=0
cc_684 N_RESET_B_M1011_g N_A_1251_463#_c_1091_n 0.0249736f $X=7.76 $Y=0.825
+ $X2=0 $Y2=0
cc_685 N_RESET_B_c_865_n N_A_1251_463#_c_1097_n 0.00484256f $X=7.46 $Y=3.15
+ $X2=0 $Y2=0
cc_686 N_RESET_B_c_865_n N_A_1251_463#_c_1098_n 0.00368249f $X=7.46 $Y=3.15
+ $X2=0 $Y2=0
cc_687 N_RESET_B_c_853_n N_A_1251_463#_c_1098_n 0.005679f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_688 N_RESET_B_c_869_n N_A_1251_463#_c_1092_n 5.45076e-19 $X=7.76 $Y=2.08
+ $X2=0 $Y2=0
cc_689 N_RESET_B_c_853_n N_A_1251_463#_c_1092_n 0.0207084f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_690 N_RESET_B_c_872_n N_A_1251_463#_c_1101_n 0.00953823f $X=7.76 $Y=2.16
+ $X2=0 $Y2=0
cc_691 N_RESET_B_c_853_n N_A_1251_463#_c_1101_n 0.011158f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_692 N_RESET_B_M1013_g N_A_1251_463#_c_1102_n 0.00933053f $X=7.535 $Y=2.525
+ $X2=0 $Y2=0
cc_693 N_RESET_B_c_872_n N_A_1251_463#_c_1102_n 0.00667846f $X=7.76 $Y=2.16
+ $X2=0 $Y2=0
cc_694 N_RESET_B_c_855_n N_A_1251_463#_c_1103_n 0.00467221f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_695 N_RESET_B_c_856_n N_A_1251_463#_c_1103_n 0.00160883f $X=8.065 $Y=1.665
+ $X2=0 $Y2=0
cc_696 N_RESET_B_c_860_n N_A_1251_463#_c_1103_n 0.00145514f $X=7.85 $Y=1.635
+ $X2=0 $Y2=0
cc_697 N_RESET_B_c_861_n N_A_1251_463#_c_1103_n 0.00585893f $X=7.85 $Y=1.635
+ $X2=0 $Y2=0
cc_698 N_RESET_B_c_869_n N_A_1251_463#_c_1093_n 0.00489681f $X=7.76 $Y=2.08
+ $X2=0 $Y2=0
cc_699 N_RESET_B_c_855_n N_A_1251_463#_c_1093_n 0.0187239f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_700 N_RESET_B_c_856_n N_A_1251_463#_c_1093_n 0.00261643f $X=8.065 $Y=1.665
+ $X2=0 $Y2=0
cc_701 N_RESET_B_c_860_n N_A_1251_463#_c_1093_n 4.84312e-19 $X=7.85 $Y=1.635
+ $X2=0 $Y2=0
cc_702 N_RESET_B_c_861_n N_A_1251_463#_c_1093_n 0.0210281f $X=7.85 $Y=1.635
+ $X2=0 $Y2=0
cc_703 N_RESET_B_c_855_n N_A_1251_463#_c_1094_n 0.00633088f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_704 N_RESET_B_c_856_n N_A_1251_463#_c_1094_n 0.00141062f $X=8.065 $Y=1.665
+ $X2=0 $Y2=0
cc_705 N_RESET_B_c_860_n N_A_1251_463#_c_1094_n 0.0219831f $X=7.85 $Y=1.635
+ $X2=0 $Y2=0
cc_706 N_RESET_B_c_861_n N_A_1251_463#_c_1094_n 0.00167181f $X=7.85 $Y=1.635
+ $X2=0 $Y2=0
cc_707 N_RESET_B_c_853_n N_A_1251_463#_c_1095_n 0.00764587f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_708 N_RESET_B_c_865_n N_A_1251_463#_c_1106_n 0.00243913f $X=7.46 $Y=3.15
+ $X2=0 $Y2=0
cc_709 N_RESET_B_c_872_n N_A_1251_463#_c_1106_n 5.5457e-19 $X=7.76 $Y=2.16 $X2=0
+ $Y2=0
cc_710 N_RESET_B_c_869_n N_A_1251_463#_c_1107_n 0.00755054f $X=7.76 $Y=2.08
+ $X2=0 $Y2=0
cc_711 N_RESET_B_c_872_n N_A_1251_463#_c_1107_n 0.00746081f $X=7.76 $Y=2.16
+ $X2=0 $Y2=0
cc_712 N_RESET_B_c_853_n N_A_1251_463#_c_1107_n 0.00513269f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_713 N_RESET_B_c_856_n N_A_1251_463#_c_1107_n 0.00138918f $X=8.065 $Y=1.665
+ $X2=0 $Y2=0
cc_714 N_RESET_B_c_860_n N_A_1251_463#_c_1107_n 0.002679f $X=7.85 $Y=1.635 $X2=0
+ $Y2=0
cc_715 N_RESET_B_c_861_n N_A_1251_463#_c_1107_n 0.0196346f $X=7.85 $Y=1.635
+ $X2=0 $Y2=0
cc_716 N_RESET_B_c_853_n N_A_854_74#_M1024_s 0.00245167f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_717 N_RESET_B_c_853_n N_A_854_74#_c_1219_n 0.0148135f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_718 N_RESET_B_c_865_n N_A_854_74#_M1028_g 0.0103562f $X=7.46 $Y=3.15 $X2=0
+ $Y2=0
cc_719 N_RESET_B_c_853_n N_A_854_74#_M1028_g 0.00487748f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_720 N_RESET_B_c_865_n N_A_854_74#_M1004_g 0.0103747f $X=7.46 $Y=3.15 $X2=0
+ $Y2=0
cc_721 N_RESET_B_c_853_n N_A_854_74#_M1004_g 0.00780418f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_722 N_RESET_B_c_853_n N_A_854_74#_c_1223_n 0.00861652f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_723 N_RESET_B_c_853_n N_A_854_74#_c_1224_n 0.00234989f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_724 N_RESET_B_M1011_g N_A_854_74#_c_1226_n 0.00994376f $X=7.76 $Y=0.825 $X2=0
+ $Y2=0
cc_725 N_RESET_B_c_855_n N_A_854_74#_c_1229_n 0.00323464f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_726 N_RESET_B_c_853_n N_A_854_74#_c_1232_n 0.00637363f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_727 N_RESET_B_c_853_n N_A_854_74#_c_1245_n 0.0123343f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_728 N_RESET_B_c_853_n N_A_854_74#_c_1246_n 0.0201134f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_729 N_RESET_B_c_853_n N_A_854_74#_c_1233_n 0.0223879f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_730 N_RESET_B_c_855_n N_A_854_74#_c_1235_n 0.0288686f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_731 N_RESET_B_c_855_n N_A_854_74#_c_1236_n 0.00214944f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_732 N_RESET_B_c_863_n N_A_854_74#_c_1237_n 0.00866981f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_733 N_RESET_B_c_855_n N_A_854_74#_c_1238_n 0.00443162f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_734 N_RESET_B_c_855_n N_A_854_74#_c_1239_n 0.0328537f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_735 N_RESET_B_c_871_n N_A_2087_410#_c_1429_n 0.00937683f $X=11.32 $Y=2.465
+ $X2=0 $Y2=0
cc_736 N_RESET_B_c_873_n N_A_2087_410#_c_1429_n 0.0129752f $X=11.25 $Y=2.375
+ $X2=0 $Y2=0
cc_737 N_RESET_B_M1007_g N_A_2087_410#_M1001_g 0.0291977f $X=11.25 $Y=0.58 $X2=0
+ $Y2=0
cc_738 N_RESET_B_c_852_n N_A_2087_410#_M1001_g 0.0115721f $X=11.25 $Y=2.285
+ $X2=0 $Y2=0
cc_739 N_RESET_B_c_855_n N_A_2087_410#_M1001_g 0.00415382f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_740 N_RESET_B_c_857_n N_A_2087_410#_M1001_g 6.26309e-19 $X=11.28 $Y=1.665
+ $X2=0 $Y2=0
cc_741 N_RESET_B_c_862_n N_A_2087_410#_M1001_g 0.0175496f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_742 N_RESET_B_c_863_n N_A_2087_410#_M1001_g 0.00267234f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_743 N_RESET_B_c_873_n N_A_2087_410#_c_1431_n 0.015263f $X=11.25 $Y=2.375
+ $X2=0 $Y2=0
cc_744 N_RESET_B_c_855_n N_A_2087_410#_c_1431_n 0.00166773f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_745 N_RESET_B_c_871_n N_A_2087_410#_c_1432_n 0.0127946f $X=11.32 $Y=2.465
+ $X2=0 $Y2=0
cc_746 N_RESET_B_c_873_n N_A_2087_410#_c_1432_n 3.39749e-19 $X=11.25 $Y=2.375
+ $X2=0 $Y2=0
cc_747 N_RESET_B_M1007_g N_A_2087_410#_c_1427_n 7.40512e-19 $X=11.25 $Y=0.58
+ $X2=0 $Y2=0
cc_748 N_RESET_B_c_852_n N_A_2087_410#_c_1435_n 8.51156e-19 $X=11.25 $Y=2.285
+ $X2=0 $Y2=0
cc_749 N_RESET_B_c_855_n N_A_2087_410#_c_1435_n 0.00135183f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_750 N_RESET_B_c_873_n N_A_2087_410#_c_1436_n 0.00255599f $X=11.25 $Y=2.375
+ $X2=0 $Y2=0
cc_751 N_RESET_B_M1007_g N_A_1827_144#_c_1517_n 0.0238259f $X=11.25 $Y=0.58
+ $X2=0 $Y2=0
cc_752 N_RESET_B_c_852_n N_A_1827_144#_c_1518_n 0.0238259f $X=11.25 $Y=2.285
+ $X2=0 $Y2=0
cc_753 N_RESET_B_c_863_n N_A_1827_144#_c_1518_n 0.00218879f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_754 N_RESET_B_c_852_n N_A_1827_144#_c_1519_n 0.0243914f $X=11.25 $Y=2.285
+ $X2=0 $Y2=0
cc_755 N_RESET_B_c_863_n N_A_1827_144#_c_1519_n 4.39803e-19 $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_756 N_RESET_B_c_873_n N_A_1827_144#_c_1531_n 0.00851518f $X=11.25 $Y=2.375
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_871_n N_A_1827_144#_c_1532_n 0.00937083f $X=11.32 $Y=2.465
+ $X2=0 $Y2=0
cc_758 N_RESET_B_c_857_n N_A_1827_144#_c_1522_n 3.16322e-19 $X=11.28 $Y=1.665
+ $X2=0 $Y2=0
cc_759 N_RESET_B_c_855_n N_A_1827_144#_c_1537_n 0.0335459f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_760 N_RESET_B_c_855_n N_A_1827_144#_c_1538_n 0.0208272f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_761 N_RESET_B_M1007_g N_A_1827_144#_c_1525_n 0.0143997f $X=11.25 $Y=0.58
+ $X2=0 $Y2=0
cc_762 N_RESET_B_c_855_n N_A_1827_144#_c_1525_n 0.0122847f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_763 N_RESET_B_c_857_n N_A_1827_144#_c_1525_n 0.00174298f $X=11.28 $Y=1.665
+ $X2=0 $Y2=0
cc_764 N_RESET_B_c_862_n N_A_1827_144#_c_1525_n 0.00126891f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_765 N_RESET_B_c_863_n N_A_1827_144#_c_1525_n 0.0296916f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_766 N_RESET_B_c_852_n N_A_1827_144#_c_1539_n 0.0105998f $X=11.25 $Y=2.285
+ $X2=0 $Y2=0
cc_767 N_RESET_B_c_873_n N_A_1827_144#_c_1539_n 0.00215447f $X=11.25 $Y=2.375
+ $X2=0 $Y2=0
cc_768 N_RESET_B_c_855_n N_A_1827_144#_c_1539_n 0.00297115f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_769 N_RESET_B_c_857_n N_A_1827_144#_c_1539_n 0.00466048f $X=11.28 $Y=1.665
+ $X2=0 $Y2=0
cc_770 N_RESET_B_c_862_n N_A_1827_144#_c_1539_n 8.68178e-19 $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_771 N_RESET_B_c_863_n N_A_1827_144#_c_1539_n 0.0158387f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_772 N_RESET_B_M1007_g N_A_1827_144#_c_1527_n 0.00109112f $X=11.25 $Y=0.58
+ $X2=0 $Y2=0
cc_773 N_RESET_B_c_852_n N_A_1827_144#_c_1527_n 0.00231391f $X=11.25 $Y=2.285
+ $X2=0 $Y2=0
cc_774 N_RESET_B_c_857_n N_A_1827_144#_c_1527_n 0.00755838f $X=11.28 $Y=1.665
+ $X2=0 $Y2=0
cc_775 N_RESET_B_c_862_n N_A_1827_144#_c_1527_n 3.9684e-19 $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_776 N_RESET_B_c_863_n N_A_1827_144#_c_1527_n 0.0432263f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_777 N_RESET_B_c_862_n N_A_1827_144#_c_1528_n 0.0238259f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_778 N_RESET_B_c_852_n N_A_1827_144#_c_1541_n 0.00258184f $X=11.25 $Y=2.285
+ $X2=0 $Y2=0
cc_779 N_RESET_B_c_855_n N_A_1827_144#_c_1541_n 0.00615148f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_780 N_RESET_B_c_857_n N_A_1827_144#_c_1541_n 0.00137624f $X=11.28 $Y=1.665
+ $X2=0 $Y2=0
cc_781 N_RESET_B_c_863_n N_A_1827_144#_c_1541_n 0.00644897f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_782 N_RESET_B_c_853_n N_VPWR_M1024_d 0.00107109f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_783 N_RESET_B_c_865_n N_VPWR_c_1723_n 0.0254401f $X=7.46 $Y=3.15 $X2=0 $Y2=0
cc_784 N_RESET_B_c_865_n N_VPWR_c_1724_n 0.0159389f $X=7.46 $Y=3.15 $X2=0 $Y2=0
cc_785 N_RESET_B_M1013_g N_VPWR_c_1724_n 0.0121568f $X=7.535 $Y=2.525 $X2=0
+ $Y2=0
cc_786 N_RESET_B_M1013_g N_VPWR_c_1725_n 0.0103331f $X=7.535 $Y=2.525 $X2=0
+ $Y2=0
cc_787 N_RESET_B_c_855_n N_VPWR_c_1725_n 0.00418607f $X=11.135 $Y=1.665 $X2=0
+ $Y2=0
cc_788 N_RESET_B_c_865_n N_VPWR_c_1728_n 0.0686175f $X=7.46 $Y=3.15 $X2=0 $Y2=0
cc_789 N_RESET_B_c_871_n N_VPWR_c_1730_n 0.00445602f $X=11.32 $Y=2.465 $X2=0
+ $Y2=0
cc_790 N_RESET_B_c_866_n N_VPWR_c_1734_n 0.0506785f $X=3.365 $Y=3.15 $X2=0 $Y2=0
cc_791 N_RESET_B_c_865_n N_VPWR_c_1735_n 0.00797417f $X=7.46 $Y=3.15 $X2=0 $Y2=0
cc_792 N_RESET_B_c_865_n N_VPWR_c_1721_n 0.167656f $X=7.46 $Y=3.15 $X2=0 $Y2=0
cc_793 N_RESET_B_c_866_n N_VPWR_c_1721_n 0.00629086f $X=3.365 $Y=3.15 $X2=0
+ $Y2=0
cc_794 N_RESET_B_c_871_n N_VPWR_c_1721_n 0.00859295f $X=11.32 $Y=2.465 $X2=0
+ $Y2=0
cc_795 N_RESET_B_c_873_n N_VPWR_c_1721_n 3.7828e-19 $X=11.25 $Y=2.375 $X2=0
+ $Y2=0
cc_796 N_RESET_B_M1039_g N_VPWR_c_1741_n 0.00829743f $X=3.29 $Y=2.64 $X2=0 $Y2=0
cc_797 N_RESET_B_c_871_n N_VPWR_c_1744_n 0.00512749f $X=11.32 $Y=2.465 $X2=0
+ $Y2=0
cc_798 N_RESET_B_M1039_g N_A_284_464#_c_1887_n 0.0140389f $X=3.29 $Y=2.64 $X2=0
+ $Y2=0
cc_799 N_RESET_B_c_849_n N_A_284_464#_c_1887_n 0.00126562f $X=3.552 $Y=1.843
+ $X2=0 $Y2=0
cc_800 N_RESET_B_c_859_n N_A_284_464#_c_1887_n 4.86356e-19 $X=3.57 $Y=1.52 $X2=0
+ $Y2=0
cc_801 N_RESET_B_M1026_g N_A_284_464#_c_1862_n 0.0166567f $X=3.445 $Y=0.615
+ $X2=0 $Y2=0
cc_802 N_RESET_B_c_853_n N_A_284_464#_c_1862_n 0.00571983f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_803 N_RESET_B_c_854_n N_A_284_464#_c_1862_n 0.00172645f $X=3.745 $Y=1.665
+ $X2=0 $Y2=0
cc_804 N_RESET_B_c_858_n N_A_284_464#_c_1862_n 0.00558289f $X=3.57 $Y=1.52 $X2=0
+ $Y2=0
cc_805 N_RESET_B_c_859_n N_A_284_464#_c_1862_n 0.0246286f $X=3.57 $Y=1.52 $X2=0
+ $Y2=0
cc_806 N_RESET_B_M1039_g N_A_284_464#_c_1868_n 0.00404939f $X=3.29 $Y=2.64 $X2=0
+ $Y2=0
cc_807 N_RESET_B_c_865_n N_A_284_464#_c_1868_n 0.00532394f $X=7.46 $Y=3.15 $X2=0
+ $Y2=0
cc_808 N_RESET_B_c_865_n N_A_284_464#_c_1870_n 0.00462388f $X=7.46 $Y=3.15 $X2=0
+ $Y2=0
cc_809 N_RESET_B_c_849_n N_A_284_464#_c_1870_n 0.00143051f $X=3.552 $Y=1.843
+ $X2=0 $Y2=0
cc_810 N_RESET_B_c_853_n N_A_284_464#_c_1870_n 0.00555136f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_811 N_RESET_B_c_854_n N_A_284_464#_c_1870_n 6.26496e-19 $X=3.745 $Y=1.665
+ $X2=0 $Y2=0
cc_812 N_RESET_B_c_859_n N_A_284_464#_c_1870_n 0.00418403f $X=3.57 $Y=1.52 $X2=0
+ $Y2=0
cc_813 N_RESET_B_M1039_g N_A_284_464#_c_1871_n 0.00547244f $X=3.29 $Y=2.64 $X2=0
+ $Y2=0
cc_814 N_RESET_B_c_849_n N_A_284_464#_c_1871_n 0.01047f $X=3.552 $Y=1.843 $X2=0
+ $Y2=0
cc_815 N_RESET_B_c_854_n N_A_284_464#_c_1871_n 0.00109964f $X=3.745 $Y=1.665
+ $X2=0 $Y2=0
cc_816 N_RESET_B_c_859_n N_A_284_464#_c_1871_n 0.0207921f $X=3.57 $Y=1.52 $X2=0
+ $Y2=0
cc_817 N_RESET_B_M1026_g N_A_284_464#_c_1946_n 0.00426885f $X=3.445 $Y=0.615
+ $X2=0 $Y2=0
cc_818 N_RESET_B_M1026_g N_A_284_464#_c_1864_n 0.00306727f $X=3.445 $Y=0.615
+ $X2=0 $Y2=0
cc_819 N_RESET_B_c_849_n N_A_284_464#_c_1864_n 0.00301402f $X=3.552 $Y=1.843
+ $X2=0 $Y2=0
cc_820 N_RESET_B_c_853_n N_A_284_464#_c_1864_n 0.0267649f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_821 N_RESET_B_c_854_n N_A_284_464#_c_1864_n 0.00260304f $X=3.745 $Y=1.665
+ $X2=0 $Y2=0
cc_822 N_RESET_B_c_858_n N_A_284_464#_c_1864_n 0.00393379f $X=3.57 $Y=1.52 $X2=0
+ $Y2=0
cc_823 N_RESET_B_c_859_n N_A_284_464#_c_1864_n 0.048278f $X=3.57 $Y=1.52 $X2=0
+ $Y2=0
cc_824 N_RESET_B_M1026_g N_A_284_464#_c_1953_n 0.00167333f $X=3.445 $Y=0.615
+ $X2=0 $Y2=0
cc_825 N_RESET_B_c_865_n N_A_284_464#_c_1873_n 0.011292f $X=7.46 $Y=3.15 $X2=0
+ $Y2=0
cc_826 N_RESET_B_c_853_n N_A_284_464#_c_1873_n 0.00702323f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_827 N_RESET_B_c_853_n N_A_284_464#_c_1874_n 0.00622113f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_828 N_RESET_B_c_865_n N_A_284_464#_c_1875_n 0.00461265f $X=7.46 $Y=3.15 $X2=0
+ $Y2=0
cc_829 N_RESET_B_c_865_n N_A_284_464#_c_1876_n 0.00410507f $X=7.46 $Y=3.15 $X2=0
+ $Y2=0
cc_830 N_RESET_B_c_849_n N_A_284_464#_c_1876_n 8.81721e-19 $X=3.552 $Y=1.843
+ $X2=0 $Y2=0
cc_831 N_RESET_B_M1011_g N_VGND_c_2037_n 0.0026133f $X=7.76 $Y=0.825 $X2=0 $Y2=0
cc_832 N_RESET_B_M1007_g N_VGND_c_2038_n 0.0154281f $X=11.25 $Y=0.58 $X2=0 $Y2=0
cc_833 N_RESET_B_M1007_g N_VGND_c_2044_n 0.00383152f $X=11.25 $Y=0.58 $X2=0
+ $Y2=0
cc_834 N_RESET_B_M1026_g N_VGND_c_2046_n 0.00463377f $X=3.445 $Y=0.615 $X2=0
+ $Y2=0
cc_835 N_RESET_B_M1011_g N_VGND_c_2046_n 7.01746e-19 $X=7.76 $Y=0.825 $X2=0
+ $Y2=0
cc_836 N_RESET_B_M1007_g N_VGND_c_2046_n 0.0075725f $X=11.25 $Y=0.58 $X2=0 $Y2=0
cc_837 N_RESET_B_M1026_g N_VGND_c_2048_n 0.00490893f $X=3.445 $Y=0.615 $X2=0
+ $Y2=0
cc_838 N_RESET_B_M1026_g N_VGND_c_2049_n 9.84134e-19 $X=3.445 $Y=0.615 $X2=0
+ $Y2=0
cc_839 N_RESET_B_M1026_g N_noxref_24_c_2154_n 0.00602133f $X=3.445 $Y=0.615
+ $X2=0 $Y2=0
cc_840 N_RESET_B_M1026_g N_noxref_24_c_2156_n 0.0110823f $X=3.445 $Y=0.615 $X2=0
+ $Y2=0
cc_841 N_A_1251_463#_c_1099_n N_A_854_74#_M1004_g 8.49757e-19 $X=6.57 $Y=2.34
+ $X2=0 $Y2=0
cc_842 N_A_1251_463#_c_1092_n N_A_854_74#_M1004_g 0.00316649f $X=6.97 $Y=2.04
+ $X2=0 $Y2=0
cc_843 N_A_1251_463#_c_1106_n N_A_854_74#_M1004_g 2.81102e-19 $X=6.97 $Y=2.125
+ $X2=0 $Y2=0
cc_844 N_A_1251_463#_c_1092_n N_A_854_74#_c_1224_n 0.00939303f $X=6.97 $Y=2.04
+ $X2=0 $Y2=0
cc_845 N_A_1251_463#_c_1092_n N_A_854_74#_M1014_g 0.00218666f $X=6.97 $Y=2.04
+ $X2=0 $Y2=0
cc_846 N_A_1251_463#_c_1095_n N_A_854_74#_M1014_g 0.010314f $X=6.97 $Y=0.91
+ $X2=0 $Y2=0
cc_847 N_A_1251_463#_c_1091_n N_A_854_74#_c_1226_n 0.00618976f $X=8.35 $Y=1.47
+ $X2=0 $Y2=0
cc_848 N_A_1251_463#_c_1091_n N_A_854_74#_M1038_g 0.0178084f $X=8.35 $Y=1.47
+ $X2=0 $Y2=0
cc_849 N_A_1251_463#_c_1092_n N_A_854_74#_c_1231_n 0.00371216f $X=6.97 $Y=2.04
+ $X2=0 $Y2=0
cc_850 N_A_1251_463#_c_1095_n N_A_854_74#_c_1231_n 0.00912217f $X=6.97 $Y=0.91
+ $X2=0 $Y2=0
cc_851 N_A_1251_463#_c_1094_n N_A_854_74#_c_1235_n 3.94236e-19 $X=8.39 $Y=1.635
+ $X2=0 $Y2=0
cc_852 N_A_1251_463#_c_1094_n N_A_854_74#_c_1236_n 0.0213826f $X=8.39 $Y=1.635
+ $X2=0 $Y2=0
cc_853 N_A_1251_463#_c_1103_n N_VPWR_M1020_s 0.00519751f $X=8.225 $Y=2.055 $X2=0
+ $Y2=0
cc_854 N_A_1251_463#_c_1097_n N_VPWR_c_1724_n 0.00721452f $X=6.405 $Y=2.545
+ $X2=0 $Y2=0
cc_855 N_A_1251_463#_c_1101_n N_VPWR_c_1724_n 0.0138919f $X=7.575 $Y=2.125 $X2=0
+ $Y2=0
cc_856 N_A_1251_463#_c_1102_n N_VPWR_c_1724_n 0.0253299f $X=7.76 $Y=2.545 $X2=0
+ $Y2=0
cc_857 N_A_1251_463#_c_1106_n N_VPWR_c_1724_n 0.00456326f $X=6.97 $Y=2.125 $X2=0
+ $Y2=0
cc_858 N_A_1251_463#_c_1096_n N_VPWR_c_1725_n 0.014528f $X=8.685 $Y=1.885 $X2=0
+ $Y2=0
cc_859 N_A_1251_463#_c_1102_n N_VPWR_c_1725_n 0.0219028f $X=7.76 $Y=2.545 $X2=0
+ $Y2=0
cc_860 N_A_1251_463#_c_1103_n N_VPWR_c_1725_n 0.0197034f $X=8.225 $Y=2.055 $X2=0
+ $Y2=0
cc_861 N_A_1251_463#_c_1094_n N_VPWR_c_1725_n 0.00249414f $X=8.39 $Y=1.635 $X2=0
+ $Y2=0
cc_862 N_A_1251_463#_c_1097_n N_VPWR_c_1728_n 0.00499897f $X=6.405 $Y=2.545
+ $X2=0 $Y2=0
cc_863 N_A_1251_463#_c_1102_n N_VPWR_c_1735_n 0.00726767f $X=7.76 $Y=2.545 $X2=0
+ $Y2=0
cc_864 N_A_1251_463#_c_1096_n N_VPWR_c_1736_n 0.00413917f $X=8.685 $Y=1.885
+ $X2=0 $Y2=0
cc_865 N_A_1251_463#_c_1096_n N_VPWR_c_1721_n 0.00822528f $X=8.685 $Y=1.885
+ $X2=0 $Y2=0
cc_866 N_A_1251_463#_c_1097_n N_VPWR_c_1721_n 0.00757479f $X=6.405 $Y=2.545
+ $X2=0 $Y2=0
cc_867 N_A_1251_463#_c_1102_n N_VPWR_c_1721_n 0.0114703f $X=7.76 $Y=2.545 $X2=0
+ $Y2=0
cc_868 N_A_1251_463#_c_1099_n N_A_284_464#_c_1874_n 0.00765126f $X=6.57 $Y=2.34
+ $X2=0 $Y2=0
cc_869 N_A_1251_463#_c_1098_n A_1341_463# 0.00247499f $X=6.885 $Y=2.34 $X2=-0.19
+ $Y2=-0.245
cc_870 N_A_1251_463#_c_1106_n A_1341_463# 0.00167209f $X=6.97 $Y=2.125 $X2=-0.19
+ $Y2=-0.245
cc_871 N_A_1251_463#_c_1091_n N_VGND_c_2037_n 8.72461e-19 $X=8.35 $Y=1.47 $X2=0
+ $Y2=0
cc_872 N_A_1251_463#_c_1091_n N_VGND_c_2046_n 9.44443e-19 $X=8.35 $Y=1.47 $X2=0
+ $Y2=0
cc_873 N_A_854_74#_c_1229_n N_A_2087_410#_c_1429_n 0.0198038f $X=10.135 $Y=2.375
+ $X2=0 $Y2=0
cc_874 N_A_854_74#_c_1244_n N_A_2087_410#_c_1429_n 0.0337673f $X=10.135 $Y=2.465
+ $X2=0 $Y2=0
cc_875 N_A_854_74#_c_1229_n N_A_2087_410#_M1001_g 0.0152759f $X=10.135 $Y=2.375
+ $X2=0 $Y2=0
cc_876 N_A_854_74#_c_1237_n N_A_2087_410#_M1001_g 0.00123274f $X=10.23 $Y=1.39
+ $X2=0 $Y2=0
cc_877 N_A_854_74#_c_1238_n N_A_2087_410#_M1001_g 0.0187349f $X=10.23 $Y=1.39
+ $X2=0 $Y2=0
cc_878 N_A_854_74#_c_1229_n N_A_2087_410#_c_1435_n 0.00116547f $X=10.135
+ $Y=2.375 $X2=0 $Y2=0
cc_879 N_A_854_74#_c_1244_n N_A_2087_410#_c_1435_n 5.72007e-19 $X=10.135
+ $Y=2.465 $X2=0 $Y2=0
cc_880 N_A_854_74#_c_1229_n N_A_1827_144#_c_1536_n 0.0141151f $X=10.135 $Y=2.375
+ $X2=0 $Y2=0
cc_881 N_A_854_74#_c_1244_n N_A_1827_144#_c_1536_n 0.0133239f $X=10.135 $Y=2.465
+ $X2=0 $Y2=0
cc_882 N_A_854_74#_c_1229_n N_A_1827_144#_c_1537_n 0.0132554f $X=10.135 $Y=2.375
+ $X2=0 $Y2=0
cc_883 N_A_854_74#_c_1237_n N_A_1827_144#_c_1537_n 0.0207258f $X=10.23 $Y=1.39
+ $X2=0 $Y2=0
cc_884 N_A_854_74#_c_1238_n N_A_1827_144#_c_1537_n 0.00380032f $X=10.23 $Y=1.39
+ $X2=0 $Y2=0
cc_885 N_A_854_74#_c_1229_n N_A_1827_144#_c_1538_n 0.00247333f $X=10.135
+ $Y=2.375 $X2=0 $Y2=0
cc_886 N_A_854_74#_c_1235_n N_A_1827_144#_c_1538_n 0.00404793f $X=9.19 $Y=1.455
+ $X2=0 $Y2=0
cc_887 N_A_854_74#_c_1239_n N_A_1827_144#_c_1538_n 0.0218019f $X=10.065 $Y=1.382
+ $X2=0 $Y2=0
cc_888 N_A_854_74#_c_1237_n N_A_1827_144#_c_1525_n 0.015537f $X=10.23 $Y=1.39
+ $X2=0 $Y2=0
cc_889 N_A_854_74#_c_1238_n N_A_1827_144#_c_1525_n 0.0017571f $X=10.23 $Y=1.39
+ $X2=0 $Y2=0
cc_890 N_A_854_74#_c_1237_n N_A_1827_144#_c_1526_n 0.00757275f $X=10.23 $Y=1.39
+ $X2=0 $Y2=0
cc_891 N_A_854_74#_c_1238_n N_A_1827_144#_c_1526_n 8.57186e-19 $X=10.23 $Y=1.39
+ $X2=0 $Y2=0
cc_892 N_A_854_74#_c_1239_n N_A_1827_144#_c_1526_n 0.00315977f $X=10.065
+ $Y=1.382 $X2=0 $Y2=0
cc_893 N_A_854_74#_M1038_g N_A_1827_144#_c_1529_n 0.0152856f $X=9.06 $Y=1.04
+ $X2=0 $Y2=0
cc_894 N_A_854_74#_c_1257_n N_VPWR_M1024_d 0.00398615f $X=4.845 $Y=1.905 $X2=0
+ $Y2=0
cc_895 N_A_854_74#_c_1245_n N_VPWR_M1024_d 9.45391e-19 $X=4.937 $Y=1.82 $X2=0
+ $Y2=0
cc_896 N_A_854_74#_M1028_g N_VPWR_c_1723_n 0.0174456f $X=5.17 $Y=2.235 $X2=0
+ $Y2=0
cc_897 N_A_854_74#_c_1244_n N_VPWR_c_1736_n 0.00456932f $X=10.135 $Y=2.465 $X2=0
+ $Y2=0
cc_898 N_A_854_74#_M1028_g N_VPWR_c_1721_n 8.51577e-19 $X=5.17 $Y=2.235 $X2=0
+ $Y2=0
cc_899 N_A_854_74#_M1004_g N_VPWR_c_1721_n 9.39239e-19 $X=6.18 $Y=2.525 $X2=0
+ $Y2=0
cc_900 N_A_854_74#_c_1244_n N_VPWR_c_1721_n 0.00929427f $X=10.135 $Y=2.465 $X2=0
+ $Y2=0
cc_901 N_A_854_74#_c_1244_n N_VPWR_c_1744_n 0.00148636f $X=10.135 $Y=2.465 $X2=0
+ $Y2=0
cc_902 N_A_854_74#_c_1246_n N_A_284_464#_c_1864_n 0.0143975f $X=4.6 $Y=1.91
+ $X2=0 $Y2=0
cc_903 N_A_854_74#_M1012_d N_A_284_464#_c_1865_n 0.00662096f $X=4.27 $Y=0.37
+ $X2=0 $Y2=0
cc_904 N_A_854_74#_c_1219_n N_A_284_464#_c_1865_n 6.22134e-19 $X=5.17 $Y=1.575
+ $X2=0 $Y2=0
cc_905 N_A_854_74#_c_1220_n N_A_284_464#_c_1865_n 0.0183388f $X=5.295 $Y=1.245
+ $X2=0 $Y2=0
cc_906 N_A_854_74#_c_1221_n N_A_284_464#_c_1865_n 0.0015961f $X=6.105 $Y=1.45
+ $X2=0 $Y2=0
cc_907 N_A_854_74#_c_1232_n N_A_284_464#_c_1865_n 0.0658405f $X=4.845 $Y=0.955
+ $X2=0 $Y2=0
cc_908 N_A_854_74#_c_1233_n N_A_284_464#_c_1865_n 0.00201511f $X=5.17 $Y=1.41
+ $X2=0 $Y2=0
cc_909 N_A_854_74#_M1024_s N_A_284_464#_c_1873_n 0.00967745f $X=4.31 $Y=1.735
+ $X2=0 $Y2=0
cc_910 N_A_854_74#_M1028_g N_A_284_464#_c_1873_n 2.98756e-19 $X=5.17 $Y=2.235
+ $X2=0 $Y2=0
cc_911 N_A_854_74#_c_1257_n N_A_284_464#_c_1873_n 0.00482813f $X=4.845 $Y=1.905
+ $X2=0 $Y2=0
cc_912 N_A_854_74#_c_1246_n N_A_284_464#_c_1873_n 0.0238186f $X=4.6 $Y=1.91
+ $X2=0 $Y2=0
cc_913 N_A_854_74#_c_1219_n N_A_284_464#_c_1874_n 2.27547e-19 $X=5.17 $Y=1.575
+ $X2=0 $Y2=0
cc_914 N_A_854_74#_M1028_g N_A_284_464#_c_1874_n 0.0180037f $X=5.17 $Y=2.235
+ $X2=0 $Y2=0
cc_915 N_A_854_74#_c_1221_n N_A_284_464#_c_1874_n 9.76613e-19 $X=6.105 $Y=1.45
+ $X2=0 $Y2=0
cc_916 N_A_854_74#_M1004_g N_A_284_464#_c_1874_n 0.0065317f $X=6.18 $Y=2.525
+ $X2=0 $Y2=0
cc_917 N_A_854_74#_c_1257_n N_A_284_464#_c_1874_n 0.0186651f $X=4.845 $Y=1.905
+ $X2=0 $Y2=0
cc_918 N_A_854_74#_c_1233_n N_A_284_464#_c_1874_n 0.00248732f $X=5.17 $Y=1.41
+ $X2=0 $Y2=0
cc_919 N_A_854_74#_M1028_g N_A_284_464#_c_1875_n 0.00923143f $X=5.17 $Y=2.235
+ $X2=0 $Y2=0
cc_920 N_A_854_74#_M1004_g N_A_284_464#_c_1875_n 0.00415617f $X=6.18 $Y=2.525
+ $X2=0 $Y2=0
cc_921 N_A_854_74#_c_1220_n N_A_284_464#_c_1866_n 0.00328335f $X=5.295 $Y=1.245
+ $X2=0 $Y2=0
cc_922 N_A_854_74#_c_1221_n N_A_284_464#_c_1866_n 0.00146926f $X=6.105 $Y=1.45
+ $X2=0 $Y2=0
cc_923 N_A_854_74#_c_1232_n N_VGND_M1010_s 0.0072067f $X=4.845 $Y=0.955 $X2=0
+ $Y2=0
cc_924 N_A_854_74#_c_1234_n N_VGND_M1010_s 0.00200761f $X=5.05 $Y=1.235 $X2=0
+ $Y2=0
cc_925 N_A_854_74#_c_1226_n N_VGND_c_2037_n 0.0254808f $X=8.985 $Y=0.2 $X2=0
+ $Y2=0
cc_926 N_A_854_74#_c_1220_n N_VGND_c_2042_n 0.0041773f $X=5.295 $Y=1.245 $X2=0
+ $Y2=0
cc_927 N_A_854_74#_c_1227_n N_VGND_c_2042_n 0.0224126f $X=7.055 $Y=0.2 $X2=0
+ $Y2=0
cc_928 N_A_854_74#_c_1226_n N_VGND_c_2043_n 0.0320058f $X=8.985 $Y=0.2 $X2=0
+ $Y2=0
cc_929 N_A_854_74#_c_1220_n N_VGND_c_2046_n 0.00537853f $X=5.295 $Y=1.245 $X2=0
+ $Y2=0
cc_930 N_A_854_74#_c_1226_n N_VGND_c_2046_n 0.0492768f $X=8.985 $Y=0.2 $X2=0
+ $Y2=0
cc_931 N_A_854_74#_c_1227_n N_VGND_c_2046_n 0.00486765f $X=7.055 $Y=0.2 $X2=0
+ $Y2=0
cc_932 N_A_854_74#_c_1220_n N_VGND_c_2050_n 0.00403889f $X=5.295 $Y=1.245 $X2=0
+ $Y2=0
cc_933 N_A_2087_410#_c_1427_n N_A_1827_144#_c_1517_n 0.0105238f $X=12.065
+ $Y=0.575 $X2=0 $Y2=0
cc_934 N_A_2087_410#_c_1428_n N_A_1827_144#_c_1517_n 0.00492805f $X=12.15
+ $Y=2.29 $X2=0 $Y2=0
cc_935 N_A_2087_410#_c_1428_n N_A_1827_144#_c_1518_n 0.00675601f $X=12.15
+ $Y=2.29 $X2=0 $Y2=0
cc_936 N_A_2087_410#_c_1428_n N_A_1827_144#_c_1519_n 0.00165643f $X=12.15
+ $Y=2.29 $X2=0 $Y2=0
cc_937 N_A_2087_410#_c_1433_n N_A_1827_144#_c_1531_n 0.00495617f $X=12.065
+ $Y=2.375 $X2=0 $Y2=0
cc_938 N_A_2087_410#_c_1428_n N_A_1827_144#_c_1531_n 0.00618531f $X=12.15
+ $Y=2.29 $X2=0 $Y2=0
cc_939 N_A_2087_410#_c_1436_n N_A_1827_144#_c_1531_n 0.00160938f $X=11.545
+ $Y=2.375 $X2=0 $Y2=0
cc_940 N_A_2087_410#_c_1432_n N_A_1827_144#_c_1532_n 0.0124831f $X=11.545
+ $Y=2.75 $X2=0 $Y2=0
cc_941 N_A_2087_410#_c_1433_n N_A_1827_144#_c_1532_n 0.00922094f $X=12.065
+ $Y=2.375 $X2=0 $Y2=0
cc_942 N_A_2087_410#_c_1436_n N_A_1827_144#_c_1532_n 0.00120418f $X=11.545
+ $Y=2.375 $X2=0 $Y2=0
cc_943 N_A_2087_410#_c_1433_n N_A_1827_144#_c_1533_n 0.00361662f $X=12.065
+ $Y=2.375 $X2=0 $Y2=0
cc_944 N_A_2087_410#_c_1428_n N_A_1827_144#_c_1533_n 0.0143738f $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_945 N_A_2087_410#_c_1427_n N_A_1827_144#_c_1520_n 0.00530055f $X=12.065
+ $Y=0.575 $X2=0 $Y2=0
cc_946 N_A_2087_410#_c_1428_n N_A_1827_144#_c_1520_n 0.0145814f $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_947 N_A_2087_410#_c_1428_n N_A_1827_144#_c_1534_n 5.01247e-19 $X=12.15
+ $Y=2.29 $X2=0 $Y2=0
cc_948 N_A_2087_410#_c_1428_n N_A_1827_144#_c_1521_n 7.30697e-19 $X=12.15
+ $Y=2.29 $X2=0 $Y2=0
cc_949 N_A_2087_410#_c_1429_n N_A_1827_144#_c_1536_n 0.00280739f $X=10.545
+ $Y=2.465 $X2=0 $Y2=0
cc_950 N_A_2087_410#_M1001_g N_A_1827_144#_c_1536_n 7.38644e-19 $X=10.69 $Y=0.58
+ $X2=0 $Y2=0
cc_951 N_A_2087_410#_c_1435_n N_A_1827_144#_c_1536_n 0.0164274f $X=10.6 $Y=2.215
+ $X2=0 $Y2=0
cc_952 N_A_2087_410#_c_1429_n N_A_1827_144#_c_1537_n 0.00124779f $X=10.545
+ $Y=2.465 $X2=0 $Y2=0
cc_953 N_A_2087_410#_M1001_g N_A_1827_144#_c_1537_n 0.0120601f $X=10.69 $Y=0.58
+ $X2=0 $Y2=0
cc_954 N_A_2087_410#_c_1431_n N_A_1827_144#_c_1537_n 0.00538841f $X=11.38
+ $Y=2.375 $X2=0 $Y2=0
cc_955 N_A_2087_410#_c_1435_n N_A_1827_144#_c_1537_n 0.017528f $X=10.6 $Y=2.215
+ $X2=0 $Y2=0
cc_956 N_A_2087_410#_M1001_g N_A_1827_144#_c_1525_n 0.0166547f $X=10.69 $Y=0.58
+ $X2=0 $Y2=0
cc_957 N_A_2087_410#_c_1427_n N_A_1827_144#_c_1525_n 0.0151071f $X=12.065
+ $Y=0.575 $X2=0 $Y2=0
cc_958 N_A_2087_410#_c_1428_n N_A_1827_144#_c_1525_n 0.0135536f $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_959 N_A_2087_410#_c_1431_n N_A_1827_144#_c_1539_n 0.024548f $X=11.38 $Y=2.375
+ $X2=0 $Y2=0
cc_960 N_A_2087_410#_c_1433_n N_A_1827_144#_c_1539_n 0.0143017f $X=12.065
+ $Y=2.375 $X2=0 $Y2=0
cc_961 N_A_2087_410#_c_1428_n N_A_1827_144#_c_1539_n 0.0135702f $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_962 N_A_2087_410#_c_1436_n N_A_1827_144#_c_1539_n 0.0286194f $X=11.545
+ $Y=2.375 $X2=0 $Y2=0
cc_963 N_A_2087_410#_c_1428_n N_A_1827_144#_c_1527_n 0.0689819f $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_964 N_A_2087_410#_c_1427_n N_A_1827_144#_c_1528_n 0.0010568f $X=12.065
+ $Y=0.575 $X2=0 $Y2=0
cc_965 N_A_2087_410#_c_1428_n N_A_1827_144#_c_1528_n 6.697e-19 $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_966 N_A_2087_410#_M1001_g N_A_1827_144#_c_1541_n 0.00514664f $X=10.69 $Y=0.58
+ $X2=0 $Y2=0
cc_967 N_A_2087_410#_c_1431_n N_A_1827_144#_c_1541_n 0.0132541f $X=11.38
+ $Y=2.375 $X2=0 $Y2=0
cc_968 N_A_2087_410#_c_1435_n N_A_1827_144#_c_1541_n 0.00515102f $X=10.6
+ $Y=2.215 $X2=0 $Y2=0
cc_969 N_A_2087_410#_c_1428_n N_A_2492_424#_c_1677_n 0.00119502f $X=12.15
+ $Y=2.29 $X2=0 $Y2=0
cc_970 N_A_2087_410#_c_1427_n N_A_2492_424#_c_1679_n 0.0191493f $X=12.065
+ $Y=0.575 $X2=0 $Y2=0
cc_971 N_A_2087_410#_c_1428_n N_A_2492_424#_c_1679_n 0.108701f $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_972 N_A_2087_410#_c_1433_n N_A_2492_424#_c_1684_n 0.013247f $X=12.065
+ $Y=2.375 $X2=0 $Y2=0
cc_973 N_A_2087_410#_c_1432_n N_VPWR_c_1726_n 0.0139233f $X=11.545 $Y=2.75 $X2=0
+ $Y2=0
cc_974 N_A_2087_410#_c_1433_n N_VPWR_c_1726_n 0.0274592f $X=12.065 $Y=2.375
+ $X2=0 $Y2=0
cc_975 N_A_2087_410#_c_1432_n N_VPWR_c_1730_n 0.0145674f $X=11.545 $Y=2.75 $X2=0
+ $Y2=0
cc_976 N_A_2087_410#_c_1429_n N_VPWR_c_1736_n 0.00415318f $X=10.545 $Y=2.465
+ $X2=0 $Y2=0
cc_977 N_A_2087_410#_c_1429_n N_VPWR_c_1721_n 0.00852129f $X=10.545 $Y=2.465
+ $X2=0 $Y2=0
cc_978 N_A_2087_410#_c_1432_n N_VPWR_c_1721_n 0.0119851f $X=11.545 $Y=2.75 $X2=0
+ $Y2=0
cc_979 N_A_2087_410#_c_1429_n N_VPWR_c_1744_n 0.0173099f $X=10.545 $Y=2.465
+ $X2=0 $Y2=0
cc_980 N_A_2087_410#_c_1431_n N_VPWR_c_1744_n 0.0390885f $X=11.38 $Y=2.375 $X2=0
+ $Y2=0
cc_981 N_A_2087_410#_c_1432_n N_VPWR_c_1744_n 0.0132487f $X=11.545 $Y=2.75 $X2=0
+ $Y2=0
cc_982 N_A_2087_410#_c_1435_n N_VPWR_c_1744_n 0.00383575f $X=10.6 $Y=2.215 $X2=0
+ $Y2=0
cc_983 N_A_2087_410#_M1001_g N_VGND_c_2038_n 0.0163013f $X=10.69 $Y=0.58 $X2=0
+ $Y2=0
cc_984 N_A_2087_410#_c_1427_n N_VGND_c_2038_n 0.00776169f $X=12.065 $Y=0.575
+ $X2=0 $Y2=0
cc_985 N_A_2087_410#_M1001_g N_VGND_c_2043_n 0.00352388f $X=10.69 $Y=0.58 $X2=0
+ $Y2=0
cc_986 N_A_2087_410#_c_1427_n N_VGND_c_2044_n 0.015221f $X=12.065 $Y=0.575 $X2=0
+ $Y2=0
cc_987 N_A_2087_410#_M1001_g N_VGND_c_2046_n 0.0069736f $X=10.69 $Y=0.58 $X2=0
+ $Y2=0
cc_988 N_A_2087_410#_c_1427_n N_VGND_c_2046_n 0.0182599f $X=12.065 $Y=0.575
+ $X2=0 $Y2=0
cc_989 N_A_1827_144#_c_1534_n N_A_2492_424#_c_1681_n 0.0112885f $X=12.83
+ $Y=2.045 $X2=0 $Y2=0
cc_990 N_A_1827_144#_c_1521_n N_A_2492_424#_M1015_g 0.0139661f $X=12.845
+ $Y=0.995 $X2=0 $Y2=0
cc_991 N_A_1827_144#_c_1518_n N_A_2492_424#_c_1677_n 0.00295561f $X=11.73
+ $Y=1.405 $X2=0 $Y2=0
cc_992 N_A_1827_144#_c_1519_n N_A_2492_424#_c_1677_n 0.00131811f $X=11.755
+ $Y=1.895 $X2=0 $Y2=0
cc_993 N_A_1827_144#_c_1533_n N_A_2492_424#_c_1677_n 0.0299671f $X=12.755
+ $Y=1.97 $X2=0 $Y2=0
cc_994 N_A_1827_144#_c_1520_n N_A_2492_424#_c_1677_n 0.030045f $X=12.77 $Y=1.07
+ $X2=0 $Y2=0
cc_995 N_A_1827_144#_c_1520_n N_A_2492_424#_c_1679_n 0.0201885f $X=12.77 $Y=1.07
+ $X2=0 $Y2=0
cc_996 N_A_1827_144#_c_1521_n N_A_2492_424#_c_1679_n 0.012287f $X=12.845
+ $Y=0.995 $X2=0 $Y2=0
cc_997 N_A_1827_144#_c_1531_n N_A_2492_424#_c_1684_n 8.46777e-19 $X=11.77
+ $Y=2.375 $X2=0 $Y2=0
cc_998 N_A_1827_144#_c_1532_n N_A_2492_424#_c_1684_n 0.00465863f $X=11.77
+ $Y=2.465 $X2=0 $Y2=0
cc_999 N_A_1827_144#_c_1533_n N_A_2492_424#_c_1684_n 0.0177354f $X=12.755
+ $Y=1.97 $X2=0 $Y2=0
cc_1000 N_A_1827_144#_c_1534_n N_A_2492_424#_c_1684_n 0.0163542f $X=12.83
+ $Y=2.045 $X2=0 $Y2=0
cc_1001 N_A_1827_144#_c_1532_n N_VPWR_c_1726_n 0.010223f $X=11.77 $Y=2.465 $X2=0
+ $Y2=0
cc_1002 N_A_1827_144#_c_1533_n N_VPWR_c_1726_n 6.69985e-19 $X=12.755 $Y=1.97
+ $X2=0 $Y2=0
cc_1003 N_A_1827_144#_c_1534_n N_VPWR_c_1726_n 0.00334683f $X=12.83 $Y=2.045
+ $X2=0 $Y2=0
cc_1004 N_A_1827_144#_c_1533_n N_VPWR_c_1727_n 0.00177592f $X=12.755 $Y=1.97
+ $X2=0 $Y2=0
cc_1005 N_A_1827_144#_c_1534_n N_VPWR_c_1727_n 0.011687f $X=12.83 $Y=2.045 $X2=0
+ $Y2=0
cc_1006 N_A_1827_144#_c_1532_n N_VPWR_c_1730_n 0.00445602f $X=11.77 $Y=2.465
+ $X2=0 $Y2=0
cc_1007 N_A_1827_144#_c_1536_n N_VPWR_c_1736_n 0.0146237f $X=9.845 $Y=2.135
+ $X2=0 $Y2=0
cc_1008 N_A_1827_144#_c_1534_n N_VPWR_c_1737_n 0.00417277f $X=12.83 $Y=2.045
+ $X2=0 $Y2=0
cc_1009 N_A_1827_144#_c_1532_n N_VPWR_c_1721_n 0.00898236f $X=11.77 $Y=2.465
+ $X2=0 $Y2=0
cc_1010 N_A_1827_144#_c_1534_n N_VPWR_c_1721_n 0.00771913f $X=12.83 $Y=2.045
+ $X2=0 $Y2=0
cc_1011 N_A_1827_144#_c_1536_n N_VPWR_c_1721_n 0.0120948f $X=9.845 $Y=2.135
+ $X2=0 $Y2=0
cc_1012 N_A_1827_144#_c_1536_n N_VPWR_c_1744_n 0.0100622f $X=9.845 $Y=2.135
+ $X2=0 $Y2=0
cc_1013 N_A_1827_144#_c_1520_n Q 2.35526e-19 $X=12.77 $Y=1.07 $X2=0 $Y2=0
cc_1014 N_A_1827_144#_c_1517_n N_VGND_c_2038_n 0.0017037f $X=11.64 $Y=0.9 $X2=0
+ $Y2=0
cc_1015 N_A_1827_144#_c_1523_n N_VGND_c_2038_n 0.00644386f $X=10.08 $Y=0.62
+ $X2=0 $Y2=0
cc_1016 N_A_1827_144#_c_1525_n N_VGND_c_2038_n 0.0305939f $X=11.565 $Y=0.955
+ $X2=0 $Y2=0
cc_1017 N_A_1827_144#_c_1521_n N_VGND_c_2039_n 0.00901588f $X=12.845 $Y=0.995
+ $X2=0 $Y2=0
cc_1018 N_A_1827_144#_c_1523_n N_VGND_c_2043_n 0.00997274f $X=10.08 $Y=0.62
+ $X2=0 $Y2=0
cc_1019 N_A_1827_144#_c_1529_n N_VGND_c_2043_n 0.0445263f $X=9.995 $Y=0.455
+ $X2=0 $Y2=0
cc_1020 N_A_1827_144#_c_1517_n N_VGND_c_2044_n 0.00435333f $X=11.64 $Y=0.9 $X2=0
+ $Y2=0
cc_1021 N_A_1827_144#_c_1521_n N_VGND_c_2044_n 0.00434272f $X=12.845 $Y=0.995
+ $X2=0 $Y2=0
cc_1022 N_A_1827_144#_c_1517_n N_VGND_c_2046_n 0.00824743f $X=11.64 $Y=0.9 $X2=0
+ $Y2=0
cc_1023 N_A_1827_144#_c_1521_n N_VGND_c_2046_n 0.00826607f $X=12.845 $Y=0.995
+ $X2=0 $Y2=0
cc_1024 N_A_1827_144#_c_1523_n N_VGND_c_2046_n 0.00649523f $X=10.08 $Y=0.62
+ $X2=0 $Y2=0
cc_1025 N_A_1827_144#_c_1529_n N_VGND_c_2046_n 0.0301144f $X=9.995 $Y=0.455
+ $X2=0 $Y2=0
cc_1026 N_A_2492_424#_c_1684_n N_VPWR_c_1726_n 0.0237277f $X=12.605 $Y=2.265
+ $X2=0 $Y2=0
cc_1027 N_A_2492_424#_c_1681_n N_VPWR_c_1727_n 0.00423469f $X=13.41 $Y=1.765
+ $X2=0 $Y2=0
cc_1028 N_A_2492_424#_c_1677_n N_VPWR_c_1727_n 0.0151403f $X=13.32 $Y=1.52 $X2=0
+ $Y2=0
cc_1029 N_A_2492_424#_c_1684_n N_VPWR_c_1727_n 0.0873946f $X=12.605 $Y=2.265
+ $X2=0 $Y2=0
cc_1030 N_A_2492_424#_c_1684_n N_VPWR_c_1737_n 0.0156346f $X=12.605 $Y=2.265
+ $X2=0 $Y2=0
cc_1031 N_A_2492_424#_c_1681_n N_VPWR_c_1738_n 0.00451267f $X=13.41 $Y=1.765
+ $X2=0 $Y2=0
cc_1032 N_A_2492_424#_c_1681_n N_VPWR_c_1721_n 0.00879786f $X=13.41 $Y=1.765
+ $X2=0 $Y2=0
cc_1033 N_A_2492_424#_c_1684_n N_VPWR_c_1721_n 0.0128494f $X=12.605 $Y=2.265
+ $X2=0 $Y2=0
cc_1034 N_A_2492_424#_c_1681_n Q 0.0160775f $X=13.41 $Y=1.765 $X2=0 $Y2=0
cc_1035 N_A_2492_424#_M1015_g Q 0.0241875f $X=13.425 $Y=0.74 $X2=0 $Y2=0
cc_1036 N_A_2492_424#_c_1678_n Q 0.0226991f $X=13.41 $Y=1.56 $X2=0 $Y2=0
cc_1037 N_A_2492_424#_c_1680_n Q 0.00799574f $X=12.645 $Y=1.52 $X2=0 $Y2=0
cc_1038 N_A_2492_424#_M1015_g N_VGND_c_2039_n 0.0060503f $X=13.425 $Y=0.74 $X2=0
+ $Y2=0
cc_1039 N_A_2492_424#_c_1677_n N_VGND_c_2039_n 0.0137394f $X=13.32 $Y=1.52 $X2=0
+ $Y2=0
cc_1040 N_A_2492_424#_c_1679_n N_VGND_c_2039_n 0.0373449f $X=12.63 $Y=0.645
+ $X2=0 $Y2=0
cc_1041 N_A_2492_424#_c_1679_n N_VGND_c_2044_n 0.0156794f $X=12.63 $Y=0.645
+ $X2=0 $Y2=0
cc_1042 N_A_2492_424#_M1015_g N_VGND_c_2045_n 0.00434272f $X=13.425 $Y=0.74
+ $X2=0 $Y2=0
cc_1043 N_A_2492_424#_M1015_g N_VGND_c_2046_n 0.00825042f $X=13.425 $Y=0.74
+ $X2=0 $Y2=0
cc_1044 N_A_2492_424#_c_1679_n N_VGND_c_2046_n 0.0129217f $X=12.63 $Y=0.645
+ $X2=0 $Y2=0
cc_1045 N_VPWR_M1016_d N_A_284_464#_c_1887_n 0.0104678f $X=2.745 $Y=2.32 $X2=0
+ $Y2=0
cc_1046 N_VPWR_c_1733_n N_A_284_464#_c_1887_n 0.0103117f $X=2.815 $Y=3.33 $X2=0
+ $Y2=0
cc_1047 N_VPWR_c_1734_n N_A_284_464#_c_1887_n 0.0043953f $X=4.78 $Y=3.33 $X2=0
+ $Y2=0
cc_1048 N_VPWR_c_1721_n N_A_284_464#_c_1887_n 0.0240636f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1049 N_VPWR_c_1741_n N_A_284_464#_c_1887_n 0.0241556f $X=2.98 $Y=3.055 $X2=0
+ $Y2=0
cc_1050 N_VPWR_c_1734_n N_A_284_464#_c_1868_n 0.0111464f $X=4.78 $Y=3.33 $X2=0
+ $Y2=0
cc_1051 N_VPWR_c_1721_n N_A_284_464#_c_1868_n 0.00823093f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1052 N_VPWR_c_1741_n N_A_284_464#_c_1868_n 5.70141e-19 $X=2.98 $Y=3.055 $X2=0
+ $Y2=0
cc_1053 N_VPWR_M1024_d N_A_284_464#_c_1874_n 0.00389705f $X=4.795 $Y=1.735 $X2=0
+ $Y2=0
cc_1054 N_VPWR_c_1723_n N_A_284_464#_c_1874_n 0.0171814f $X=4.945 $Y=2.585 $X2=0
+ $Y2=0
cc_1055 N_VPWR_c_1728_n N_A_284_464#_c_1875_n 0.00478298f $X=7.225 $Y=3.33 $X2=0
+ $Y2=0
cc_1056 N_VPWR_c_1721_n N_A_284_464#_c_1875_n 0.00695772f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1057 N_VPWR_c_1722_n N_A_284_464#_c_1884_n 0.0106407f $X=0.73 $Y=2.805 $X2=0
+ $Y2=0
cc_1058 N_VPWR_c_1733_n N_A_284_464#_c_1884_n 0.0290068f $X=2.815 $Y=3.33 $X2=0
+ $Y2=0
cc_1059 N_VPWR_c_1721_n N_A_284_464#_c_1884_n 0.0288251f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1060 N_VPWR_c_1727_n Q 0.0451069f $X=13.14 $Y=1.985 $X2=0 $Y2=0
cc_1061 N_VPWR_c_1738_n Q 0.0146088f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1062 N_VPWR_c_1721_n Q 0.0120707f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1063 N_A_284_464#_c_1887_n A_471_464# 0.00325808f $X=3.43 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_1064 N_A_284_464#_c_1862_n N_VGND_M1026_d 8.85948e-19 $X=3.905 $Y=1.1 $X2=0
+ $Y2=0
cc_1065 N_A_284_464#_c_1946_n N_VGND_M1026_d 0.00597038f $X=3.99 $Y=1.015 $X2=0
+ $Y2=0
cc_1066 N_A_284_464#_c_1953_n N_VGND_M1026_d 0.00458913f $X=4.075 $Y=0.615 $X2=0
+ $Y2=0
cc_1067 N_A_284_464#_c_1867_n N_VGND_M1026_d 8.30808e-19 $X=3.99 $Y=1.1 $X2=0
+ $Y2=0
cc_1068 N_A_284_464#_c_1865_n N_VGND_M1010_s 0.00878709f $X=5.905 $Y=0.615 $X2=0
+ $Y2=0
cc_1069 N_A_284_464#_c_1865_n N_VGND_c_2041_n 0.0154055f $X=5.905 $Y=0.615 $X2=0
+ $Y2=0
cc_1070 N_A_284_464#_c_1865_n N_VGND_c_2042_n 0.0218488f $X=5.905 $Y=0.615 $X2=0
+ $Y2=0
cc_1071 N_A_284_464#_c_1865_n N_VGND_c_2046_n 0.0548314f $X=5.905 $Y=0.615 $X2=0
+ $Y2=0
cc_1072 N_A_284_464#_c_1953_n N_VGND_c_2046_n 0.00133036f $X=4.075 $Y=0.615
+ $X2=0 $Y2=0
cc_1073 N_A_284_464#_c_1862_n N_VGND_c_2049_n 0.00983574f $X=3.905 $Y=1.1 $X2=0
+ $Y2=0
cc_1074 N_A_284_464#_c_1953_n N_VGND_c_2049_n 0.0128556f $X=4.075 $Y=0.615 $X2=0
+ $Y2=0
cc_1075 N_A_284_464#_c_1865_n N_VGND_c_2050_n 0.0263497f $X=5.905 $Y=0.615 $X2=0
+ $Y2=0
cc_1076 N_A_284_464#_c_1877_n N_noxref_24_c_2153_n 0.00596172f $X=2.72 $Y=0.68
+ $X2=0 $Y2=0
cc_1077 N_A_284_464#_M1022_d N_noxref_24_c_2154_n 0.00467414f $X=1.98 $Y=0.405
+ $X2=0 $Y2=0
cc_1078 N_A_284_464#_c_1877_n N_noxref_24_c_2154_n 0.0511317f $X=2.72 $Y=0.68
+ $X2=0 $Y2=0
cc_1079 N_A_284_464#_c_1862_n N_noxref_24_c_2154_n 0.00375974f $X=3.905 $Y=1.1
+ $X2=0 $Y2=0
cc_1080 N_A_284_464#_c_1861_n N_noxref_24_c_2156_n 0.00371663f $X=2.805 $Y=1.015
+ $X2=0 $Y2=0
cc_1081 N_A_284_464#_c_1862_n N_noxref_24_c_2156_n 0.0270682f $X=3.905 $Y=1.1
+ $X2=0 $Y2=0
cc_1082 N_A_284_464#_c_1946_n N_noxref_24_c_2156_n 0.00449664f $X=3.99 $Y=1.015
+ $X2=0 $Y2=0
cc_1083 N_A_284_464#_c_1953_n N_noxref_24_c_2156_n 0.0059249f $X=4.075 $Y=0.615
+ $X2=0 $Y2=0
cc_1084 N_A_284_464#_c_1877_n noxref_26 0.00135313f $X=2.72 $Y=0.68 $X2=-0.19
+ $Y2=-0.245
cc_1085 Q N_VGND_c_2039_n 0.0308485f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1086 Q N_VGND_c_2045_n 0.0145639f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1087 Q N_VGND_c_2046_n 0.0119984f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1088 N_VGND_c_2036_n N_noxref_24_c_2153_n 0.0236042f $X=0.78 $Y=0.65 $X2=0
+ $Y2=0
cc_1089 N_VGND_c_2046_n N_noxref_24_c_2154_n 0.071615f $X=13.68 $Y=0 $X2=0 $Y2=0
cc_1090 N_VGND_c_2048_n N_noxref_24_c_2154_n 0.124162f $X=3.575 $Y=0.137 $X2=0
+ $Y2=0
cc_1091 N_VGND_c_2049_n N_noxref_24_c_2154_n 0.00856573f $X=4.065 $Y=0.137 $X2=0
+ $Y2=0
cc_1092 N_VGND_c_2036_n N_noxref_24_c_2155_n 0.0125438f $X=0.78 $Y=0.65 $X2=0
+ $Y2=0
cc_1093 N_VGND_c_2046_n N_noxref_24_c_2155_n 0.0127354f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1094 N_VGND_c_2048_n N_noxref_24_c_2155_n 0.0231539f $X=3.575 $Y=0.137 $X2=0
+ $Y2=0
cc_1095 N_noxref_24_c_2154_n noxref_25 0.00366293f $X=3.06 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1096 N_noxref_24_c_2154_n noxref_26 0.0013394f $X=3.06 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
