* File: sky130_fd_sc_ls__a32oi_2.pex.spice
* Created: Wed Sep  2 10:53:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A32OI_2%B2 3 5 7 10 12 14 17 20 25 30
r48 25 26 3.59701 $w=4.02e-07 $l=3e-08 $layer=POLY_cond $X=0.975 $Y=1.532
+ $X2=1.005 $Y2=1.532
r49 22 23 1.79851 $w=4.02e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.532
+ $X2=0.51 $Y2=1.532
r50 20 30 4.04332 $w=4.78e-07 $l=1.15e-07 $layer=LI1_cond $X=0.24 $Y=1.54
+ $X2=0.355 $Y2=1.54
r51 18 25 5.99502 $w=4.02e-07 $l=5e-08 $layer=POLY_cond $X=0.925 $Y=1.532
+ $X2=0.975 $Y2=1.532
r52 18 23 49.7587 $w=4.02e-07 $l=4.15e-07 $layer=POLY_cond $X=0.925 $Y=1.532
+ $X2=0.51 $Y2=1.532
r53 17 30 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=0.925 $Y=1.465
+ $X2=0.355 $Y2=1.465
r54 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.925
+ $Y=1.465 $X2=0.925 $Y2=1.465
r55 12 26 25.9839 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=1.532
r56 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r57 8 25 25.9839 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.975 $Y=1.3
+ $X2=0.975 $Y2=1.532
r58 8 10 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.975 $Y=1.3
+ $X2=0.975 $Y2=0.74
r59 5 23 25.9839 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.532
r60 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r61 1 22 25.9839 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.532
r62 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A32OI_2%B1 1 3 4 6 7 9 10 12 13 14 20
c56 7 0 1.33933e-19 $X=1.835 $Y=1.22
c57 1 0 8.87788e-21 $X=1.405 $Y=1.22
r58 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.01
+ $Y=1.385 $X2=2.01 $Y2=1.385
r59 20 22 0.598015 $w=4.03e-07 $l=5e-09 $layer=POLY_cond $X=2.005 $Y=1.492
+ $X2=2.01 $Y2=1.492
r60 19 20 20.3325 $w=4.03e-07 $l=1.7e-07 $layer=POLY_cond $X=1.835 $Y=1.492
+ $X2=2.005 $Y2=1.492
r61 18 19 39.469 $w=4.03e-07 $l=3.3e-07 $layer=POLY_cond $X=1.505 $Y=1.492
+ $X2=1.835 $Y2=1.492
r62 14 23 4.67207 $w=3.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.16 $Y=1.365
+ $X2=2.01 $Y2=1.365
r63 13 23 10.2785 $w=3.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=2.01 $Y2=1.365
r64 10 20 26.0447 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.005 $Y=1.765
+ $X2=2.005 $Y2=1.492
r65 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.005 $Y=1.765
+ $X2=2.005 $Y2=2.4
r66 7 19 26.0447 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.835 $Y=1.22
+ $X2=1.835 $Y2=1.492
r67 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.835 $Y=1.22 $X2=1.835
+ $Y2=0.74
r68 4 18 26.0447 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=1.492
r69 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=2.4
r70 1 18 11.9603 $w=4.03e-07 $l=3.18094e-07 $layer=POLY_cond $X=1.405 $Y=1.22
+ $X2=1.505 $Y2=1.492
r71 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.405 $Y=1.22 $X2=1.405
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A32OI_2%A1 1 3 4 6 7 9 10 12 13 20
c55 13 0 1.33933e-19 $X=2.64 $Y=1.295
c56 10 0 2.88763e-19 $X=3.345 $Y=1.765
r57 20 21 2.38025 $w=4.05e-07 $l=2e-08 $layer=POLY_cond $X=3.325 $Y=1.492
+ $X2=3.345 $Y2=1.492
r58 19 20 51.1753 $w=4.05e-07 $l=4.3e-07 $layer=POLY_cond $X=2.895 $Y=1.492
+ $X2=3.325 $Y2=1.492
r59 17 19 33.9185 $w=4.05e-07 $l=2.85e-07 $layer=POLY_cond $X=2.61 $Y=1.492
+ $X2=2.895 $Y2=1.492
r60 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.385 $X2=2.61 $Y2=1.385
r61 15 17 12.4963 $w=4.05e-07 $l=1.05e-07 $layer=POLY_cond $X=2.505 $Y=1.492
+ $X2=2.61 $Y2=1.492
r62 13 18 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.61 $Y=1.295 $X2=2.61
+ $Y2=1.385
r63 10 21 26.1659 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.345 $Y=1.765
+ $X2=3.345 $Y2=1.492
r64 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.345 $Y=1.765
+ $X2=3.345 $Y2=2.4
r65 7 20 26.1659 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.325 $Y=1.22
+ $X2=3.325 $Y2=1.492
r66 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.325 $Y=1.22 $X2=3.325
+ $Y2=0.74
r67 4 19 26.1659 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.895 $Y=1.22
+ $X2=2.895 $Y2=1.492
r68 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.895 $Y=1.22 $X2=2.895
+ $Y2=0.74
r69 1 15 26.1659 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.505 $Y=1.765
+ $X2=2.505 $Y2=1.492
r70 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.505 $Y=1.765
+ $X2=2.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A32OI_2%A2 3 5 7 8 10 13 16 17 18 19 20 25
c58 25 0 1.42489e-19 $X=4.21 $Y=1.515
c59 16 0 1.39445e-19 $X=3.795 $Y=1.557
c60 8 0 1.85225e-19 $X=4.31 $Y=1.765
c61 3 0 5.89156e-20 $X=3.78 $Y=0.74
r62 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.21
+ $Y=1.515 $X2=4.21 $Y2=1.515
r63 20 25 3.48413 $w=4.28e-07 $l=1.3e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=4.21 $Y2=1.565
r64 19 20 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=4.08 $Y2=1.565
r65 17 24 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=4.22 $Y=1.515 $X2=4.21
+ $Y2=1.515
r66 17 18 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=4.22 $Y=1.515
+ $X2=4.31 $Y2=1.557
r67 15 24 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=3.885 $Y=1.515
+ $X2=4.21 $Y2=1.515
r68 15 16 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=3.885 $Y=1.515
+ $X2=3.795 $Y2=1.557
r69 11 18 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=4.325 $Y=1.35
+ $X2=4.31 $Y2=1.557
r70 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.325 $Y=1.35
+ $X2=4.325 $Y2=0.74
r71 8 18 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.31 $Y=1.765
+ $X2=4.31 $Y2=1.557
r72 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.31 $Y=1.765
+ $X2=4.31 $Y2=2.4
r73 5 16 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.795 $Y=1.765
+ $X2=3.795 $Y2=1.557
r74 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.795 $Y=1.765
+ $X2=3.795 $Y2=2.4
r75 1 16 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=3.78 $Y=1.35
+ $X2=3.795 $Y2=1.557
r76 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.78 $Y=1.35 $X2=3.78
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__A32OI_2%A3 1 3 4 6 7 9 10 12 13 18
c41 1 0 1.0634e-20 $X=4.935 $Y=1.765
r42 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.95
+ $Y=1.385 $X2=5.95 $Y2=1.385
r43 18 20 25.3359 $w=3.9e-07 $l=2.05e-07 $layer=POLY_cond $X=5.745 $Y=1.492
+ $X2=5.95 $Y2=1.492
r44 17 18 32.1333 $w=3.9e-07 $l=2.6e-07 $layer=POLY_cond $X=5.485 $Y=1.492
+ $X2=5.745 $Y2=1.492
r45 16 17 21.0103 $w=3.9e-07 $l=1.7e-07 $layer=POLY_cond $X=5.315 $Y=1.492
+ $X2=5.485 $Y2=1.492
r46 15 16 46.9641 $w=3.9e-07 $l=3.8e-07 $layer=POLY_cond $X=4.935 $Y=1.492
+ $X2=5.315 $Y2=1.492
r47 13 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.95 $Y=1.295 $X2=5.95
+ $Y2=1.385
r48 10 18 25.2441 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=5.745 $Y=1.22
+ $X2=5.745 $Y2=1.492
r49 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.745 $Y=1.22
+ $X2=5.745 $Y2=0.74
r50 7 17 25.2441 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=5.485 $Y=1.765
+ $X2=5.485 $Y2=1.492
r51 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.485 $Y=1.765
+ $X2=5.485 $Y2=2.4
r52 4 16 25.2441 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=5.315 $Y=1.22
+ $X2=5.315 $Y2=1.492
r53 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.315 $Y=1.22 $X2=5.315
+ $Y2=0.74
r54 1 15 25.2441 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.935 $Y=1.765
+ $X2=4.935 $Y2=1.492
r55 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.935 $Y=1.765
+ $X2=4.935 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LS__A32OI_2%A_27_368# 1 2 3 4 5 6 21 25 26 29 31 33 37
+ 41 43 45 47 49 53 57 60
c87 41 0 3.42133e-19 $X=3.57 $Y=2.465
r88 68 69 1.59269 $w=3.83e-07 $l=5e-08 $layer=LI1_cond $X=4.647 $Y=1.985
+ $X2=4.647 $Y2=2.035
r89 66 68 5.73368 $w=3.83e-07 $l=1.8e-07 $layer=LI1_cond $X=4.647 $Y=1.805
+ $X2=4.647 $Y2=1.985
r90 64 65 3.21434 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=2.145
+ $X2=3.57 $Y2=2.23
r91 63 64 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=3.57 $Y=2.115 $X2=3.57
+ $Y2=2.145
r92 60 63 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.57 $Y=2.035 $X2=3.57
+ $Y2=2.115
r93 53 55 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.71 $Y=1.985
+ $X2=5.71 $Y2=2.815
r94 51 53 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.71 $Y=1.89
+ $X2=5.71 $Y2=1.985
r95 50 66 5.51523 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=4.875 $Y=1.805
+ $X2=4.647 $Y2=1.805
r96 49 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.545 $Y=1.805
+ $X2=5.71 $Y2=1.89
r97 49 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.545 $Y=1.805
+ $X2=4.875 $Y2=1.805
r98 45 69 2.6202 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.647 $Y=2.12
+ $X2=4.647 $Y2=2.035
r99 45 47 7.36048 $w=4.53e-07 $l=2.8e-07 $layer=LI1_cond $X=4.647 $Y=2.12
+ $X2=4.647 $Y2=2.4
r100 44 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.735 $Y=2.035
+ $X2=3.57 $Y2=2.035
r101 43 69 5.51523 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=4.42 $Y=2.035
+ $X2=4.647 $Y2=2.035
r102 43 44 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.42 $Y=2.035
+ $X2=3.735 $Y2=2.035
r103 41 65 9.5026 $w=2.83e-07 $l=2.35e-07 $layer=LI1_cond $X=3.592 $Y=2.465
+ $X2=3.592 $Y2=2.23
r104 38 59 4.64039 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=2.4 $Y=2.145
+ $X2=2.257 $Y2=2.145
r105 37 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=2.145
+ $X2=3.57 $Y2=2.145
r106 37 38 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=3.405 $Y=2.145
+ $X2=2.4 $Y2=2.145
r107 34 36 16.579 $w=2.83e-07 $l=4.1e-07 $layer=LI1_cond $X=2.257 $Y=2.905
+ $X2=2.257 $Y2=2.495
r108 33 59 2.75828 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.257 $Y=2.23
+ $X2=2.257 $Y2=2.145
r109 33 36 10.7157 $w=2.83e-07 $l=2.65e-07 $layer=LI1_cond $X=2.257 $Y=2.23
+ $X2=2.257 $Y2=2.495
r110 32 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=2.99
+ $X2=1.28 $Y2=2.99
r111 31 34 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=2.115 $Y=2.99
+ $X2=2.257 $Y2=2.905
r112 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=2.99
+ $X2=1.445 $Y2=2.99
r113 27 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=2.905
+ $X2=1.28 $Y2=2.99
r114 27 29 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.28 $Y=2.905
+ $X2=1.28 $Y2=2.27
r115 25 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=1.28 $Y2=2.99
r116 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=0.445 $Y2=2.99
r117 21 24 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115
+ $X2=0.28 $Y2=2.815
r118 19 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r119 19 24 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.28 $Y2=2.815
r120 6 55 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.56
+ $Y=1.84 $X2=5.71 $Y2=2.815
r121 6 53 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.56
+ $Y=1.84 $X2=5.71 $Y2=1.985
r122 5 68 600 $w=1.7e-07 $l=3.90832e-07 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.84 $X2=4.71 $Y2=1.985
r123 5 47 300 $w=1.7e-07 $l=6.5238e-07 $layer=licon1_PDIFF $count=2 $X=4.385
+ $Y=1.84 $X2=4.585 $Y2=2.4
r124 4 63 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.84 $X2=3.57 $Y2=2.115
r125 4 41 300 $w=1.7e-07 $l=6.95971e-07 $layer=licon1_PDIFF $count=2 $X=3.42
+ $Y=1.84 $X2=3.57 $Y2=2.465
r126 3 59 600 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.84 $X2=2.28 $Y2=2.145
r127 3 36 300 $w=1.7e-07 $l=7.48348e-07 $layer=licon1_PDIFF $count=2 $X=2.08
+ $Y=1.84 $X2=2.28 $Y2=2.495
r128 2 29 300 $w=1.7e-07 $l=5.20481e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.84 $X2=1.28 $Y2=2.27
r129 1 24 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r130 1 21 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__A32OI_2%Y 1 2 3 4 13 15 17 23 25 27 29 34 38 42 43
+ 44 47 50
c80 44 0 1.39445e-19 $X=3.035 $Y=1.58
c81 43 0 5.89156e-20 $X=3.12 $Y=1.235
c82 25 0 8.87788e-21 $X=3.005 $Y=0.925
r83 47 50 2.75584 $w=2.28e-07 $l=5.5e-08 $layer=LI1_cond $X=3.12 $Y=1.72
+ $X2=3.12 $Y2=1.665
r84 44 47 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=1.805 $X2=3.12
+ $Y2=1.72
r85 44 50 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.12 $Y=1.65
+ $X2=3.12 $Y2=1.665
r86 42 44 15.0319 $w=2.28e-07 $l=3e-07 $layer=LI1_cond $X=3.12 $Y=1.35 $X2=3.12
+ $Y2=1.65
r87 42 43 5.98911 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.35
+ $X2=3.12 $Y2=1.235
r88 40 41 10.3763 $w=1.94e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=0.76
+ $X2=3.105 $Y2=0.925
r89 34 36 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.62 $Y=0.8
+ $X2=1.62 $Y2=0.925
r90 29 41 5.185 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=1.01 $X2=3.105
+ $Y2=0.925
r91 29 43 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=3.105 $Y=1.01
+ $X2=3.105 $Y2=1.235
r92 28 38 8.61065 $w=1.7e-07 $l=1.83916e-07 $layer=LI1_cond $X=1.945 $Y=1.805
+ $X2=1.78 $Y2=1.845
r93 27 44 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.005 $Y=1.805
+ $X2=3.12 $Y2=1.805
r94 27 28 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=3.005 $Y=1.805
+ $X2=1.945 $Y2=1.805
r95 26 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0.925
+ $X2=1.62 $Y2=0.925
r96 25 41 1.50975 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.005 $Y=0.925
+ $X2=3.105 $Y2=0.925
r97 25 26 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=3.005 $Y=0.925
+ $X2=1.785 $Y2=0.925
r98 21 38 0.89609 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=1.78 $Y=1.97
+ $X2=1.78 $Y2=1.845
r99 21 23 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.78 $Y=1.97
+ $X2=1.78 $Y2=2.65
r100 18 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=1.885
+ $X2=0.78 $Y2=1.885
r101 17 38 8.61065 $w=1.7e-07 $l=1.83916e-07 $layer=LI1_cond $X=1.615 $Y=1.885
+ $X2=1.78 $Y2=1.845
r102 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=1.885
+ $X2=0.945 $Y2=1.885
r103 13 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=1.97 $X2=0.78
+ $Y2=1.885
r104 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.78 $Y=1.97
+ $X2=0.78 $Y2=2.645
r105 4 23 400 $w=1.7e-07 $l=9.04489e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.78 $Y2=2.65
r106 4 21 400 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.78 $Y2=1.97
r107 3 32 400 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.78 $Y2=1.965
r108 3 15 400 $w=1.7e-07 $l=8.97218e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.78 $Y2=2.645
r109 2 40 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=2.97
+ $Y=0.37 $X2=3.11 $Y2=0.76
r110 1 34 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=1.48
+ $Y=0.37 $X2=1.62 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LS__A32OI_2%VPWR 1 2 3 12 16 20 25 26 27 29 34 44 45 48
+ 53
r69 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r70 48 51 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r71 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r72 42 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r73 42 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r74 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r75 39 53 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=4.25 $Y=3.33
+ $X2=4.077 $Y2=3.33
r76 39 41 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.25 $Y=3.33
+ $X2=5.04 $Y2=3.33
r77 38 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r78 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r79 35 48 13.764 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=3.28 $Y=3.33
+ $X2=2.925 $Y2=3.33
r80 35 37 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.28 $Y=3.33 $X2=3.6
+ $Y2=3.33
r81 34 53 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=4.077 $Y2=3.33
r82 34 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=3.6 $Y2=3.33
r83 32 51 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.64 $Y2=3.33
r84 31 32 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r85 29 48 13.764 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=2.57 $Y=3.33
+ $X2=2.925 $Y2=3.33
r86 29 31 152.011 $w=1.68e-07 $l=2.33e-06 $layer=LI1_cond $X=2.57 $Y=3.33
+ $X2=0.24 $Y2=3.33
r87 27 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r88 27 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r89 27 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r90 25 41 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.045 $Y=3.33
+ $X2=5.04 $Y2=3.33
r91 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=3.33
+ $X2=5.21 $Y2=3.33
r92 24 44 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=5.375 $Y=3.33 $X2=6
+ $Y2=3.33
r93 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.375 $Y=3.33
+ $X2=5.21 $Y2=3.33
r94 20 23 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.21 $Y=2.155
+ $X2=5.21 $Y2=2.835
r95 18 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.21 $Y=3.245
+ $X2=5.21 $Y2=3.33
r96 18 23 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.21 $Y=3.245
+ $X2=5.21 $Y2=2.835
r97 14 53 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.077 $Y=3.245
+ $X2=4.077 $Y2=3.33
r98 14 16 29.0616 $w=3.43e-07 $l=8.7e-07 $layer=LI1_cond $X=4.077 $Y=3.245
+ $X2=4.077 $Y2=2.375
r99 10 48 2.89202 $w=7.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=3.245
+ $X2=2.925 $Y2=3.33
r100 10 12 12.6346 $w=7.08e-07 $l=7.5e-07 $layer=LI1_cond $X=2.925 $Y=3.245
+ $X2=2.925 $Y2=2.495
r101 3 23 400 $w=1.7e-07 $l=1.09042e-06 $layer=licon1_PDIFF $count=1 $X=5.01
+ $Y=1.84 $X2=5.21 $Y2=2.835
r102 3 20 400 $w=1.7e-07 $l=4.02772e-07 $layer=licon1_PDIFF $count=1 $X=5.01
+ $Y=1.84 $X2=5.21 $Y2=2.155
r103 2 16 300 $w=1.7e-07 $l=6.29206e-07 $layer=licon1_PDIFF $count=2 $X=3.87
+ $Y=1.84 $X2=4.075 $Y2=2.375
r104 1 12 150 $w=1.7e-07 $l=8.82865e-07 $layer=licon1_PDIFF $count=4 $X=2.58
+ $Y=1.84 $X2=3.115 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LS__A32OI_2%A_27_74# 1 2 3 12 14 15 20 21 22
r37 22 25 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.12 $Y=0.34
+ $X2=2.12 $Y2=0.55
r38 20 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=0.34
+ $X2=2.12 $Y2=0.34
r39 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.955 $Y=0.34
+ $X2=1.275 $Y2=0.34
r40 17 19 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.19 $Y=0.96
+ $X2=1.19 $Y2=0.515
r41 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.19 $Y=0.425
+ $X2=1.275 $Y2=0.34
r42 16 19 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.19 $Y=0.425 $X2=1.19
+ $Y2=0.515
r43 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.105 $Y=1.045
+ $X2=1.19 $Y2=0.96
r44 14 15 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.105 $Y=1.045
+ $X2=0.365 $Y2=1.045
r45 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.365 $Y2=1.045
r46 10 12 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.24 $Y2=0.515
r47 3 25 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=1.91
+ $Y=0.37 $X2=2.12 $Y2=0.55
r48 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.05
+ $Y=0.37 $X2=1.19 $Y2=0.515
r49 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__A32OI_2%VGND 1 2 3 12 16 18 20 22 24 29 37 43 46 50
r67 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r68 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r69 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r70 41 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r71 41 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r72 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r73 38 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.185 $Y=0 $X2=5.06
+ $Y2=0
r74 38 40 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.185 $Y=0 $X2=5.52
+ $Y2=0
r75 37 49 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.795 $Y=0 $X2=6.017
+ $Y2=0
r76 37 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.795 $Y=0 $X2=5.52
+ $Y2=0
r77 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r78 35 36 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r79 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r80 32 35 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.56
+ $Y2=0
r81 32 33 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r82 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r83 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r84 29 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.935 $Y=0 $X2=5.06
+ $Y2=0
r85 29 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.935 $Y=0 $X2=4.56
+ $Y2=0
r86 27 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r87 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r88 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r89 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r90 22 36 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r91 22 33 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=1.2
+ $Y2=0
r92 18 49 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.96 $Y=0.085
+ $X2=6.017 $Y2=0
r93 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.96 $Y=0.085
+ $X2=5.96 $Y2=0.515
r94 14 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.06 $Y=0.085
+ $X2=5.06 $Y2=0
r95 14 16 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=5.06 $Y=0.085
+ $X2=5.06 $Y2=0.675
r96 10 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r97 10 12 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.625
r98 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.82
+ $Y=0.37 $X2=5.96 $Y2=0.515
r99 2 16 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.37 $X2=5.1 $Y2=0.675
r100 1 12 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_LS__A32OI_2%A_507_74# 1 2 3 10 14 16 20 22 27
r44 22 25 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.68 $Y=0.34
+ $X2=2.68 $Y2=0.55
r45 18 20 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=4.54 $Y=0.425
+ $X2=4.54 $Y2=0.675
r46 17 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=0.34
+ $X2=3.54 $Y2=0.34
r47 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.375 $Y=0.34
+ $X2=4.54 $Y2=0.425
r48 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.375 $Y=0.34
+ $X2=3.705 $Y2=0.34
r49 12 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=0.425
+ $X2=3.54 $Y2=0.34
r50 12 14 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.54 $Y=0.425 $X2=3.54
+ $Y2=0.515
r51 11 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=0.34
+ $X2=2.68 $Y2=0.34
r52 10 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=0.34
+ $X2=3.54 $Y2=0.34
r53 10 11 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.375 $Y=0.34
+ $X2=2.845 $Y2=0.34
r54 3 20 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=4.4
+ $Y=0.37 $X2=4.54 $Y2=0.675
r55 2 14 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.4
+ $Y=0.37 $X2=3.54 $Y2=0.515
r56 1 25 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.37 $X2=2.68 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LS__A32OI_2%A_771_74# 1 2 9 11 12 15
r28 13 15 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=5.49 $Y=1.01
+ $X2=5.49 $Y2=0.515
r29 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.365 $Y=1.095
+ $X2=5.49 $Y2=1.01
r30 11 12 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=5.365 $Y=1.095
+ $X2=4.205 $Y2=1.095
r31 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.04 $Y=1.01
+ $X2=4.205 $Y2=1.095
r32 7 9 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=4.04 $Y=1.01 $X2=4.04
+ $Y2=0.76
r33 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.39
+ $Y=0.37 $X2=5.53 $Y2=0.515
r34 1 9 182 $w=1.7e-07 $l=4.7355e-07 $layer=licon1_NDIFF $count=1 $X=3.855
+ $Y=0.37 $X2=4.04 $Y2=0.76
.ends

