* NGSPICE file created from sky130_fd_sc_ls__and4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__and4b_2 A_N B C D VGND VNB VPB VPWR X
M1000 a_537_74# C a_459_74# VNB nshort w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=1.776e+11p ps=1.96e+06u
M1001 a_459_74# D VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=7.2205e+11p ps=4.95e+06u
M1002 a_186_48# D VPWR VPB phighvt w=1e+06u l=150000u
+  ad=6.65e+11p pd=5.33e+06u as=1.86225e+12p ps=1.232e+07u
M1003 VGND a_186_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1004 a_645_74# B a_537_74# VNB nshort w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=0p ps=0u
M1005 VGND A_N a_27_112# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1006 a_186_48# B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_186_48# a_27_112# a_645_74# VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 VPWR A_N a_27_112# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1009 X a_186_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1010 VPWR C a_186_48# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_186_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_186_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_27_112# a_186_48# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

