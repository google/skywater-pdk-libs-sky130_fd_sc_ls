* File: sky130_fd_sc_ls__o22a_2.spice
* Created: Wed Sep  2 11:19:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o22a_2.pex.spice"
.subckt sky130_fd_sc_ls__o22a_2  VNB VPB B1 B2 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_X_M1006_d N_A_82_48#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2035 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1008 N_X_M1006_d N_A_82_48#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.19325 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_82_48#_M1002_d N_B1_M1002_g N_A_307_74#_M1002_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1147 AS=0.195 PD=1.05 PS=2.03 NRD=2.424 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1011 N_A_307_74#_M1011_d N_B2_M1011_g N_A_82_48#_M1002_d VNB NSHORT L=0.15
+ W=0.74 AD=0.1295 AS=0.1147 PD=1.09 PS=1.05 NRD=11.34 NRS=2.424 M=1 R=4.93333
+ SA=75000.6 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g N_A_307_74#_M1011_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1007 N_A_307_74#_M1007_d N_A1_M1007_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_A_82_48#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.3 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1003_d N_A_82_48#_M1003_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.369811 AS=0.168 PD=1.88604 PS=1.42 NRD=48.4029 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1001 A_383_384# N_B1_M1001_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1 AD=0.15
+ AS=0.330189 PD=1.3 PS=1.68396 NRD=18.6953 NRS=54.1947 M=1 R=6.66667 SA=75001.5
+ SB=75001.7 A=0.15 P=2.3 MULT=1
MM1004 N_A_82_48#_M1004_d N_B2_M1004_g A_383_384# VPB PHIGHVT L=0.15 W=1 AD=0.18
+ AS=0.15 PD=1.36 PS=1.3 NRD=1.9503 NRS=18.6953 M=1 R=6.66667 SA=75002
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1005 A_575_384# N_A2_M1005_g N_A_82_48#_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.18 PD=1.39 PS=1.36 NRD=27.5603 NRS=13.7703 M=1 R=6.66667
+ SA=75002.5 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g A_575_384# VPB PHIGHVT L=0.15 W=1 AD=0.29
+ AS=0.195 PD=2.58 PS=1.39 NRD=1.9503 NRS=27.5603 M=1 R=6.66667 SA=75003
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ls__o22a_2.pxi.spice"
*
.ends
*
*
