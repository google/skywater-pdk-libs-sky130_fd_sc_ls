* File: sky130_fd_sc_ls__bufbuf_16.pxi.spice
* Created: Wed Sep  2 10:56:57 2020
* 
x_PM_SKY130_FD_SC_LS__BUFBUF_16%A N_A_c_235_n N_A_M1030_g N_A_M1049_g A
+ N_A_c_237_n PM_SKY130_FD_SC_LS__BUFBUF_16%A
x_PM_SKY130_FD_SC_LS__BUFBUF_16%A_27_368# N_A_27_368#_M1049_s
+ N_A_27_368#_M1030_s N_A_27_368#_M1025_g N_A_27_368#_c_278_n
+ N_A_27_368#_M1001_g N_A_27_368#_M1029_g N_A_27_368#_c_279_n
+ N_A_27_368#_M1031_g N_A_27_368#_M1050_g N_A_27_368#_c_280_n
+ N_A_27_368#_M1043_g N_A_27_368#_c_281_n N_A_27_368#_c_282_n
+ N_A_27_368#_c_270_n N_A_27_368#_c_271_n N_A_27_368#_c_272_n
+ N_A_27_368#_c_296_n N_A_27_368#_c_273_n N_A_27_368#_c_274_n
+ N_A_27_368#_c_275_n N_A_27_368#_c_276_n N_A_27_368#_c_277_n
+ PM_SKY130_FD_SC_LS__BUFBUF_16%A_27_368#
x_PM_SKY130_FD_SC_LS__BUFBUF_16%A_203_74# N_A_203_74#_M1025_s
+ N_A_203_74#_M1050_s N_A_203_74#_M1001_d N_A_203_74#_M1043_d
+ N_A_203_74#_M1000_g N_A_203_74#_c_393_n N_A_203_74#_M1005_g
+ N_A_203_74#_M1006_g N_A_203_74#_c_394_n N_A_203_74#_M1016_g
+ N_A_203_74#_c_395_n N_A_203_74#_M1028_g N_A_203_74#_M1023_g
+ N_A_203_74#_M1027_g N_A_203_74#_c_396_n N_A_203_74#_M1032_g
+ N_A_203_74#_c_397_n N_A_203_74#_M1036_g N_A_203_74#_M1041_g
+ N_A_203_74#_c_398_n N_A_203_74#_M1046_g N_A_203_74#_M1048_g
+ N_A_203_74#_c_399_n N_A_203_74#_c_383_n N_A_203_74#_c_384_n
+ N_A_203_74#_c_385_n N_A_203_74#_c_400_n N_A_203_74#_c_401_n
+ N_A_203_74#_c_386_n N_A_203_74#_c_402_n N_A_203_74#_c_387_n
+ N_A_203_74#_c_388_n N_A_203_74#_c_389_n N_A_203_74#_c_390_n
+ N_A_203_74#_c_404_n N_A_203_74#_c_391_n N_A_203_74#_c_392_n
+ PM_SKY130_FD_SC_LS__BUFBUF_16%A_203_74#
x_PM_SKY130_FD_SC_LS__BUFBUF_16%A_588_74# N_A_588_74#_M1000_d
+ N_A_588_74#_M1023_d N_A_588_74#_M1041_d N_A_588_74#_M1005_s
+ N_A_588_74#_M1028_s N_A_588_74#_M1036_s N_A_588_74#_M1002_g
+ N_A_588_74#_c_606_n N_A_588_74#_M1003_g N_A_588_74#_M1004_g
+ N_A_588_74#_c_607_n N_A_588_74#_M1008_g N_A_588_74#_M1007_g
+ N_A_588_74#_c_608_n N_A_588_74#_M1009_g N_A_588_74#_M1011_g
+ N_A_588_74#_c_609_n N_A_588_74#_M1010_g N_A_588_74#_M1012_g
+ N_A_588_74#_c_610_n N_A_588_74#_M1015_g N_A_588_74#_M1013_g
+ N_A_588_74#_c_611_n N_A_588_74#_M1017_g N_A_588_74#_M1014_g
+ N_A_588_74#_c_612_n N_A_588_74#_M1019_g N_A_588_74#_M1018_g
+ N_A_588_74#_c_613_n N_A_588_74#_M1020_g N_A_588_74#_M1021_g
+ N_A_588_74#_c_614_n N_A_588_74#_M1026_g N_A_588_74#_M1022_g
+ N_A_588_74#_c_615_n N_A_588_74#_M1033_g N_A_588_74#_M1024_g
+ N_A_588_74#_c_616_n N_A_588_74#_M1035_g N_A_588_74#_M1034_g
+ N_A_588_74#_c_617_n N_A_588_74#_M1038_g N_A_588_74#_M1037_g
+ N_A_588_74#_c_618_n N_A_588_74#_M1039_g N_A_588_74#_M1040_g
+ N_A_588_74#_c_619_n N_A_588_74#_M1044_g N_A_588_74#_c_620_n
+ N_A_588_74#_M1047_g N_A_588_74#_M1042_g N_A_588_74#_M1045_g
+ N_A_588_74#_c_621_n N_A_588_74#_M1051_g N_A_588_74#_c_587_n
+ N_A_588_74#_c_622_n N_A_588_74#_c_623_n N_A_588_74#_c_588_n
+ N_A_588_74#_c_589_n N_A_588_74#_c_624_n N_A_588_74#_c_625_n
+ N_A_588_74#_c_590_n N_A_588_74#_c_591_n N_A_588_74#_c_626_n
+ N_A_588_74#_c_592_n N_A_588_74#_c_628_n N_A_588_74#_c_593_n
+ N_A_588_74#_c_594_n N_A_588_74#_c_629_n N_A_588_74#_c_595_n
+ N_A_588_74#_c_596_n N_A_588_74#_c_597_n N_A_588_74#_c_598_n
+ N_A_588_74#_c_599_n N_A_588_74#_c_600_n N_A_588_74#_c_601_n
+ N_A_588_74#_c_602_n N_A_588_74#_c_603_n N_A_588_74#_c_604_n
+ N_A_588_74#_c_605_n PM_SKY130_FD_SC_LS__BUFBUF_16%A_588_74#
x_PM_SKY130_FD_SC_LS__BUFBUF_16%VPWR N_VPWR_M1030_d N_VPWR_M1031_s
+ N_VPWR_M1005_d N_VPWR_M1016_d N_VPWR_M1032_d N_VPWR_M1046_d N_VPWR_M1008_s
+ N_VPWR_M1010_s N_VPWR_M1017_s N_VPWR_M1020_s N_VPWR_M1033_s N_VPWR_M1038_s
+ N_VPWR_M1044_s N_VPWR_M1051_s N_VPWR_c_1054_n N_VPWR_c_1055_n N_VPWR_c_1056_n
+ N_VPWR_c_1057_n N_VPWR_c_1058_n N_VPWR_c_1059_n N_VPWR_c_1060_n
+ N_VPWR_c_1061_n N_VPWR_c_1062_n N_VPWR_c_1063_n N_VPWR_c_1064_n
+ N_VPWR_c_1065_n N_VPWR_c_1066_n N_VPWR_c_1067_n N_VPWR_c_1068_n
+ N_VPWR_c_1069_n N_VPWR_c_1070_n N_VPWR_c_1071_n N_VPWR_c_1072_n
+ N_VPWR_c_1073_n N_VPWR_c_1074_n N_VPWR_c_1075_n N_VPWR_c_1076_n
+ N_VPWR_c_1077_n N_VPWR_c_1078_n N_VPWR_c_1079_n N_VPWR_c_1080_n
+ N_VPWR_c_1081_n N_VPWR_c_1082_n N_VPWR_c_1083_n N_VPWR_c_1084_n
+ N_VPWR_c_1085_n N_VPWR_c_1086_n VPWR N_VPWR_c_1087_n N_VPWR_c_1088_n
+ N_VPWR_c_1089_n N_VPWR_c_1090_n N_VPWR_c_1091_n N_VPWR_c_1092_n
+ N_VPWR_c_1093_n N_VPWR_c_1094_n N_VPWR_c_1053_n
+ PM_SKY130_FD_SC_LS__BUFBUF_16%VPWR
x_PM_SKY130_FD_SC_LS__BUFBUF_16%X N_X_M1002_s N_X_M1007_s N_X_M1012_s
+ N_X_M1014_s N_X_M1021_s N_X_M1024_s N_X_M1037_s N_X_M1042_s N_X_M1003_d
+ N_X_M1009_d N_X_M1015_d N_X_M1019_d N_X_M1026_d N_X_M1035_d N_X_M1039_d
+ N_X_M1047_d N_X_c_1285_n N_X_c_1296_n N_X_c_1297_n N_X_c_1286_n N_X_c_1298_n
+ N_X_c_1287_n N_X_c_1299_n N_X_c_1288_n N_X_c_1300_n N_X_c_1289_n N_X_c_1301_n
+ N_X_c_1290_n N_X_c_1302_n N_X_c_1291_n N_X_c_1304_n N_X_c_1292_n N_X_c_1293_n
+ N_X_c_1306_n N_X_c_1391_n N_X_c_1393_n N_X_c_1395_n N_X_c_1397_n N_X_c_1399_n
+ N_X_c_1294_n X N_X_c_1403_n N_X_c_1307_n N_X_c_1414_n N_X_c_1308_n
+ N_X_c_1424_n N_X_c_1309_n N_X_c_1434_n N_X_c_1310_n N_X_c_1444_n N_X_c_1311_n
+ N_X_c_1454_n N_X_c_1459_n N_X_c_1461_n PM_SKY130_FD_SC_LS__BUFBUF_16%X
x_PM_SKY130_FD_SC_LS__BUFBUF_16%VGND N_VGND_M1049_d N_VGND_M1029_d
+ N_VGND_M1000_s N_VGND_M1006_s N_VGND_M1027_s N_VGND_M1048_s N_VGND_M1004_d
+ N_VGND_M1011_d N_VGND_M1013_d N_VGND_M1018_d N_VGND_M1022_d N_VGND_M1034_d
+ N_VGND_M1040_d N_VGND_M1045_d N_VGND_c_1568_n N_VGND_c_1569_n N_VGND_c_1570_n
+ N_VGND_c_1571_n N_VGND_c_1572_n N_VGND_c_1573_n N_VGND_c_1574_n
+ N_VGND_c_1575_n N_VGND_c_1576_n N_VGND_c_1577_n N_VGND_c_1578_n
+ N_VGND_c_1579_n N_VGND_c_1580_n N_VGND_c_1581_n N_VGND_c_1582_n
+ N_VGND_c_1583_n N_VGND_c_1584_n N_VGND_c_1585_n N_VGND_c_1586_n
+ N_VGND_c_1587_n N_VGND_c_1588_n N_VGND_c_1589_n N_VGND_c_1590_n
+ N_VGND_c_1591_n N_VGND_c_1592_n N_VGND_c_1593_n N_VGND_c_1594_n
+ N_VGND_c_1595_n N_VGND_c_1596_n VGND N_VGND_c_1597_n N_VGND_c_1598_n
+ N_VGND_c_1599_n N_VGND_c_1600_n N_VGND_c_1601_n N_VGND_c_1602_n
+ N_VGND_c_1603_n N_VGND_c_1604_n N_VGND_c_1605_n N_VGND_c_1606_n
+ N_VGND_c_1607_n N_VGND_c_1608_n N_VGND_c_1609_n N_VGND_c_1610_n
+ PM_SKY130_FD_SC_LS__BUFBUF_16%VGND
cc_1 VNB N_A_c_235_n 0.0469497f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_A_M1049_g 0.0292035f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_3 VNB N_A_c_237_n 0.0164929f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_4 VNB N_A_27_368#_M1025_g 0.0208235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_A_27_368#_M1029_g 0.0203832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_368#_M1050_g 0.0236987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_368#_c_270_n 0.0247745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_368#_c_271_n 0.00328084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_368#_c_272_n 0.00880147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_368#_c_273_n 0.00305978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_368#_c_274_n 4.30494e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_368#_c_275_n 9.89968e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_368#_c_276_n 0.00196276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_368#_c_277_n 0.075733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_203_74#_M1000_g 0.0249724f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.665
cc_16 VNB N_A_203_74#_M1006_g 0.0221345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_203_74#_M1023_g 0.0226903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_203_74#_M1027_g 0.0221052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_203_74#_M1041_g 0.0226392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_203_74#_M1048_g 0.0218922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_203_74#_c_383_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_203_74#_c_384_n 0.00278048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_203_74#_c_385_n 0.00140582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_203_74#_c_386_n 0.00886931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_203_74#_c_387_n 0.00537054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_203_74#_c_388_n 2.51917e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_203_74#_c_389_n 0.0289582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_203_74#_c_390_n 0.00384974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_203_74#_c_391_n 0.00554308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_203_74#_c_392_n 0.153349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_588_74#_M1002_g 0.0218098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_588_74#_M1004_g 0.0214105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_588_74#_M1007_g 0.0221679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_588_74#_M1011_g 0.0221649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_588_74#_M1012_g 0.0221667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_588_74#_M1013_g 0.0221573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_588_74#_M1014_g 0.0221554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_588_74#_M1018_g 0.0230696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_588_74#_M1021_g 0.0221575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_588_74#_M1022_g 0.0223217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_588_74#_M1024_g 0.0221589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_588_74#_M1034_g 0.0223264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_588_74#_M1037_g 0.0230747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_588_74#_M1040_g 0.0224479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_588_74#_M1042_g 0.0229374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_588_74#_M1045_g 0.0275406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_588_74#_c_587_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_588_74#_c_588_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_588_74#_c_589_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_588_74#_c_590_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_588_74#_c_591_n 0.00394887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_588_74#_c_592_n 0.00512973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_588_74#_c_593_n 0.00207939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_588_74#_c_594_n 0.00160381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_588_74#_c_595_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_588_74#_c_596_n 6.82873e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_588_74#_c_597_n 0.00256367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_588_74#_c_598_n 0.00101348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_588_74#_c_599_n 0.00102104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_588_74#_c_600_n 0.00169752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_588_74#_c_601_n 0.00169308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_588_74#_c_602_n 0.00168836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_588_74#_c_603_n 0.00167714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_588_74#_c_604_n 0.00173951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_588_74#_c_605_n 0.460539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VPWR_c_1053_n 0.541827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_X_c_1285_n 0.00387206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_X_c_1286_n 0.00613809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_X_c_1287_n 0.00430032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_X_c_1288_n 0.00427247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_X_c_1289_n 0.00400922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_X_c_1290_n 0.00403739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_X_c_1291_n 0.00624928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_X_c_1292_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_X_c_1293_n 0.00177005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_X_c_1294_n 8.14549e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1568_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1569_n 0.00487792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1570_n 0.0194176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1571_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1572_n 0.00508214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1573_n 0.00907711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1574_n 0.00610153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1575_n 0.0185633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1576_n 0.00914547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1577_n 0.0191273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1578_n 0.00977395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1579_n 0.0103321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1580_n 0.00733316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1581_n 0.00738619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1582_n 0.00814903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1583_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1584_n 0.0551309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1585_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1586_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1587_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1588_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1589_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1590_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1591_n 0.0193197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1592_n 0.00346226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1593_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1594_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1595_n 0.0172076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1596_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1597_n 0.0178682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1598_n 0.0208471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1599_n 0.0178544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1600_n 0.0174535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1601_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1602_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1603_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1604_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1605_n 0.00413547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1606_n 0.00509721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1607_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1608_n 0.00579171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1609_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1610_n 0.677396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VPB N_A_c_235_n 0.0289679f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_121 VPB N_A_c_237_n 0.0073823f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_122 VPB N_A_27_368#_c_278_n 0.0157325f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_123 VPB N_A_27_368#_c_279_n 0.0152259f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_27_368#_c_280_n 0.0174767f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_27_368#_c_281_n 0.00758177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_27_368#_c_282_n 0.035396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_27_368#_c_274_n 0.00282546f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_27_368#_c_277_n 0.0201051f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_203_74#_c_393_n 0.016706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_203_74#_c_394_n 0.0154142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_203_74#_c_395_n 0.0154142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_203_74#_c_396_n 0.0154714f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_203_74#_c_397_n 0.0154739f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_203_74#_c_398_n 0.015613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_203_74#_c_399_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_203_74#_c_400_n 0.00179527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_203_74#_c_401_n 0.00183475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_203_74#_c_402_n 0.0119925f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_203_74#_c_388_n 0.00389907f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_203_74#_c_404_n 0.00354092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_203_74#_c_392_n 0.0392138f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_588_74#_c_606_n 0.0155965f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_588_74#_c_607_n 0.0158608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_588_74#_c_608_n 0.0156169f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_588_74#_c_609_n 0.0154857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_588_74#_c_610_n 0.0152381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_588_74#_c_611_n 0.0154857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_588_74#_c_612_n 0.0152381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_588_74#_c_613_n 0.0154857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_588_74#_c_614_n 0.0152381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_588_74#_c_615_n 0.0154857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_588_74#_c_616_n 0.0152381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_588_74#_c_617_n 0.0154849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_588_74#_c_618_n 0.015238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_588_74#_c_619_n 0.0154847f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_588_74#_c_620_n 0.0154624f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_588_74#_c_621_n 0.018112f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_588_74#_c_622_n 0.00183525f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_588_74#_c_623_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_588_74#_c_624_n 0.00179576f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_588_74#_c_625_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_588_74#_c_626_n 0.00225253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_588_74#_c_592_n 0.00383306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_588_74#_c_628_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_588_74#_c_629_n 0.00183525f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_588_74#_c_597_n 0.0203553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_588_74#_c_598_n 0.00140185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_588_74#_c_599_n 0.001404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_588_74#_c_600_n 0.001404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_588_74#_c_601_n 0.00146853f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_588_74#_c_602_n 0.00153061f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_588_74#_c_603_n 0.00193852f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_588_74#_c_604_n 0.00154468f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_588_74#_c_605_n 0.0968951f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1054_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1055_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1056_n 0.0224094f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1057_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1058_n 0.00799791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1059_n 0.00799791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1060_n 0.00886117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1061_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1062_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1063_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1064_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1065_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1066_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1067_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1068_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1069_n 0.0108116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1070_n 0.0645842f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1071_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1072_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1073_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1074_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1075_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1076_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1077_n 0.0209223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1078_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1079_n 0.0199677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1080_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1081_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1082_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1083_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1084_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1085_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1086_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1087_n 0.0220361f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1088_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1089_n 0.0194914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1090_n 0.0233502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1091_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1092_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1093_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1094_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1053_n 0.155444f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_X_c_1285_n 6.16092e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_X_c_1296_n 6.42544e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_X_c_1297_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_X_c_1298_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_X_c_1299_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_X_c_1300_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_X_c_1301_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_X_c_1302_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_X_c_1291_n 0.00126227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_X_c_1304_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_X_c_1293_n 0.0028678f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_X_c_1306_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_X_c_1307_n 0.0012582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_X_c_1308_n 0.0012582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_X_c_1309_n 0.0012582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_X_c_1310_n 0.0012582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_X_c_1311_n 0.00125958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 N_A_M1049_g N_A_27_368#_M1025_g 0.0271299f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A_c_235_n N_A_27_368#_c_278_n 0.0214583f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_236 N_A_c_235_n N_A_27_368#_c_281_n 0.0016558f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A_c_237_n N_A_27_368#_c_281_n 0.0258609f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_238 N_A_c_235_n N_A_27_368#_c_282_n 0.0104891f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A_M1049_g N_A_27_368#_c_270_n 0.00159319f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A_c_235_n N_A_27_368#_c_271_n 7.76566e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A_M1049_g N_A_27_368#_c_271_n 0.0147297f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A_c_237_n N_A_27_368#_c_271_n 0.00934403f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_243 N_A_c_235_n N_A_27_368#_c_272_n 0.00162252f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_244 N_A_c_237_n N_A_27_368#_c_272_n 0.0219376f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_245 N_A_c_235_n N_A_27_368#_c_296_n 0.0139266f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_246 N_A_c_237_n N_A_27_368#_c_296_n 0.00433199f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_247 N_A_M1049_g N_A_27_368#_c_273_n 0.00383985f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A_c_235_n N_A_27_368#_c_274_n 0.0048739f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_249 N_A_c_237_n N_A_27_368#_c_274_n 0.0113191f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_250 N_A_c_235_n N_A_27_368#_c_276_n 0.00282733f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_251 N_A_c_237_n N_A_27_368#_c_276_n 0.0280981f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_252 N_A_c_235_n N_A_27_368#_c_277_n 0.0201541f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_253 N_A_c_237_n N_A_27_368#_c_277_n 3.07734e-19 $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_254 N_A_c_235_n N_A_203_74#_c_399_n 7.53836e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_255 N_A_c_235_n N_VPWR_c_1054_n 0.00486623f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_256 N_A_c_235_n N_VPWR_c_1090_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_257 N_A_c_235_n N_VPWR_c_1053_n 0.00861168f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_258 N_A_M1049_g N_VGND_c_1568_n 0.0125189f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A_M1049_g N_VGND_c_1597_n 0.00383152f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A_M1049_g N_VGND_c_1610_n 0.00761248f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_27_368#_c_278_n N_A_203_74#_c_399_n 0.0123949f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_262 N_A_27_368#_c_279_n N_A_203_74#_c_399_n 0.0125029f $X=1.405 $Y=1.765
+ $X2=0 $Y2=0
cc_263 N_A_27_368#_c_280_n N_A_203_74#_c_399_n 6.9119e-19 $X=1.855 $Y=1.765
+ $X2=0 $Y2=0
cc_264 N_A_27_368#_c_282_n N_A_203_74#_c_399_n 0.00469517f $X=0.28 $Y=2.815
+ $X2=0 $Y2=0
cc_265 N_A_27_368#_M1025_g N_A_203_74#_c_383_n 3.92313e-19 $X=0.94 $Y=0.74 $X2=0
+ $Y2=0
cc_266 N_A_27_368#_M1029_g N_A_203_74#_c_383_n 3.92313e-19 $X=1.37 $Y=0.74 $X2=0
+ $Y2=0
cc_267 N_A_27_368#_M1029_g N_A_203_74#_c_384_n 0.0124689f $X=1.37 $Y=0.74 $X2=0
+ $Y2=0
cc_268 N_A_27_368#_M1050_g N_A_203_74#_c_384_n 0.0111329f $X=1.805 $Y=0.74 $X2=0
+ $Y2=0
cc_269 N_A_27_368#_c_275_n N_A_203_74#_c_384_n 0.045124f $X=1.71 $Y=1.465 $X2=0
+ $Y2=0
cc_270 N_A_27_368#_c_277_n N_A_203_74#_c_384_n 0.00235416f $X=1.805 $Y=1.532
+ $X2=0 $Y2=0
cc_271 N_A_27_368#_c_271_n N_A_203_74#_c_385_n 0.00146386f $X=0.675 $Y=1.045
+ $X2=0 $Y2=0
cc_272 N_A_27_368#_c_275_n N_A_203_74#_c_385_n 0.0143381f $X=1.71 $Y=1.465 $X2=0
+ $Y2=0
cc_273 N_A_27_368#_c_277_n N_A_203_74#_c_385_n 0.00232957f $X=1.805 $Y=1.532
+ $X2=0 $Y2=0
cc_274 N_A_27_368#_c_279_n N_A_203_74#_c_400_n 0.0120074f $X=1.405 $Y=1.765
+ $X2=0 $Y2=0
cc_275 N_A_27_368#_c_280_n N_A_203_74#_c_400_n 0.0124959f $X=1.855 $Y=1.765
+ $X2=0 $Y2=0
cc_276 N_A_27_368#_c_275_n N_A_203_74#_c_400_n 0.0389377f $X=1.71 $Y=1.465 $X2=0
+ $Y2=0
cc_277 N_A_27_368#_c_277_n N_A_203_74#_c_400_n 0.00763082f $X=1.805 $Y=1.532
+ $X2=0 $Y2=0
cc_278 N_A_27_368#_c_278_n N_A_203_74#_c_401_n 0.00232081f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_279 N_A_27_368#_c_279_n N_A_203_74#_c_401_n 9.3899e-19 $X=1.405 $Y=1.765
+ $X2=0 $Y2=0
cc_280 N_A_27_368#_c_274_n N_A_203_74#_c_401_n 0.00779207f $X=0.76 $Y=1.95 $X2=0
+ $Y2=0
cc_281 N_A_27_368#_c_275_n N_A_203_74#_c_401_n 0.0276943f $X=1.71 $Y=1.465 $X2=0
+ $Y2=0
cc_282 N_A_27_368#_c_277_n N_A_203_74#_c_401_n 0.00792231f $X=1.805 $Y=1.532
+ $X2=0 $Y2=0
cc_283 N_A_27_368#_M1029_g N_A_203_74#_c_386_n 6.2115e-19 $X=1.37 $Y=0.74 $X2=0
+ $Y2=0
cc_284 N_A_27_368#_M1050_g N_A_203_74#_c_386_n 0.00965297f $X=1.805 $Y=0.74
+ $X2=0 $Y2=0
cc_285 N_A_27_368#_c_279_n N_A_203_74#_c_402_n 6.9119e-19 $X=1.405 $Y=1.765
+ $X2=0 $Y2=0
cc_286 N_A_27_368#_c_280_n N_A_203_74#_c_402_n 0.013033f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_287 N_A_27_368#_M1050_g N_A_203_74#_c_387_n 0.00581735f $X=1.805 $Y=0.74
+ $X2=0 $Y2=0
cc_288 N_A_27_368#_c_275_n N_A_203_74#_c_387_n 0.00148049f $X=1.71 $Y=1.465
+ $X2=0 $Y2=0
cc_289 N_A_27_368#_c_277_n N_A_203_74#_c_387_n 5.85517e-19 $X=1.805 $Y=1.532
+ $X2=0 $Y2=0
cc_290 N_A_27_368#_c_280_n N_A_203_74#_c_388_n 0.00125956f $X=1.855 $Y=1.765
+ $X2=0 $Y2=0
cc_291 N_A_27_368#_c_277_n N_A_203_74#_c_388_n 0.00440021f $X=1.805 $Y=1.532
+ $X2=0 $Y2=0
cc_292 N_A_27_368#_M1050_g N_A_203_74#_c_390_n 0.00121029f $X=1.805 $Y=0.74
+ $X2=0 $Y2=0
cc_293 N_A_27_368#_c_275_n N_A_203_74#_c_390_n 0.00159649f $X=1.71 $Y=1.465
+ $X2=0 $Y2=0
cc_294 N_A_27_368#_c_277_n N_A_203_74#_c_390_n 0.00218305f $X=1.805 $Y=1.532
+ $X2=0 $Y2=0
cc_295 N_A_27_368#_c_280_n N_A_203_74#_c_404_n 0.00140967f $X=1.855 $Y=1.765
+ $X2=0 $Y2=0
cc_296 N_A_27_368#_c_277_n N_A_203_74#_c_404_n 5.72167e-19 $X=1.805 $Y=1.532
+ $X2=0 $Y2=0
cc_297 N_A_27_368#_c_275_n N_A_203_74#_c_391_n 0.0275462f $X=1.71 $Y=1.465 $X2=0
+ $Y2=0
cc_298 N_A_27_368#_c_277_n N_A_203_74#_c_391_n 0.0101009f $X=1.805 $Y=1.532
+ $X2=0 $Y2=0
cc_299 N_A_27_368#_c_296_n N_VPWR_M1030_d 0.00457874f $X=0.675 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_300 N_A_27_368#_c_274_n N_VPWR_M1030_d 0.0015936f $X=0.76 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_301 N_A_27_368#_c_278_n N_VPWR_c_1054_n 0.00486623f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_A_27_368#_c_282_n N_VPWR_c_1054_n 0.0449718f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_303 N_A_27_368#_c_296_n N_VPWR_c_1054_n 0.0148103f $X=0.675 $Y=2.035 $X2=0
+ $Y2=0
cc_304 N_A_27_368#_c_279_n N_VPWR_c_1055_n 0.00586501f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_305 N_A_27_368#_c_280_n N_VPWR_c_1055_n 0.00586501f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_306 N_A_27_368#_c_280_n N_VPWR_c_1056_n 0.0046855f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_307 N_A_27_368#_c_278_n N_VPWR_c_1071_n 0.00445602f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_308 N_A_27_368#_c_279_n N_VPWR_c_1071_n 0.00445602f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_309 N_A_27_368#_c_280_n N_VPWR_c_1087_n 0.00445602f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_310 N_A_27_368#_c_282_n N_VPWR_c_1090_n 0.0145938f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_311 N_A_27_368#_c_278_n N_VPWR_c_1053_n 0.00857673f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_312 N_A_27_368#_c_279_n N_VPWR_c_1053_n 0.00857589f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_313 N_A_27_368#_c_280_n N_VPWR_c_1053_n 0.00862391f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_314 N_A_27_368#_c_282_n N_VPWR_c_1053_n 0.0120466f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_315 N_A_27_368#_c_271_n N_VGND_M1049_d 0.00214519f $X=0.675 $Y=1.045
+ $X2=-0.19 $Y2=-0.245
cc_316 N_A_27_368#_M1025_g N_VGND_c_1568_n 0.00978365f $X=0.94 $Y=0.74 $X2=0
+ $Y2=0
cc_317 N_A_27_368#_M1029_g N_VGND_c_1568_n 4.56715e-19 $X=1.37 $Y=0.74 $X2=0
+ $Y2=0
cc_318 N_A_27_368#_c_270_n N_VGND_c_1568_n 0.0164982f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_319 N_A_27_368#_c_271_n N_VGND_c_1568_n 0.016426f $X=0.675 $Y=1.045 $X2=0
+ $Y2=0
cc_320 N_A_27_368#_c_275_n N_VGND_c_1568_n 0.00113213f $X=1.71 $Y=1.465 $X2=0
+ $Y2=0
cc_321 N_A_27_368#_M1025_g N_VGND_c_1569_n 4.57991e-19 $X=0.94 $Y=0.74 $X2=0
+ $Y2=0
cc_322 N_A_27_368#_M1029_g N_VGND_c_1569_n 0.0090301f $X=1.37 $Y=0.74 $X2=0
+ $Y2=0
cc_323 N_A_27_368#_M1050_g N_VGND_c_1569_n 0.00455924f $X=1.805 $Y=0.74 $X2=0
+ $Y2=0
cc_324 N_A_27_368#_M1050_g N_VGND_c_1570_n 0.00414085f $X=1.805 $Y=0.74 $X2=0
+ $Y2=0
cc_325 N_A_27_368#_M1025_g N_VGND_c_1585_n 0.00383152f $X=0.94 $Y=0.74 $X2=0
+ $Y2=0
cc_326 N_A_27_368#_M1029_g N_VGND_c_1585_n 0.00383152f $X=1.37 $Y=0.74 $X2=0
+ $Y2=0
cc_327 N_A_27_368#_c_270_n N_VGND_c_1597_n 0.011066f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_328 N_A_27_368#_M1050_g N_VGND_c_1598_n 0.00434272f $X=1.805 $Y=0.74 $X2=0
+ $Y2=0
cc_329 N_A_27_368#_M1025_g N_VGND_c_1610_n 0.0075754f $X=0.94 $Y=0.74 $X2=0
+ $Y2=0
cc_330 N_A_27_368#_M1029_g N_VGND_c_1610_n 0.0075754f $X=1.37 $Y=0.74 $X2=0
+ $Y2=0
cc_331 N_A_27_368#_M1050_g N_VGND_c_1610_n 0.00825445f $X=1.805 $Y=0.74 $X2=0
+ $Y2=0
cc_332 N_A_27_368#_c_270_n N_VGND_c_1610_n 0.00915947f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_333 N_A_203_74#_M1048_g N_A_588_74#_M1002_g 0.0171756f $X=5.155 $Y=0.74 $X2=0
+ $Y2=0
cc_334 N_A_203_74#_c_398_n N_A_588_74#_c_606_n 0.00875024f $X=5.14 $Y=1.765
+ $X2=0 $Y2=0
cc_335 N_A_203_74#_M1000_g N_A_588_74#_c_587_n 0.00765982f $X=2.865 $Y=0.74
+ $X2=0 $Y2=0
cc_336 N_A_203_74#_M1006_g N_A_588_74#_c_587_n 3.97481e-19 $X=3.295 $Y=0.74
+ $X2=0 $Y2=0
cc_337 N_A_203_74#_c_393_n N_A_588_74#_c_622_n 0.0022934f $X=2.88 $Y=1.765 $X2=0
+ $Y2=0
cc_338 N_A_203_74#_c_394_n N_A_588_74#_c_622_n 6.83942e-19 $X=3.33 $Y=1.765
+ $X2=0 $Y2=0
cc_339 N_A_203_74#_c_389_n N_A_588_74#_c_622_n 0.0276944f $X=4.315 $Y=1.485
+ $X2=0 $Y2=0
cc_340 N_A_203_74#_c_392_n N_A_588_74#_c_622_n 0.00789892f $X=5.14 $Y=1.542
+ $X2=0 $Y2=0
cc_341 N_A_203_74#_c_393_n N_A_588_74#_c_623_n 0.0116424f $X=2.88 $Y=1.765 $X2=0
+ $Y2=0
cc_342 N_A_203_74#_c_394_n N_A_588_74#_c_623_n 0.0123f $X=3.33 $Y=1.765 $X2=0
+ $Y2=0
cc_343 N_A_203_74#_c_395_n N_A_588_74#_c_623_n 6.8511e-19 $X=3.78 $Y=1.765 $X2=0
+ $Y2=0
cc_344 N_A_203_74#_M1006_g N_A_588_74#_c_588_n 0.0131239f $X=3.295 $Y=0.74 $X2=0
+ $Y2=0
cc_345 N_A_203_74#_M1023_g N_A_588_74#_c_588_n 0.0114885f $X=3.795 $Y=0.74 $X2=0
+ $Y2=0
cc_346 N_A_203_74#_c_389_n N_A_588_74#_c_588_n 0.0500092f $X=4.315 $Y=1.485
+ $X2=0 $Y2=0
cc_347 N_A_203_74#_c_392_n N_A_588_74#_c_588_n 0.00381149f $X=5.14 $Y=1.542
+ $X2=0 $Y2=0
cc_348 N_A_203_74#_M1000_g N_A_588_74#_c_589_n 0.00337781f $X=2.865 $Y=0.74
+ $X2=0 $Y2=0
cc_349 N_A_203_74#_c_389_n N_A_588_74#_c_589_n 0.0209731f $X=4.315 $Y=1.485
+ $X2=0 $Y2=0
cc_350 N_A_203_74#_c_392_n N_A_588_74#_c_589_n 0.00232957f $X=5.14 $Y=1.542
+ $X2=0 $Y2=0
cc_351 N_A_203_74#_c_394_n N_A_588_74#_c_624_n 0.0120074f $X=3.33 $Y=1.765 $X2=0
+ $Y2=0
cc_352 N_A_203_74#_c_395_n N_A_588_74#_c_624_n 0.0120074f $X=3.78 $Y=1.765 $X2=0
+ $Y2=0
cc_353 N_A_203_74#_c_389_n N_A_588_74#_c_624_n 0.0417603f $X=4.315 $Y=1.485
+ $X2=0 $Y2=0
cc_354 N_A_203_74#_c_392_n N_A_588_74#_c_624_n 0.00735278f $X=5.14 $Y=1.542
+ $X2=0 $Y2=0
cc_355 N_A_203_74#_c_394_n N_A_588_74#_c_625_n 6.8511e-19 $X=3.33 $Y=1.765 $X2=0
+ $Y2=0
cc_356 N_A_203_74#_c_395_n N_A_588_74#_c_625_n 0.0123f $X=3.78 $Y=1.765 $X2=0
+ $Y2=0
cc_357 N_A_203_74#_c_396_n N_A_588_74#_c_625_n 0.0123512f $X=4.23 $Y=1.765 $X2=0
+ $Y2=0
cc_358 N_A_203_74#_c_397_n N_A_588_74#_c_625_n 6.81182e-19 $X=4.69 $Y=1.765
+ $X2=0 $Y2=0
cc_359 N_A_203_74#_M1006_g N_A_588_74#_c_590_n 8.89165e-19 $X=3.295 $Y=0.74
+ $X2=0 $Y2=0
cc_360 N_A_203_74#_M1023_g N_A_588_74#_c_590_n 0.00882909f $X=3.795 $Y=0.74
+ $X2=0 $Y2=0
cc_361 N_A_203_74#_M1027_g N_A_588_74#_c_590_n 3.97481e-19 $X=4.225 $Y=0.74
+ $X2=0 $Y2=0
cc_362 N_A_203_74#_M1027_g N_A_588_74#_c_591_n 0.0131239f $X=4.225 $Y=0.74 $X2=0
+ $Y2=0
cc_363 N_A_203_74#_M1041_g N_A_588_74#_c_591_n 0.0133559f $X=4.725 $Y=0.74 $X2=0
+ $Y2=0
cc_364 N_A_203_74#_c_389_n N_A_588_74#_c_591_n 0.0283384f $X=4.315 $Y=1.485
+ $X2=0 $Y2=0
cc_365 N_A_203_74#_c_392_n N_A_588_74#_c_591_n 0.00420544f $X=5.14 $Y=1.542
+ $X2=0 $Y2=0
cc_366 N_A_203_74#_c_396_n N_A_588_74#_c_626_n 0.012065f $X=4.23 $Y=1.765 $X2=0
+ $Y2=0
cc_367 N_A_203_74#_c_397_n N_A_588_74#_c_626_n 0.0140404f $X=4.69 $Y=1.765 $X2=0
+ $Y2=0
cc_368 N_A_203_74#_c_389_n N_A_588_74#_c_626_n 0.0227591f $X=4.315 $Y=1.485
+ $X2=0 $Y2=0
cc_369 N_A_203_74#_c_392_n N_A_588_74#_c_626_n 0.00829792f $X=5.14 $Y=1.542
+ $X2=0 $Y2=0
cc_370 N_A_203_74#_c_397_n N_A_588_74#_c_592_n 0.00225922f $X=4.69 $Y=1.765
+ $X2=0 $Y2=0
cc_371 N_A_203_74#_c_398_n N_A_588_74#_c_592_n 0.00416027f $X=5.14 $Y=1.765
+ $X2=0 $Y2=0
cc_372 N_A_203_74#_c_389_n N_A_588_74#_c_592_n 0.0147393f $X=4.315 $Y=1.485
+ $X2=0 $Y2=0
cc_373 N_A_203_74#_c_392_n N_A_588_74#_c_592_n 0.050143f $X=5.14 $Y=1.542 $X2=0
+ $Y2=0
cc_374 N_A_203_74#_c_396_n N_A_588_74#_c_628_n 6.92433e-19 $X=4.23 $Y=1.765
+ $X2=0 $Y2=0
cc_375 N_A_203_74#_c_397_n N_A_588_74#_c_628_n 0.0125421f $X=4.69 $Y=1.765 $X2=0
+ $Y2=0
cc_376 N_A_203_74#_c_398_n N_A_588_74#_c_628_n 0.011073f $X=5.14 $Y=1.765 $X2=0
+ $Y2=0
cc_377 N_A_203_74#_M1027_g N_A_588_74#_c_593_n 8.89165e-19 $X=4.225 $Y=0.74
+ $X2=0 $Y2=0
cc_378 N_A_203_74#_M1041_g N_A_588_74#_c_593_n 0.00882909f $X=4.725 $Y=0.74
+ $X2=0 $Y2=0
cc_379 N_A_203_74#_M1048_g N_A_588_74#_c_593_n 4.18373e-19 $X=5.155 $Y=0.74
+ $X2=0 $Y2=0
cc_380 N_A_203_74#_M1041_g N_A_588_74#_c_594_n 0.00440835f $X=4.725 $Y=0.74
+ $X2=0 $Y2=0
cc_381 N_A_203_74#_M1048_g N_A_588_74#_c_594_n 0.00450088f $X=5.155 $Y=0.74
+ $X2=0 $Y2=0
cc_382 N_A_203_74#_c_395_n N_A_588_74#_c_629_n 6.83942e-19 $X=3.78 $Y=1.765
+ $X2=0 $Y2=0
cc_383 N_A_203_74#_c_396_n N_A_588_74#_c_629_n 6.83942e-19 $X=4.23 $Y=1.765
+ $X2=0 $Y2=0
cc_384 N_A_203_74#_c_389_n N_A_588_74#_c_629_n 0.0276944f $X=4.315 $Y=1.485
+ $X2=0 $Y2=0
cc_385 N_A_203_74#_c_392_n N_A_588_74#_c_629_n 0.00789892f $X=5.14 $Y=1.542
+ $X2=0 $Y2=0
cc_386 N_A_203_74#_M1023_g N_A_588_74#_c_595_n 0.00121617f $X=3.795 $Y=0.74
+ $X2=0 $Y2=0
cc_387 N_A_203_74#_c_389_n N_A_588_74#_c_595_n 0.0209731f $X=4.315 $Y=1.485
+ $X2=0 $Y2=0
cc_388 N_A_203_74#_c_392_n N_A_588_74#_c_595_n 0.00232957f $X=5.14 $Y=1.542
+ $X2=0 $Y2=0
cc_389 N_A_203_74#_M1041_g N_A_588_74#_c_596_n 0.00150479f $X=4.725 $Y=0.74
+ $X2=0 $Y2=0
cc_390 N_A_203_74#_M1048_g N_A_588_74#_c_596_n 0.00358809f $X=5.155 $Y=0.74
+ $X2=0 $Y2=0
cc_391 N_A_203_74#_c_398_n N_A_588_74#_c_597_n 0.00472284f $X=5.14 $Y=1.765
+ $X2=0 $Y2=0
cc_392 N_A_203_74#_c_392_n N_A_588_74#_c_597_n 2.6189e-19 $X=5.14 $Y=1.542 $X2=0
+ $Y2=0
cc_393 N_A_203_74#_c_392_n N_A_588_74#_c_605_n 0.0171756f $X=5.14 $Y=1.542 $X2=0
+ $Y2=0
cc_394 N_A_203_74#_c_400_n N_VPWR_M1031_s 0.00247267f $X=1.915 $Y=1.885 $X2=0
+ $Y2=0
cc_395 N_A_203_74#_c_399_n N_VPWR_c_1054_n 0.0449718f $X=1.18 $Y=1.985 $X2=0
+ $Y2=0
cc_396 N_A_203_74#_c_399_n N_VPWR_c_1055_n 0.0547423f $X=1.18 $Y=1.985 $X2=0
+ $Y2=0
cc_397 N_A_203_74#_c_400_n N_VPWR_c_1055_n 0.0136682f $X=1.915 $Y=1.885 $X2=0
+ $Y2=0
cc_398 N_A_203_74#_c_402_n N_VPWR_c_1055_n 0.0547423f $X=2.08 $Y=1.985 $X2=0
+ $Y2=0
cc_399 N_A_203_74#_c_393_n N_VPWR_c_1056_n 0.0100889f $X=2.88 $Y=1.765 $X2=0
+ $Y2=0
cc_400 N_A_203_74#_c_402_n N_VPWR_c_1056_n 0.0638129f $X=2.08 $Y=1.985 $X2=0
+ $Y2=0
cc_401 N_A_203_74#_c_389_n N_VPWR_c_1056_n 0.0219385f $X=4.315 $Y=1.485 $X2=0
+ $Y2=0
cc_402 N_A_203_74#_c_404_n N_VPWR_c_1056_n 0.0100711f $X=2.08 $Y=1.885 $X2=0
+ $Y2=0
cc_403 N_A_203_74#_c_394_n N_VPWR_c_1057_n 0.00571432f $X=3.33 $Y=1.765 $X2=0
+ $Y2=0
cc_404 N_A_203_74#_c_395_n N_VPWR_c_1057_n 0.00571432f $X=3.78 $Y=1.765 $X2=0
+ $Y2=0
cc_405 N_A_203_74#_c_396_n N_VPWR_c_1058_n 0.00574346f $X=4.23 $Y=1.765 $X2=0
+ $Y2=0
cc_406 N_A_203_74#_c_397_n N_VPWR_c_1058_n 0.00575951f $X=4.69 $Y=1.765 $X2=0
+ $Y2=0
cc_407 N_A_203_74#_c_398_n N_VPWR_c_1059_n 0.00603309f $X=5.14 $Y=1.765 $X2=0
+ $Y2=0
cc_408 N_A_203_74#_c_399_n N_VPWR_c_1071_n 0.014552f $X=1.18 $Y=1.985 $X2=0
+ $Y2=0
cc_409 N_A_203_74#_c_393_n N_VPWR_c_1073_n 0.00445602f $X=2.88 $Y=1.765 $X2=0
+ $Y2=0
cc_410 N_A_203_74#_c_394_n N_VPWR_c_1073_n 0.00445602f $X=3.33 $Y=1.765 $X2=0
+ $Y2=0
cc_411 N_A_203_74#_c_395_n N_VPWR_c_1075_n 0.00445602f $X=3.78 $Y=1.765 $X2=0
+ $Y2=0
cc_412 N_A_203_74#_c_396_n N_VPWR_c_1075_n 0.00445602f $X=4.23 $Y=1.765 $X2=0
+ $Y2=0
cc_413 N_A_203_74#_c_397_n N_VPWR_c_1077_n 0.00445602f $X=4.69 $Y=1.765 $X2=0
+ $Y2=0
cc_414 N_A_203_74#_c_398_n N_VPWR_c_1077_n 0.00445602f $X=5.14 $Y=1.765 $X2=0
+ $Y2=0
cc_415 N_A_203_74#_c_402_n N_VPWR_c_1087_n 0.0145938f $X=2.08 $Y=1.985 $X2=0
+ $Y2=0
cc_416 N_A_203_74#_c_393_n N_VPWR_c_1053_n 0.00862391f $X=2.88 $Y=1.765 $X2=0
+ $Y2=0
cc_417 N_A_203_74#_c_394_n N_VPWR_c_1053_n 0.00857589f $X=3.33 $Y=1.765 $X2=0
+ $Y2=0
cc_418 N_A_203_74#_c_395_n N_VPWR_c_1053_n 0.00857589f $X=3.78 $Y=1.765 $X2=0
+ $Y2=0
cc_419 N_A_203_74#_c_396_n N_VPWR_c_1053_n 0.00857685f $X=4.23 $Y=1.765 $X2=0
+ $Y2=0
cc_420 N_A_203_74#_c_397_n N_VPWR_c_1053_n 0.00857909f $X=4.69 $Y=1.765 $X2=0
+ $Y2=0
cc_421 N_A_203_74#_c_398_n N_VPWR_c_1053_n 0.00857762f $X=5.14 $Y=1.765 $X2=0
+ $Y2=0
cc_422 N_A_203_74#_c_399_n N_VPWR_c_1053_n 0.0119791f $X=1.18 $Y=1.985 $X2=0
+ $Y2=0
cc_423 N_A_203_74#_c_402_n N_VPWR_c_1053_n 0.0120466f $X=2.08 $Y=1.985 $X2=0
+ $Y2=0
cc_424 N_A_203_74#_M1048_g N_X_c_1285_n 7.91799e-19 $X=5.155 $Y=0.74 $X2=0 $Y2=0
cc_425 N_A_203_74#_c_392_n N_X_c_1285_n 4.82789e-19 $X=5.14 $Y=1.542 $X2=0 $Y2=0
cc_426 N_A_203_74#_c_398_n N_X_c_1296_n 3.77031e-19 $X=5.14 $Y=1.765 $X2=0 $Y2=0
cc_427 N_A_203_74#_c_384_n N_VGND_M1029_d 0.00177524f $X=1.855 $Y=1.045 $X2=0
+ $Y2=0
cc_428 N_A_203_74#_c_383_n N_VGND_c_1568_n 0.0164567f $X=1.155 $Y=0.515 $X2=0
+ $Y2=0
cc_429 N_A_203_74#_c_383_n N_VGND_c_1569_n 0.0157999f $X=1.155 $Y=0.515 $X2=0
+ $Y2=0
cc_430 N_A_203_74#_c_384_n N_VGND_c_1569_n 0.015373f $X=1.855 $Y=1.045 $X2=0
+ $Y2=0
cc_431 N_A_203_74#_c_386_n N_VGND_c_1569_n 0.0315611f $X=2.02 $Y=0.515 $X2=0
+ $Y2=0
cc_432 N_A_203_74#_M1000_g N_VGND_c_1570_n 0.018401f $X=2.865 $Y=0.74 $X2=0
+ $Y2=0
cc_433 N_A_203_74#_c_386_n N_VGND_c_1570_n 0.0455802f $X=2.02 $Y=0.515 $X2=0
+ $Y2=0
cc_434 N_A_203_74#_c_389_n N_VGND_c_1570_n 0.0268194f $X=4.315 $Y=1.485 $X2=0
+ $Y2=0
cc_435 N_A_203_74#_c_390_n N_VGND_c_1570_n 0.0134079f $X=2.035 $Y=1.045 $X2=0
+ $Y2=0
cc_436 N_A_203_74#_M1000_g N_VGND_c_1571_n 5.08869e-19 $X=2.865 $Y=0.74 $X2=0
+ $Y2=0
cc_437 N_A_203_74#_M1006_g N_VGND_c_1571_n 0.0101377f $X=3.295 $Y=0.74 $X2=0
+ $Y2=0
cc_438 N_A_203_74#_M1023_g N_VGND_c_1571_n 0.00408259f $X=3.795 $Y=0.74 $X2=0
+ $Y2=0
cc_439 N_A_203_74#_M1023_g N_VGND_c_1572_n 5.08869e-19 $X=3.795 $Y=0.74 $X2=0
+ $Y2=0
cc_440 N_A_203_74#_M1027_g N_VGND_c_1572_n 0.0101377f $X=4.225 $Y=0.74 $X2=0
+ $Y2=0
cc_441 N_A_203_74#_M1041_g N_VGND_c_1572_n 0.00417204f $X=4.725 $Y=0.74 $X2=0
+ $Y2=0
cc_442 N_A_203_74#_M1048_g N_VGND_c_1573_n 0.00183296f $X=5.155 $Y=0.74 $X2=0
+ $Y2=0
cc_443 N_A_203_74#_c_383_n N_VGND_c_1585_n 0.00749631f $X=1.155 $Y=0.515 $X2=0
+ $Y2=0
cc_444 N_A_203_74#_M1000_g N_VGND_c_1587_n 0.00434272f $X=2.865 $Y=0.74 $X2=0
+ $Y2=0
cc_445 N_A_203_74#_M1006_g N_VGND_c_1587_n 0.00383152f $X=3.295 $Y=0.74 $X2=0
+ $Y2=0
cc_446 N_A_203_74#_M1023_g N_VGND_c_1589_n 0.00434272f $X=3.795 $Y=0.74 $X2=0
+ $Y2=0
cc_447 N_A_203_74#_M1027_g N_VGND_c_1589_n 0.00383152f $X=4.225 $Y=0.74 $X2=0
+ $Y2=0
cc_448 N_A_203_74#_M1041_g N_VGND_c_1591_n 0.00434272f $X=4.725 $Y=0.74 $X2=0
+ $Y2=0
cc_449 N_A_203_74#_M1048_g N_VGND_c_1591_n 0.00461464f $X=5.155 $Y=0.74 $X2=0
+ $Y2=0
cc_450 N_A_203_74#_c_386_n N_VGND_c_1598_n 0.0159025f $X=2.02 $Y=0.515 $X2=0
+ $Y2=0
cc_451 N_A_203_74#_M1000_g N_VGND_c_1610_n 0.00825059f $X=2.865 $Y=0.74 $X2=0
+ $Y2=0
cc_452 N_A_203_74#_M1006_g N_VGND_c_1610_n 0.0075754f $X=3.295 $Y=0.74 $X2=0
+ $Y2=0
cc_453 N_A_203_74#_M1023_g N_VGND_c_1610_n 0.00820718f $X=3.795 $Y=0.74 $X2=0
+ $Y2=0
cc_454 N_A_203_74#_M1027_g N_VGND_c_1610_n 0.0075754f $X=4.225 $Y=0.74 $X2=0
+ $Y2=0
cc_455 N_A_203_74#_M1041_g N_VGND_c_1610_n 0.00820718f $X=4.725 $Y=0.74 $X2=0
+ $Y2=0
cc_456 N_A_203_74#_M1048_g N_VGND_c_1610_n 0.00908206f $X=5.155 $Y=0.74 $X2=0
+ $Y2=0
cc_457 N_A_203_74#_c_383_n N_VGND_c_1610_n 0.0062048f $X=1.155 $Y=0.515 $X2=0
+ $Y2=0
cc_458 N_A_203_74#_c_386_n N_VGND_c_1610_n 0.0131064f $X=2.02 $Y=0.515 $X2=0
+ $Y2=0
cc_459 N_A_588_74#_c_624_n N_VPWR_M1016_d 0.00247267f $X=3.84 $Y=1.905 $X2=0
+ $Y2=0
cc_460 N_A_588_74#_c_626_n N_VPWR_M1032_d 0.00285423f $X=4.75 $Y=1.905 $X2=0
+ $Y2=0
cc_461 N_A_588_74#_c_622_n N_VPWR_c_1056_n 0.0121319f $X=3.105 $Y=1.99 $X2=0
+ $Y2=0
cc_462 N_A_588_74#_c_623_n N_VPWR_c_1056_n 0.0663772f $X=3.105 $Y=2.815 $X2=0
+ $Y2=0
cc_463 N_A_588_74#_c_623_n N_VPWR_c_1057_n 0.0534396f $X=3.105 $Y=2.815 $X2=0
+ $Y2=0
cc_464 N_A_588_74#_c_624_n N_VPWR_c_1057_n 0.0136682f $X=3.84 $Y=1.905 $X2=0
+ $Y2=0
cc_465 N_A_588_74#_c_625_n N_VPWR_c_1057_n 0.0534396f $X=4.005 $Y=2.815 $X2=0
+ $Y2=0
cc_466 N_A_588_74#_c_625_n N_VPWR_c_1058_n 0.0534396f $X=4.005 $Y=2.815 $X2=0
+ $Y2=0
cc_467 N_A_588_74#_c_626_n N_VPWR_c_1058_n 0.0136682f $X=4.75 $Y=1.905 $X2=0
+ $Y2=0
cc_468 N_A_588_74#_c_628_n N_VPWR_c_1058_n 0.0514755f $X=4.915 $Y=2.815 $X2=0
+ $Y2=0
cc_469 N_A_588_74#_c_606_n N_VPWR_c_1059_n 0.00607438f $X=5.6 $Y=1.765 $X2=0
+ $Y2=0
cc_470 N_A_588_74#_c_592_n N_VPWR_c_1059_n 0.0133926f $X=4.915 $Y=1.99 $X2=0
+ $Y2=0
cc_471 N_A_588_74#_c_628_n N_VPWR_c_1059_n 0.0644799f $X=4.915 $Y=2.815 $X2=0
+ $Y2=0
cc_472 N_A_588_74#_c_597_n N_VPWR_c_1059_n 0.00610188f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_473 N_A_588_74#_c_607_n N_VPWR_c_1060_n 0.00879286f $X=6.05 $Y=1.765 $X2=0
+ $Y2=0
cc_474 N_A_588_74#_c_608_n N_VPWR_c_1060_n 0.00783147f $X=6.55 $Y=1.765 $X2=0
+ $Y2=0
cc_475 N_A_588_74#_c_597_n N_VPWR_c_1060_n 0.00101965f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_476 N_A_588_74#_c_598_n N_VPWR_c_1060_n 0.0139369f $X=6.21 $Y=1.485 $X2=0
+ $Y2=0
cc_477 N_A_588_74#_c_605_n N_VPWR_c_1060_n 0.00225562f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_478 N_A_588_74#_c_609_n N_VPWR_c_1061_n 0.00711256f $X=7 $Y=1.765 $X2=0 $Y2=0
cc_479 N_A_588_74#_c_610_n N_VPWR_c_1061_n 0.00711256f $X=7.45 $Y=1.765 $X2=0
+ $Y2=0
cc_480 N_A_588_74#_c_597_n N_VPWR_c_1061_n 9.65229e-19 $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_481 N_A_588_74#_c_599_n N_VPWR_c_1061_n 0.00513697f $X=7.085 $Y=1.485 $X2=0
+ $Y2=0
cc_482 N_A_588_74#_c_605_n N_VPWR_c_1061_n 0.00295615f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_483 N_A_588_74#_c_611_n N_VPWR_c_1062_n 0.00590719f $X=7.9 $Y=1.765 $X2=0
+ $Y2=0
cc_484 N_A_588_74#_c_612_n N_VPWR_c_1062_n 0.00590719f $X=8.35 $Y=1.765 $X2=0
+ $Y2=0
cc_485 N_A_588_74#_c_597_n N_VPWR_c_1062_n 9.65229e-19 $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_486 N_A_588_74#_c_600_n N_VPWR_c_1062_n 0.00513697f $X=7.985 $Y=1.485 $X2=0
+ $Y2=0
cc_487 N_A_588_74#_c_605_n N_VPWR_c_1062_n 0.00295817f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_488 N_A_588_74#_c_613_n N_VPWR_c_1063_n 0.00590719f $X=8.8 $Y=1.765 $X2=0
+ $Y2=0
cc_489 N_A_588_74#_c_614_n N_VPWR_c_1063_n 0.00590719f $X=9.25 $Y=1.765 $X2=0
+ $Y2=0
cc_490 N_A_588_74#_c_597_n N_VPWR_c_1063_n 8.37589e-19 $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_491 N_A_588_74#_c_601_n N_VPWR_c_1063_n 0.00724805f $X=8.905 $Y=1.485 $X2=0
+ $Y2=0
cc_492 N_A_588_74#_c_605_n N_VPWR_c_1063_n 0.00229926f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_493 N_A_588_74#_c_614_n N_VPWR_c_1064_n 0.00445602f $X=9.25 $Y=1.765 $X2=0
+ $Y2=0
cc_494 N_A_588_74#_c_615_n N_VPWR_c_1064_n 0.00445602f $X=9.7 $Y=1.765 $X2=0
+ $Y2=0
cc_495 N_A_588_74#_c_615_n N_VPWR_c_1065_n 0.00590719f $X=9.7 $Y=1.765 $X2=0
+ $Y2=0
cc_496 N_A_588_74#_c_616_n N_VPWR_c_1065_n 0.00590719f $X=10.15 $Y=1.765 $X2=0
+ $Y2=0
cc_497 N_A_588_74#_c_597_n N_VPWR_c_1065_n 7.09949e-19 $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_498 N_A_588_74#_c_602_n N_VPWR_c_1065_n 0.00935913f $X=9.815 $Y=1.485 $X2=0
+ $Y2=0
cc_499 N_A_588_74#_c_605_n N_VPWR_c_1065_n 0.00164034f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_500 N_A_588_74#_c_616_n N_VPWR_c_1066_n 0.00445602f $X=10.15 $Y=1.765 $X2=0
+ $Y2=0
cc_501 N_A_588_74#_c_617_n N_VPWR_c_1066_n 0.00445602f $X=10.6 $Y=1.765 $X2=0
+ $Y2=0
cc_502 N_A_588_74#_c_617_n N_VPWR_c_1067_n 0.00590719f $X=10.6 $Y=1.765 $X2=0
+ $Y2=0
cc_503 N_A_588_74#_c_618_n N_VPWR_c_1067_n 0.00590719f $X=11.05 $Y=1.765 $X2=0
+ $Y2=0
cc_504 N_A_588_74#_c_597_n N_VPWR_c_1067_n 5.61035e-19 $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_505 N_A_588_74#_c_603_n N_VPWR_c_1067_n 0.0118221f $X=10.76 $Y=1.485 $X2=0
+ $Y2=0
cc_506 N_A_588_74#_c_605_n N_VPWR_c_1067_n 8.71254e-19 $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_507 N_A_588_74#_c_619_n N_VPWR_c_1068_n 0.00637352f $X=11.5 $Y=1.765 $X2=0
+ $Y2=0
cc_508 N_A_588_74#_c_620_n N_VPWR_c_1068_n 0.0129659f $X=11.95 $Y=1.765 $X2=0
+ $Y2=0
cc_509 N_A_588_74#_c_621_n N_VPWR_c_1068_n 8.16443e-19 $X=12.45 $Y=1.765 $X2=0
+ $Y2=0
cc_510 N_A_588_74#_c_597_n N_VPWR_c_1068_n 6.31165e-19 $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_511 N_A_588_74#_c_604_n N_VPWR_c_1068_n 0.0163224f $X=11.685 $Y=1.485 $X2=0
+ $Y2=0
cc_512 N_A_588_74#_c_605_n N_VPWR_c_1068_n 0.00148663f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_513 N_A_588_74#_c_621_n N_VPWR_c_1070_n 0.0102292f $X=12.45 $Y=1.765 $X2=0
+ $Y2=0
cc_514 N_A_588_74#_c_623_n N_VPWR_c_1073_n 0.014552f $X=3.105 $Y=2.815 $X2=0
+ $Y2=0
cc_515 N_A_588_74#_c_625_n N_VPWR_c_1075_n 0.014552f $X=4.005 $Y=2.815 $X2=0
+ $Y2=0
cc_516 N_A_588_74#_c_628_n N_VPWR_c_1077_n 0.014552f $X=4.915 $Y=2.815 $X2=0
+ $Y2=0
cc_517 N_A_588_74#_c_606_n N_VPWR_c_1079_n 0.00445602f $X=5.6 $Y=1.765 $X2=0
+ $Y2=0
cc_518 N_A_588_74#_c_607_n N_VPWR_c_1079_n 0.00445602f $X=6.05 $Y=1.765 $X2=0
+ $Y2=0
cc_519 N_A_588_74#_c_608_n N_VPWR_c_1081_n 0.00445602f $X=6.55 $Y=1.765 $X2=0
+ $Y2=0
cc_520 N_A_588_74#_c_609_n N_VPWR_c_1081_n 0.00445602f $X=7 $Y=1.765 $X2=0 $Y2=0
cc_521 N_A_588_74#_c_610_n N_VPWR_c_1083_n 0.00445602f $X=7.45 $Y=1.765 $X2=0
+ $Y2=0
cc_522 N_A_588_74#_c_611_n N_VPWR_c_1083_n 0.00445602f $X=7.9 $Y=1.765 $X2=0
+ $Y2=0
cc_523 N_A_588_74#_c_612_n N_VPWR_c_1085_n 0.00445602f $X=8.35 $Y=1.765 $X2=0
+ $Y2=0
cc_524 N_A_588_74#_c_613_n N_VPWR_c_1085_n 0.00445602f $X=8.8 $Y=1.765 $X2=0
+ $Y2=0
cc_525 N_A_588_74#_c_618_n N_VPWR_c_1088_n 0.00445602f $X=11.05 $Y=1.765 $X2=0
+ $Y2=0
cc_526 N_A_588_74#_c_619_n N_VPWR_c_1088_n 0.00445602f $X=11.5 $Y=1.765 $X2=0
+ $Y2=0
cc_527 N_A_588_74#_c_620_n N_VPWR_c_1089_n 0.00413917f $X=11.95 $Y=1.765 $X2=0
+ $Y2=0
cc_528 N_A_588_74#_c_621_n N_VPWR_c_1089_n 0.00445602f $X=12.45 $Y=1.765 $X2=0
+ $Y2=0
cc_529 N_A_588_74#_c_606_n N_VPWR_c_1053_n 0.00857986f $X=5.6 $Y=1.765 $X2=0
+ $Y2=0
cc_530 N_A_588_74#_c_607_n N_VPWR_c_1053_n 0.00857378f $X=6.05 $Y=1.765 $X2=0
+ $Y2=0
cc_531 N_A_588_74#_c_608_n N_VPWR_c_1053_n 0.0085805f $X=6.55 $Y=1.765 $X2=0
+ $Y2=0
cc_532 N_A_588_74#_c_609_n N_VPWR_c_1053_n 0.00857589f $X=7 $Y=1.765 $X2=0 $Y2=0
cc_533 N_A_588_74#_c_610_n N_VPWR_c_1053_n 0.00857589f $X=7.45 $Y=1.765 $X2=0
+ $Y2=0
cc_534 N_A_588_74#_c_611_n N_VPWR_c_1053_n 0.00857589f $X=7.9 $Y=1.765 $X2=0
+ $Y2=0
cc_535 N_A_588_74#_c_612_n N_VPWR_c_1053_n 0.00857589f $X=8.35 $Y=1.765 $X2=0
+ $Y2=0
cc_536 N_A_588_74#_c_613_n N_VPWR_c_1053_n 0.00857589f $X=8.8 $Y=1.765 $X2=0
+ $Y2=0
cc_537 N_A_588_74#_c_614_n N_VPWR_c_1053_n 0.00857589f $X=9.25 $Y=1.765 $X2=0
+ $Y2=0
cc_538 N_A_588_74#_c_615_n N_VPWR_c_1053_n 0.00857589f $X=9.7 $Y=1.765 $X2=0
+ $Y2=0
cc_539 N_A_588_74#_c_616_n N_VPWR_c_1053_n 0.00857589f $X=10.15 $Y=1.765 $X2=0
+ $Y2=0
cc_540 N_A_588_74#_c_617_n N_VPWR_c_1053_n 0.00857589f $X=10.6 $Y=1.765 $X2=0
+ $Y2=0
cc_541 N_A_588_74#_c_618_n N_VPWR_c_1053_n 0.00857589f $X=11.05 $Y=1.765 $X2=0
+ $Y2=0
cc_542 N_A_588_74#_c_619_n N_VPWR_c_1053_n 0.00857589f $X=11.5 $Y=1.765 $X2=0
+ $Y2=0
cc_543 N_A_588_74#_c_620_n N_VPWR_c_1053_n 0.00818187f $X=11.95 $Y=1.765 $X2=0
+ $Y2=0
cc_544 N_A_588_74#_c_621_n N_VPWR_c_1053_n 0.00861561f $X=12.45 $Y=1.765 $X2=0
+ $Y2=0
cc_545 N_A_588_74#_c_623_n N_VPWR_c_1053_n 0.0119791f $X=3.105 $Y=2.815 $X2=0
+ $Y2=0
cc_546 N_A_588_74#_c_625_n N_VPWR_c_1053_n 0.0119791f $X=4.005 $Y=2.815 $X2=0
+ $Y2=0
cc_547 N_A_588_74#_c_628_n N_VPWR_c_1053_n 0.0119791f $X=4.915 $Y=2.815 $X2=0
+ $Y2=0
cc_548 N_A_588_74#_M1002_g N_X_c_1285_n 0.0142206f $X=5.585 $Y=0.74 $X2=0 $Y2=0
cc_549 N_A_588_74#_M1004_g N_X_c_1285_n 0.00312902f $X=6.015 $Y=0.74 $X2=0 $Y2=0
cc_550 N_A_588_74#_c_592_n N_X_c_1285_n 0.0255489f $X=4.915 $Y=1.99 $X2=0 $Y2=0
cc_551 N_A_588_74#_c_594_n N_X_c_1285_n 0.00478929f $X=4.975 $Y=1.32 $X2=0 $Y2=0
cc_552 N_A_588_74#_c_596_n N_X_c_1285_n 6.148e-19 $X=4.94 $Y=1.065 $X2=0 $Y2=0
cc_553 N_A_588_74#_c_597_n N_X_c_1285_n 0.0256633f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_554 N_A_588_74#_c_598_n N_X_c_1285_n 0.0301658f $X=6.21 $Y=1.485 $X2=0 $Y2=0
cc_555 N_A_588_74#_c_605_n N_X_c_1285_n 0.0251451f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_556 N_A_588_74#_c_606_n N_X_c_1296_n 0.00631728f $X=5.6 $Y=1.765 $X2=0 $Y2=0
cc_557 N_A_588_74#_c_607_n N_X_c_1296_n 0.00465475f $X=6.05 $Y=1.765 $X2=0 $Y2=0
cc_558 N_A_588_74#_c_592_n N_X_c_1296_n 0.00418771f $X=4.915 $Y=1.99 $X2=0 $Y2=0
cc_559 N_A_588_74#_c_597_n N_X_c_1296_n 0.00716941f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_560 N_A_588_74#_c_605_n N_X_c_1296_n 0.00215402f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_561 N_A_588_74#_c_606_n N_X_c_1297_n 0.00999652f $X=5.6 $Y=1.765 $X2=0 $Y2=0
cc_562 N_A_588_74#_c_607_n N_X_c_1297_n 0.00901091f $X=6.05 $Y=1.765 $X2=0 $Y2=0
cc_563 N_A_588_74#_M1007_g N_X_c_1286_n 0.00340636f $X=6.445 $Y=0.74 $X2=0 $Y2=0
cc_564 N_A_588_74#_M1011_g N_X_c_1286_n 0.00324826f $X=6.875 $Y=0.74 $X2=0 $Y2=0
cc_565 N_A_588_74#_c_598_n N_X_c_1286_n 0.0232726f $X=6.21 $Y=1.485 $X2=0 $Y2=0
cc_566 N_A_588_74#_c_599_n N_X_c_1286_n 0.0298139f $X=7.085 $Y=1.485 $X2=0 $Y2=0
cc_567 N_A_588_74#_c_605_n N_X_c_1286_n 0.0129665f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_568 N_A_588_74#_c_608_n N_X_c_1298_n 0.00969223f $X=6.55 $Y=1.765 $X2=0 $Y2=0
cc_569 N_A_588_74#_c_609_n N_X_c_1298_n 0.00961693f $X=7 $Y=1.765 $X2=0 $Y2=0
cc_570 N_A_588_74#_M1012_g N_X_c_1287_n 0.00345711f $X=7.305 $Y=0.74 $X2=0 $Y2=0
cc_571 N_A_588_74#_M1013_g N_X_c_1287_n 0.0143082f $X=7.735 $Y=0.74 $X2=0 $Y2=0
cc_572 N_A_588_74#_M1014_g N_X_c_1287_n 7.58559e-19 $X=8.235 $Y=0.74 $X2=0 $Y2=0
cc_573 N_A_588_74#_c_599_n N_X_c_1287_n 0.0233075f $X=7.085 $Y=1.485 $X2=0 $Y2=0
cc_574 N_A_588_74#_c_600_n N_X_c_1287_n 0.030056f $X=7.985 $Y=1.485 $X2=0 $Y2=0
cc_575 N_A_588_74#_c_605_n N_X_c_1287_n 0.0126181f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_576 N_A_588_74#_c_610_n N_X_c_1299_n 0.00961693f $X=7.45 $Y=1.765 $X2=0 $Y2=0
cc_577 N_A_588_74#_c_611_n N_X_c_1299_n 0.00961693f $X=7.9 $Y=1.765 $X2=0 $Y2=0
cc_578 N_A_588_74#_M1013_g N_X_c_1288_n 7.66254e-19 $X=7.735 $Y=0.74 $X2=0 $Y2=0
cc_579 N_A_588_74#_M1014_g N_X_c_1288_n 0.0146643f $X=8.235 $Y=0.74 $X2=0 $Y2=0
cc_580 N_A_588_74#_M1018_g N_X_c_1288_n 0.00346402f $X=8.665 $Y=0.74 $X2=0 $Y2=0
cc_581 N_A_588_74#_c_600_n N_X_c_1288_n 0.0233075f $X=7.985 $Y=1.485 $X2=0 $Y2=0
cc_582 N_A_588_74#_c_601_n N_X_c_1288_n 0.0302001f $X=8.905 $Y=1.485 $X2=0 $Y2=0
cc_583 N_A_588_74#_c_605_n N_X_c_1288_n 0.0126023f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_584 N_A_588_74#_c_612_n N_X_c_1300_n 0.00961693f $X=8.35 $Y=1.765 $X2=0 $Y2=0
cc_585 N_A_588_74#_c_613_n N_X_c_1300_n 0.00961693f $X=8.8 $Y=1.765 $X2=0 $Y2=0
cc_586 N_A_588_74#_M1018_g N_X_c_1289_n 7.72776e-19 $X=8.665 $Y=0.74 $X2=0 $Y2=0
cc_587 N_A_588_74#_M1021_g N_X_c_1289_n 0.0145949f $X=9.165 $Y=0.74 $X2=0 $Y2=0
cc_588 N_A_588_74#_M1022_g N_X_c_1289_n 0.00328496f $X=9.595 $Y=0.74 $X2=0 $Y2=0
cc_589 N_A_588_74#_c_601_n N_X_c_1289_n 0.0233081f $X=8.905 $Y=1.485 $X2=0 $Y2=0
cc_590 N_A_588_74#_c_602_n N_X_c_1289_n 0.0301915f $X=9.815 $Y=1.485 $X2=0 $Y2=0
cc_591 N_A_588_74#_c_605_n N_X_c_1289_n 0.0128404f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_592 N_A_588_74#_c_614_n N_X_c_1301_n 0.00961693f $X=9.25 $Y=1.765 $X2=0 $Y2=0
cc_593 N_A_588_74#_c_615_n N_X_c_1301_n 0.00961693f $X=9.7 $Y=1.765 $X2=0 $Y2=0
cc_594 N_A_588_74#_M1022_g N_X_c_1290_n 8.2524e-19 $X=9.595 $Y=0.74 $X2=0 $Y2=0
cc_595 N_A_588_74#_M1024_g N_X_c_1290_n 0.0145943f $X=10.095 $Y=0.74 $X2=0 $Y2=0
cc_596 N_A_588_74#_M1034_g N_X_c_1290_n 0.00541965f $X=10.525 $Y=0.74 $X2=0
+ $Y2=0
cc_597 N_A_588_74#_c_602_n N_X_c_1290_n 0.023362f $X=9.815 $Y=1.485 $X2=0 $Y2=0
cc_598 N_A_588_74#_c_603_n N_X_c_1290_n 0.0303238f $X=10.76 $Y=1.485 $X2=0 $Y2=0
cc_599 N_A_588_74#_c_605_n N_X_c_1290_n 0.0129045f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_600 N_A_588_74#_c_616_n N_X_c_1302_n 0.00961693f $X=10.15 $Y=1.765 $X2=0
+ $Y2=0
cc_601 N_A_588_74#_c_617_n N_X_c_1302_n 0.00961693f $X=10.6 $Y=1.765 $X2=0 $Y2=0
cc_602 N_A_588_74#_c_617_n N_X_c_1291_n 0.0011387f $X=10.6 $Y=1.765 $X2=0 $Y2=0
cc_603 N_A_588_74#_M1037_g N_X_c_1291_n 0.00562543f $X=11.025 $Y=0.74 $X2=0
+ $Y2=0
cc_604 N_A_588_74#_c_618_n N_X_c_1291_n 0.00331751f $X=11.05 $Y=1.765 $X2=0
+ $Y2=0
cc_605 N_A_588_74#_M1040_g N_X_c_1291_n 0.00527627f $X=11.455 $Y=0.74 $X2=0
+ $Y2=0
cc_606 N_A_588_74#_c_619_n N_X_c_1291_n 0.00327622f $X=11.5 $Y=1.765 $X2=0 $Y2=0
cc_607 N_A_588_74#_c_597_n N_X_c_1291_n 0.0256842f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_608 N_A_588_74#_c_603_n N_X_c_1291_n 0.0302662f $X=10.76 $Y=1.485 $X2=0 $Y2=0
cc_609 N_A_588_74#_c_604_n N_X_c_1291_n 0.0302916f $X=11.685 $Y=1.485 $X2=0
+ $Y2=0
cc_610 N_A_588_74#_c_605_n N_X_c_1291_n 0.025039f $X=12.395 $Y=1.542 $X2=0 $Y2=0
cc_611 N_A_588_74#_c_618_n N_X_c_1304_n 0.00961693f $X=11.05 $Y=1.765 $X2=0
+ $Y2=0
cc_612 N_A_588_74#_c_619_n N_X_c_1304_n 0.00961693f $X=11.5 $Y=1.765 $X2=0 $Y2=0
cc_613 N_A_588_74#_M1040_g N_X_c_1292_n 2.35461e-19 $X=11.455 $Y=0.74 $X2=0
+ $Y2=0
cc_614 N_A_588_74#_M1042_g N_X_c_1292_n 0.0078247f $X=11.965 $Y=0.74 $X2=0 $Y2=0
cc_615 N_A_588_74#_M1045_g N_X_c_1292_n 0.00794138f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_616 N_A_588_74#_c_620_n N_X_c_1293_n 0.00836331f $X=11.95 $Y=1.765 $X2=0
+ $Y2=0
cc_617 N_A_588_74#_M1042_g N_X_c_1293_n 0.00465421f $X=11.965 $Y=0.74 $X2=0
+ $Y2=0
cc_618 N_A_588_74#_M1045_g N_X_c_1293_n 0.00881083f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_619 N_A_588_74#_c_621_n N_X_c_1293_n 0.00192244f $X=12.45 $Y=1.765 $X2=0
+ $Y2=0
cc_620 N_A_588_74#_c_597_n N_X_c_1293_n 0.00283069f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_621 N_A_588_74#_c_604_n N_X_c_1293_n 0.0314793f $X=11.685 $Y=1.485 $X2=0
+ $Y2=0
cc_622 N_A_588_74#_c_605_n N_X_c_1293_n 0.0411045f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_623 N_A_588_74#_c_621_n N_X_c_1306_n 0.00943968f $X=12.45 $Y=1.765 $X2=0
+ $Y2=0
cc_624 N_A_588_74#_c_597_n N_X_c_1391_n 0.0192444f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_625 N_A_588_74#_c_605_n N_X_c_1391_n 0.0101332f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_626 N_A_588_74#_c_597_n N_X_c_1393_n 0.023376f $X=11.685 $Y=1.665 $X2=0 $Y2=0
cc_627 N_A_588_74#_c_605_n N_X_c_1393_n 0.0133147f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_628 N_A_588_74#_c_597_n N_X_c_1395_n 0.023376f $X=11.685 $Y=1.665 $X2=0 $Y2=0
cc_629 N_A_588_74#_c_605_n N_X_c_1395_n 0.0132989f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_630 N_A_588_74#_c_597_n N_X_c_1397_n 0.0208971f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_631 N_A_588_74#_c_605_n N_X_c_1397_n 0.0113574f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_632 N_A_588_74#_c_597_n N_X_c_1399_n 0.0194235f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_633 N_A_588_74#_c_605_n N_X_c_1399_n 0.0104676f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_634 N_A_588_74#_M1042_g N_X_c_1294_n 0.00358838f $X=11.965 $Y=0.74 $X2=0
+ $Y2=0
cc_635 N_A_588_74#_M1045_g N_X_c_1294_n 0.00288102f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_636 N_A_588_74#_c_608_n N_X_c_1403_n 0.001146f $X=6.55 $Y=1.765 $X2=0 $Y2=0
cc_637 N_A_588_74#_c_609_n N_X_c_1403_n 0.00145229f $X=7 $Y=1.765 $X2=0 $Y2=0
cc_638 N_A_588_74#_c_610_n N_X_c_1403_n 4.2577e-19 $X=7.45 $Y=1.765 $X2=0 $Y2=0
cc_639 N_A_588_74#_c_597_n N_X_c_1403_n 0.00136816f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_640 N_A_588_74#_c_605_n N_X_c_1403_n 0.00366161f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_641 N_A_588_74#_c_607_n N_X_c_1307_n 0.00113009f $X=6.05 $Y=1.765 $X2=0 $Y2=0
cc_642 N_A_588_74#_c_608_n N_X_c_1307_n 0.00327936f $X=6.55 $Y=1.765 $X2=0 $Y2=0
cc_643 N_A_588_74#_c_609_n N_X_c_1307_n 0.00295629f $X=7 $Y=1.765 $X2=0 $Y2=0
cc_644 N_A_588_74#_c_597_n N_X_c_1307_n 0.00869127f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_645 N_A_588_74#_c_598_n N_X_c_1307_n 0.00464651f $X=6.21 $Y=1.485 $X2=0 $Y2=0
cc_646 N_A_588_74#_c_605_n N_X_c_1307_n 0.00339568f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_647 N_A_588_74#_c_610_n N_X_c_1414_n 0.00114251f $X=7.45 $Y=1.765 $X2=0 $Y2=0
cc_648 N_A_588_74#_c_611_n N_X_c_1414_n 0.00145229f $X=7.9 $Y=1.765 $X2=0 $Y2=0
cc_649 N_A_588_74#_c_597_n N_X_c_1414_n 0.00136816f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_650 N_A_588_74#_c_605_n N_X_c_1414_n 0.00366161f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_651 N_A_588_74#_c_609_n N_X_c_1308_n 0.00120072f $X=7 $Y=1.765 $X2=0 $Y2=0
cc_652 N_A_588_74#_c_610_n N_X_c_1308_n 0.00318335f $X=7.45 $Y=1.765 $X2=0 $Y2=0
cc_653 N_A_588_74#_c_611_n N_X_c_1308_n 0.00295629f $X=7.9 $Y=1.765 $X2=0 $Y2=0
cc_654 N_A_588_74#_c_597_n N_X_c_1308_n 0.00888655f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_655 N_A_588_74#_c_599_n N_X_c_1308_n 0.00378597f $X=7.085 $Y=1.485 $X2=0
+ $Y2=0
cc_656 N_A_588_74#_c_605_n N_X_c_1308_n 0.00351046f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_657 N_A_588_74#_c_612_n N_X_c_1424_n 0.00114251f $X=8.35 $Y=1.765 $X2=0 $Y2=0
cc_658 N_A_588_74#_c_613_n N_X_c_1424_n 0.00145229f $X=8.8 $Y=1.765 $X2=0 $Y2=0
cc_659 N_A_588_74#_c_597_n N_X_c_1424_n 0.00136816f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_660 N_A_588_74#_c_605_n N_X_c_1424_n 0.00366161f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_661 N_A_588_74#_c_611_n N_X_c_1309_n 0.00113893f $X=7.9 $Y=1.765 $X2=0 $Y2=0
cc_662 N_A_588_74#_c_612_n N_X_c_1309_n 0.00318335f $X=8.35 $Y=1.765 $X2=0 $Y2=0
cc_663 N_A_588_74#_c_613_n N_X_c_1309_n 0.00295629f $X=8.8 $Y=1.765 $X2=0 $Y2=0
cc_664 N_A_588_74#_c_597_n N_X_c_1309_n 0.00888655f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_665 N_A_588_74#_c_600_n N_X_c_1309_n 0.00378597f $X=7.985 $Y=1.485 $X2=0
+ $Y2=0
cc_666 N_A_588_74#_c_605_n N_X_c_1309_n 0.00351046f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_667 N_A_588_74#_c_614_n N_X_c_1434_n 0.00114251f $X=9.25 $Y=1.765 $X2=0 $Y2=0
cc_668 N_A_588_74#_c_615_n N_X_c_1434_n 0.00145229f $X=9.7 $Y=1.765 $X2=0 $Y2=0
cc_669 N_A_588_74#_c_597_n N_X_c_1434_n 0.00136816f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_670 N_A_588_74#_c_605_n N_X_c_1434_n 0.00366161f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_671 N_A_588_74#_c_613_n N_X_c_1310_n 0.00113893f $X=8.8 $Y=1.765 $X2=0 $Y2=0
cc_672 N_A_588_74#_c_614_n N_X_c_1310_n 0.00318335f $X=9.25 $Y=1.765 $X2=0 $Y2=0
cc_673 N_A_588_74#_c_615_n N_X_c_1310_n 0.00295629f $X=9.7 $Y=1.765 $X2=0 $Y2=0
cc_674 N_A_588_74#_c_597_n N_X_c_1310_n 0.00877275f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_675 N_A_588_74#_c_601_n N_X_c_1310_n 0.00426873f $X=8.905 $Y=1.485 $X2=0
+ $Y2=0
cc_676 N_A_588_74#_c_605_n N_X_c_1310_n 0.00345221f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_677 N_A_588_74#_c_616_n N_X_c_1444_n 0.00114251f $X=10.15 $Y=1.765 $X2=0
+ $Y2=0
cc_678 N_A_588_74#_c_617_n N_X_c_1444_n 0.00145229f $X=10.6 $Y=1.765 $X2=0 $Y2=0
cc_679 N_A_588_74#_c_597_n N_X_c_1444_n 0.00125217f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_680 N_A_588_74#_c_605_n N_X_c_1444_n 0.00325044f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_681 N_A_588_74#_c_615_n N_X_c_1311_n 0.00113884f $X=9.7 $Y=1.765 $X2=0 $Y2=0
cc_682 N_A_588_74#_c_616_n N_X_c_1311_n 0.00323056f $X=10.15 $Y=1.765 $X2=0
+ $Y2=0
cc_683 N_A_588_74#_c_617_n N_X_c_1311_n 0.00306306f $X=10.6 $Y=1.765 $X2=0 $Y2=0
cc_684 N_A_588_74#_c_597_n N_X_c_1311_n 0.00907039f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_685 N_A_588_74#_c_602_n N_X_c_1311_n 0.00486082f $X=9.815 $Y=1.485 $X2=0
+ $Y2=0
cc_686 N_A_588_74#_c_605_n N_X_c_1311_n 0.00347167f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_687 N_A_588_74#_c_618_n N_X_c_1454_n 0.00114251f $X=11.05 $Y=1.765 $X2=0
+ $Y2=0
cc_688 N_A_588_74#_c_619_n N_X_c_1454_n 0.00145586f $X=11.5 $Y=1.765 $X2=0 $Y2=0
cc_689 N_A_588_74#_c_620_n N_X_c_1454_n 4.18597e-19 $X=11.95 $Y=1.765 $X2=0
+ $Y2=0
cc_690 N_A_588_74#_c_597_n N_X_c_1454_n 0.00102018f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_691 N_A_588_74#_c_605_n N_X_c_1454_n 0.00242812f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_692 N_A_588_74#_c_621_n N_X_c_1459_n 0.00230104f $X=12.45 $Y=1.765 $X2=0
+ $Y2=0
cc_693 N_A_588_74#_c_605_n N_X_c_1459_n 8.23484e-19 $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_694 N_A_588_74#_c_607_n N_X_c_1461_n 0.00863624f $X=6.05 $Y=1.765 $X2=0 $Y2=0
cc_695 N_A_588_74#_c_608_n N_X_c_1461_n 0.0083567f $X=6.55 $Y=1.765 $X2=0 $Y2=0
cc_696 N_A_588_74#_c_609_n N_X_c_1461_n 0.00808368f $X=7 $Y=1.765 $X2=0 $Y2=0
cc_697 N_A_588_74#_c_610_n N_X_c_1461_n 0.00801383f $X=7.45 $Y=1.765 $X2=0 $Y2=0
cc_698 N_A_588_74#_c_611_n N_X_c_1461_n 0.00671038f $X=7.9 $Y=1.765 $X2=0 $Y2=0
cc_699 N_A_588_74#_c_612_n N_X_c_1461_n 0.00663712f $X=8.35 $Y=1.765 $X2=0 $Y2=0
cc_700 N_A_588_74#_c_613_n N_X_c_1461_n 0.00671038f $X=8.8 $Y=1.765 $X2=0 $Y2=0
cc_701 N_A_588_74#_c_614_n N_X_c_1461_n 0.00672667f $X=9.25 $Y=1.765 $X2=0 $Y2=0
cc_702 N_A_588_74#_c_615_n N_X_c_1461_n 0.00671038f $X=9.7 $Y=1.765 $X2=0 $Y2=0
cc_703 N_A_588_74#_c_616_n N_X_c_1461_n 0.00681622f $X=10.15 $Y=1.765 $X2=0
+ $Y2=0
cc_704 N_A_588_74#_c_617_n N_X_c_1461_n 0.0067616f $X=10.6 $Y=1.765 $X2=0 $Y2=0
cc_705 N_A_588_74#_c_618_n N_X_c_1461_n 0.00701605f $X=11.05 $Y=1.765 $X2=0
+ $Y2=0
cc_706 N_A_588_74#_c_619_n N_X_c_1461_n 0.00686404f $X=11.5 $Y=1.765 $X2=0 $Y2=0
cc_707 N_A_588_74#_c_620_n N_X_c_1461_n 0.0135342f $X=11.95 $Y=1.765 $X2=0 $Y2=0
cc_708 N_A_588_74#_c_621_n N_X_c_1461_n 9.10578e-19 $X=12.45 $Y=1.765 $X2=0
+ $Y2=0
cc_709 N_A_588_74#_c_597_n N_X_c_1461_n 0.609641f $X=11.685 $Y=1.665 $X2=0 $Y2=0
cc_710 N_A_588_74#_c_598_n N_X_c_1461_n 0.0021687f $X=6.21 $Y=1.485 $X2=0 $Y2=0
cc_711 N_A_588_74#_c_599_n N_X_c_1461_n 0.00287155f $X=7.085 $Y=1.485 $X2=0
+ $Y2=0
cc_712 N_A_588_74#_c_600_n N_X_c_1461_n 0.00286681f $X=7.985 $Y=1.485 $X2=0
+ $Y2=0
cc_713 N_A_588_74#_c_601_n N_X_c_1461_n 0.00296141f $X=8.905 $Y=1.485 $X2=0
+ $Y2=0
cc_714 N_A_588_74#_c_602_n N_X_c_1461_n 0.00305601f $X=9.815 $Y=1.485 $X2=0
+ $Y2=0
cc_715 N_A_588_74#_c_603_n N_X_c_1461_n 0.00313509f $X=10.76 $Y=1.485 $X2=0
+ $Y2=0
cc_716 N_A_588_74#_c_604_n N_X_c_1461_n 0.00404503f $X=11.685 $Y=1.485 $X2=0
+ $Y2=0
cc_717 N_A_588_74#_c_605_n N_X_c_1461_n 0.00627731f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_718 N_A_588_74#_c_588_n N_VGND_M1006_s 0.00250873f $X=3.845 $Y=1.065 $X2=0
+ $Y2=0
cc_719 N_A_588_74#_c_591_n N_VGND_M1027_s 0.00250873f $X=4.775 $Y=1.065 $X2=0
+ $Y2=0
cc_720 N_A_588_74#_c_587_n N_VGND_c_1570_n 0.023409f $X=3.08 $Y=0.515 $X2=0
+ $Y2=0
cc_721 N_A_588_74#_c_589_n N_VGND_c_1570_n 0.00711243f $X=3.165 $Y=1.065 $X2=0
+ $Y2=0
cc_722 N_A_588_74#_c_587_n N_VGND_c_1571_n 0.017215f $X=3.08 $Y=0.515 $X2=0
+ $Y2=0
cc_723 N_A_588_74#_c_588_n N_VGND_c_1571_n 0.0209867f $X=3.845 $Y=1.065 $X2=0
+ $Y2=0
cc_724 N_A_588_74#_c_590_n N_VGND_c_1571_n 0.0173318f $X=4.01 $Y=0.515 $X2=0
+ $Y2=0
cc_725 N_A_588_74#_c_590_n N_VGND_c_1572_n 0.017215f $X=4.01 $Y=0.515 $X2=0
+ $Y2=0
cc_726 N_A_588_74#_c_591_n N_VGND_c_1572_n 0.0209867f $X=4.775 $Y=1.065 $X2=0
+ $Y2=0
cc_727 N_A_588_74#_c_593_n N_VGND_c_1572_n 0.0173318f $X=4.94 $Y=0.515 $X2=0
+ $Y2=0
cc_728 N_A_588_74#_M1002_g N_VGND_c_1573_n 0.00171481f $X=5.585 $Y=0.74 $X2=0
+ $Y2=0
cc_729 N_A_588_74#_c_592_n N_VGND_c_1573_n 0.0101469f $X=4.915 $Y=1.99 $X2=0
+ $Y2=0
cc_730 N_A_588_74#_c_593_n N_VGND_c_1573_n 0.00112941f $X=4.94 $Y=0.515 $X2=0
+ $Y2=0
cc_731 N_A_588_74#_c_596_n N_VGND_c_1573_n 0.00704273f $X=4.94 $Y=1.065 $X2=0
+ $Y2=0
cc_732 N_A_588_74#_c_597_n N_VGND_c_1573_n 0.00278617f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_733 N_A_588_74#_M1002_g N_VGND_c_1574_n 6.16849e-19 $X=5.585 $Y=0.74 $X2=0
+ $Y2=0
cc_734 N_A_588_74#_M1004_g N_VGND_c_1574_n 0.0128539f $X=6.015 $Y=0.74 $X2=0
+ $Y2=0
cc_735 N_A_588_74#_M1007_g N_VGND_c_1574_n 0.00204911f $X=6.445 $Y=0.74 $X2=0
+ $Y2=0
cc_736 N_A_588_74#_c_597_n N_VGND_c_1574_n 0.00128328f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_737 N_A_588_74#_c_598_n N_VGND_c_1574_n 0.0183169f $X=6.21 $Y=1.485 $X2=0
+ $Y2=0
cc_738 N_A_588_74#_c_605_n N_VGND_c_1574_n 7.80261e-19 $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_739 N_A_588_74#_M1007_g N_VGND_c_1575_n 0.00461464f $X=6.445 $Y=0.74 $X2=0
+ $Y2=0
cc_740 N_A_588_74#_M1011_g N_VGND_c_1575_n 0.00461464f $X=6.875 $Y=0.74 $X2=0
+ $Y2=0
cc_741 N_A_588_74#_M1011_g N_VGND_c_1576_n 0.00217717f $X=6.875 $Y=0.74 $X2=0
+ $Y2=0
cc_742 N_A_588_74#_M1012_g N_VGND_c_1576_n 0.00203758f $X=7.305 $Y=0.74 $X2=0
+ $Y2=0
cc_743 N_A_588_74#_c_597_n N_VGND_c_1576_n 0.00111156f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_744 N_A_588_74#_c_599_n N_VGND_c_1576_n 0.0158153f $X=7.085 $Y=1.485 $X2=0
+ $Y2=0
cc_745 N_A_588_74#_c_605_n N_VGND_c_1576_n 7.76654e-19 $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_746 N_A_588_74#_M1012_g N_VGND_c_1577_n 0.00461464f $X=7.305 $Y=0.74 $X2=0
+ $Y2=0
cc_747 N_A_588_74#_M1013_g N_VGND_c_1577_n 0.00439937f $X=7.735 $Y=0.74 $X2=0
+ $Y2=0
cc_748 N_A_588_74#_M1013_g N_VGND_c_1578_n 0.00232598f $X=7.735 $Y=0.74 $X2=0
+ $Y2=0
cc_749 N_A_588_74#_M1014_g N_VGND_c_1578_n 0.00579981f $X=8.235 $Y=0.74 $X2=0
+ $Y2=0
cc_750 N_A_588_74#_c_597_n N_VGND_c_1578_n 0.00137249f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_751 N_A_588_74#_c_600_n N_VGND_c_1578_n 0.019527f $X=7.985 $Y=1.485 $X2=0
+ $Y2=0
cc_752 N_A_588_74#_c_605_n N_VGND_c_1578_n 0.0013193f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_753 N_A_588_74#_M1018_g N_VGND_c_1579_n 0.00245186f $X=8.665 $Y=0.74 $X2=0
+ $Y2=0
cc_754 N_A_588_74#_M1021_g N_VGND_c_1579_n 0.00580958f $X=9.165 $Y=0.74 $X2=0
+ $Y2=0
cc_755 N_A_588_74#_c_597_n N_VGND_c_1579_n 0.00152905f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_756 N_A_588_74#_c_601_n N_VGND_c_1579_n 0.0217547f $X=8.905 $Y=1.485 $X2=0
+ $Y2=0
cc_757 N_A_588_74#_c_605_n N_VGND_c_1579_n 0.00132195f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_758 N_A_588_74#_M1021_g N_VGND_c_1580_n 5.94534e-19 $X=9.165 $Y=0.74 $X2=0
+ $Y2=0
cc_759 N_A_588_74#_M1022_g N_VGND_c_1580_n 0.0114917f $X=9.595 $Y=0.74 $X2=0
+ $Y2=0
cc_760 N_A_588_74#_M1024_g N_VGND_c_1580_n 0.00579705f $X=10.095 $Y=0.74 $X2=0
+ $Y2=0
cc_761 N_A_588_74#_c_597_n N_VGND_c_1580_n 0.00160551f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_762 N_A_588_74#_c_602_n N_VGND_c_1580_n 0.0228524f $X=9.815 $Y=1.485 $X2=0
+ $Y2=0
cc_763 N_A_588_74#_c_605_n N_VGND_c_1580_n 0.00132461f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_764 N_A_588_74#_M1024_g N_VGND_c_1581_n 6.13445e-19 $X=10.095 $Y=0.74 $X2=0
+ $Y2=0
cc_765 N_A_588_74#_M1034_g N_VGND_c_1581_n 0.0134511f $X=10.525 $Y=0.74 $X2=0
+ $Y2=0
cc_766 N_A_588_74#_M1037_g N_VGND_c_1581_n 0.00583686f $X=11.025 $Y=0.74 $X2=0
+ $Y2=0
cc_767 N_A_588_74#_c_597_n N_VGND_c_1581_n 0.00170077f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_768 N_A_588_74#_c_603_n N_VGND_c_1581_n 0.0242563f $X=10.76 $Y=1.485 $X2=0
+ $Y2=0
cc_769 N_A_588_74#_c_605_n N_VGND_c_1581_n 0.00132644f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_770 N_A_588_74#_M1037_g N_VGND_c_1582_n 5.68036e-19 $X=11.025 $Y=0.74 $X2=0
+ $Y2=0
cc_771 N_A_588_74#_M1040_g N_VGND_c_1582_n 0.0134929f $X=11.455 $Y=0.74 $X2=0
+ $Y2=0
cc_772 N_A_588_74#_M1042_g N_VGND_c_1582_n 0.00727688f $X=11.965 $Y=0.74 $X2=0
+ $Y2=0
cc_773 N_A_588_74#_c_597_n N_VGND_c_1582_n 0.00167989f $X=11.685 $Y=1.665 $X2=0
+ $Y2=0
cc_774 N_A_588_74#_c_604_n N_VGND_c_1582_n 0.0242765f $X=11.685 $Y=1.485 $X2=0
+ $Y2=0
cc_775 N_A_588_74#_c_605_n N_VGND_c_1582_n 0.00140447f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_776 N_A_588_74#_M1045_g N_VGND_c_1584_n 0.0198727f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_777 N_A_588_74#_c_605_n N_VGND_c_1584_n 0.00109954f $X=12.395 $Y=1.542 $X2=0
+ $Y2=0
cc_778 N_A_588_74#_c_587_n N_VGND_c_1587_n 0.0109942f $X=3.08 $Y=0.515 $X2=0
+ $Y2=0
cc_779 N_A_588_74#_c_590_n N_VGND_c_1589_n 0.0109942f $X=4.01 $Y=0.515 $X2=0
+ $Y2=0
cc_780 N_A_588_74#_c_593_n N_VGND_c_1591_n 0.0109942f $X=4.94 $Y=0.515 $X2=0
+ $Y2=0
cc_781 N_A_588_74#_M1002_g N_VGND_c_1593_n 0.00434272f $X=5.585 $Y=0.74 $X2=0
+ $Y2=0
cc_782 N_A_588_74#_M1004_g N_VGND_c_1593_n 0.00383152f $X=6.015 $Y=0.74 $X2=0
+ $Y2=0
cc_783 N_A_588_74#_M1037_g N_VGND_c_1595_n 0.00461464f $X=11.025 $Y=0.74 $X2=0
+ $Y2=0
cc_784 N_A_588_74#_M1040_g N_VGND_c_1595_n 0.00383152f $X=11.455 $Y=0.74 $X2=0
+ $Y2=0
cc_785 N_A_588_74#_M1014_g N_VGND_c_1599_n 0.00434272f $X=8.235 $Y=0.74 $X2=0
+ $Y2=0
cc_786 N_A_588_74#_M1018_g N_VGND_c_1599_n 0.00461464f $X=8.665 $Y=0.74 $X2=0
+ $Y2=0
cc_787 N_A_588_74#_M1021_g N_VGND_c_1600_n 0.00434272f $X=9.165 $Y=0.74 $X2=0
+ $Y2=0
cc_788 N_A_588_74#_M1022_g N_VGND_c_1600_n 0.00444681f $X=9.595 $Y=0.74 $X2=0
+ $Y2=0
cc_789 N_A_588_74#_M1024_g N_VGND_c_1601_n 0.00434272f $X=10.095 $Y=0.74 $X2=0
+ $Y2=0
cc_790 N_A_588_74#_M1034_g N_VGND_c_1601_n 0.00383152f $X=10.525 $Y=0.74 $X2=0
+ $Y2=0
cc_791 N_A_588_74#_M1042_g N_VGND_c_1602_n 0.00434272f $X=11.965 $Y=0.74 $X2=0
+ $Y2=0
cc_792 N_A_588_74#_M1045_g N_VGND_c_1602_n 0.00434272f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_793 N_A_588_74#_M1002_g N_VGND_c_1610_n 0.00820382f $X=5.585 $Y=0.74 $X2=0
+ $Y2=0
cc_794 N_A_588_74#_M1004_g N_VGND_c_1610_n 0.0075754f $X=6.015 $Y=0.74 $X2=0
+ $Y2=0
cc_795 N_A_588_74#_M1007_g N_VGND_c_1610_n 0.00908333f $X=6.445 $Y=0.74 $X2=0
+ $Y2=0
cc_796 N_A_588_74#_M1011_g N_VGND_c_1610_n 0.00907324f $X=6.875 $Y=0.74 $X2=0
+ $Y2=0
cc_797 N_A_588_74#_M1012_g N_VGND_c_1610_n 0.00908333f $X=7.305 $Y=0.74 $X2=0
+ $Y2=0
cc_798 N_A_588_74#_M1013_g N_VGND_c_1610_n 0.0083895f $X=7.735 $Y=0.74 $X2=0
+ $Y2=0
cc_799 N_A_588_74#_M1014_g N_VGND_c_1610_n 0.00820718f $X=8.235 $Y=0.74 $X2=0
+ $Y2=0
cc_800 N_A_588_74#_M1018_g N_VGND_c_1610_n 0.00907983f $X=8.665 $Y=0.74 $X2=0
+ $Y2=0
cc_801 N_A_588_74#_M1021_g N_VGND_c_1610_n 0.00820718f $X=9.165 $Y=0.74 $X2=0
+ $Y2=0
cc_802 N_A_588_74#_M1022_g N_VGND_c_1610_n 0.00877518f $X=9.595 $Y=0.74 $X2=0
+ $Y2=0
cc_803 N_A_588_74#_M1024_g N_VGND_c_1610_n 0.00820718f $X=10.095 $Y=0.74 $X2=0
+ $Y2=0
cc_804 N_A_588_74#_M1034_g N_VGND_c_1610_n 0.0075754f $X=10.525 $Y=0.74 $X2=0
+ $Y2=0
cc_805 N_A_588_74#_M1037_g N_VGND_c_1610_n 0.00908767f $X=11.025 $Y=0.74 $X2=0
+ $Y2=0
cc_806 N_A_588_74#_M1040_g N_VGND_c_1610_n 0.0075754f $X=11.455 $Y=0.74 $X2=0
+ $Y2=0
cc_807 N_A_588_74#_M1042_g N_VGND_c_1610_n 0.00821029f $X=11.965 $Y=0.74 $X2=0
+ $Y2=0
cc_808 N_A_588_74#_M1045_g N_VGND_c_1610_n 0.00823934f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_809 N_A_588_74#_c_587_n N_VGND_c_1610_n 0.00904371f $X=3.08 $Y=0.515 $X2=0
+ $Y2=0
cc_810 N_A_588_74#_c_590_n N_VGND_c_1610_n 0.00904371f $X=4.01 $Y=0.515 $X2=0
+ $Y2=0
cc_811 N_A_588_74#_c_593_n N_VGND_c_1610_n 0.00904371f $X=4.94 $Y=0.515 $X2=0
+ $Y2=0
cc_812 N_VPWR_c_1059_n N_X_c_1296_n 0.00897508f $X=5.365 $Y=2.09 $X2=0 $Y2=0
cc_813 N_VPWR_c_1060_n N_X_c_1296_n 0.00812812f $X=6.325 $Y=2.325 $X2=0 $Y2=0
cc_814 N_VPWR_c_1059_n N_X_c_1297_n 0.0556989f $X=5.365 $Y=2.09 $X2=0 $Y2=0
cc_815 N_VPWR_c_1060_n N_X_c_1297_n 0.0351499f $X=6.325 $Y=2.325 $X2=0 $Y2=0
cc_816 N_VPWR_c_1079_n N_X_c_1297_n 0.014552f $X=6.16 $Y=3.33 $X2=0 $Y2=0
cc_817 N_VPWR_c_1053_n N_X_c_1297_n 0.0119791f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_818 N_VPWR_c_1081_n N_X_c_1298_n 0.014552f $X=7.14 $Y=3.33 $X2=0 $Y2=0
cc_819 N_VPWR_c_1053_n N_X_c_1298_n 0.0119791f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_820 N_VPWR_c_1083_n N_X_c_1299_n 0.014552f $X=8.04 $Y=3.33 $X2=0 $Y2=0
cc_821 N_VPWR_c_1053_n N_X_c_1299_n 0.0119791f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_822 N_VPWR_c_1085_n N_X_c_1300_n 0.014552f $X=8.94 $Y=3.33 $X2=0 $Y2=0
cc_823 N_VPWR_c_1053_n N_X_c_1300_n 0.0119791f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_824 N_VPWR_c_1064_n N_X_c_1301_n 0.014552f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_825 N_VPWR_c_1053_n N_X_c_1301_n 0.0119791f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_826 N_VPWR_c_1066_n N_X_c_1302_n 0.014552f $X=10.74 $Y=3.33 $X2=0 $Y2=0
cc_827 N_VPWR_c_1053_n N_X_c_1302_n 0.0119791f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_828 N_VPWR_c_1088_n N_X_c_1304_n 0.014552f $X=11.64 $Y=3.33 $X2=0 $Y2=0
cc_829 N_VPWR_c_1053_n N_X_c_1304_n 0.0119791f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_830 N_VPWR_c_1068_n N_X_c_1293_n 0.0419868f $X=11.725 $Y=2.09 $X2=0 $Y2=0
cc_831 N_VPWR_c_1070_n N_X_c_1293_n 0.00687696f $X=12.675 $Y=1.985 $X2=0 $Y2=0
cc_832 N_VPWR_c_1089_n N_X_c_1306_n 0.0145938f $X=12.59 $Y=3.33 $X2=0 $Y2=0
cc_833 N_VPWR_c_1053_n N_X_c_1306_n 0.0120466f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_834 N_VPWR_c_1060_n N_X_c_1403_n 0.0683802f $X=6.325 $Y=2.325 $X2=0 $Y2=0
cc_835 N_VPWR_c_1061_n N_X_c_1403_n 0.0667435f $X=7.225 $Y=2.325 $X2=0 $Y2=0
cc_836 N_VPWR_c_1061_n N_X_c_1414_n 0.0667435f $X=7.225 $Y=2.325 $X2=0 $Y2=0
cc_837 N_VPWR_c_1062_n N_X_c_1414_n 0.0667435f $X=8.125 $Y=2.09 $X2=0 $Y2=0
cc_838 N_VPWR_c_1062_n N_X_c_1424_n 0.0667435f $X=8.125 $Y=2.09 $X2=0 $Y2=0
cc_839 N_VPWR_c_1063_n N_X_c_1424_n 0.0667435f $X=9.025 $Y=2.09 $X2=0 $Y2=0
cc_840 N_VPWR_c_1063_n N_X_c_1434_n 0.0667435f $X=9.025 $Y=2.09 $X2=0 $Y2=0
cc_841 N_VPWR_c_1065_n N_X_c_1434_n 0.0667435f $X=9.925 $Y=2.09 $X2=0 $Y2=0
cc_842 N_VPWR_c_1065_n N_X_c_1444_n 0.0667435f $X=9.925 $Y=2.09 $X2=0 $Y2=0
cc_843 N_VPWR_c_1067_n N_X_c_1444_n 0.0667435f $X=10.825 $Y=2.09 $X2=0 $Y2=0
cc_844 N_VPWR_c_1067_n N_X_c_1454_n 0.0667435f $X=10.825 $Y=2.09 $X2=0 $Y2=0
cc_845 N_VPWR_c_1068_n N_X_c_1454_n 0.0683802f $X=11.725 $Y=2.09 $X2=0 $Y2=0
cc_846 N_VPWR_c_1070_n N_X_c_1459_n 0.0633666f $X=12.675 $Y=1.985 $X2=0 $Y2=0
cc_847 N_VPWR_M1008_s N_X_c_1461_n 0.00574927f $X=6.125 $Y=1.84 $X2=0 $Y2=0
cc_848 N_VPWR_M1010_s N_X_c_1461_n 0.00688909f $X=7.075 $Y=1.84 $X2=0 $Y2=0
cc_849 N_VPWR_M1017_s N_X_c_1461_n 0.00687795f $X=7.975 $Y=1.84 $X2=0 $Y2=0
cc_850 N_VPWR_M1020_s N_X_c_1461_n 0.00680435f $X=8.875 $Y=1.84 $X2=0 $Y2=0
cc_851 N_VPWR_M1033_s N_X_c_1461_n 0.00673074f $X=9.775 $Y=1.84 $X2=0 $Y2=0
cc_852 N_VPWR_M1038_s N_X_c_1461_n 0.00657127f $X=10.675 $Y=1.84 $X2=0 $Y2=0
cc_853 N_VPWR_M1044_s N_X_c_1461_n 0.00406632f $X=11.575 $Y=1.84 $X2=0 $Y2=0
cc_854 N_VPWR_c_1059_n N_X_c_1461_n 0.00144666f $X=5.365 $Y=2.09 $X2=0 $Y2=0
cc_855 N_VPWR_c_1060_n N_X_c_1461_n 0.0256929f $X=6.325 $Y=2.325 $X2=0 $Y2=0
cc_856 N_VPWR_c_1061_n N_X_c_1461_n 0.0198929f $X=7.225 $Y=2.325 $X2=0 $Y2=0
cc_857 N_VPWR_c_1062_n N_X_c_1461_n 0.0198929f $X=8.125 $Y=2.09 $X2=0 $Y2=0
cc_858 N_VPWR_c_1063_n N_X_c_1461_n 0.0195347f $X=9.025 $Y=2.09 $X2=0 $Y2=0
cc_859 N_VPWR_c_1065_n N_X_c_1461_n 0.0191765f $X=9.925 $Y=2.09 $X2=0 $Y2=0
cc_860 N_VPWR_c_1067_n N_X_c_1461_n 0.0187586f $X=10.825 $Y=2.09 $X2=0 $Y2=0
cc_861 N_VPWR_c_1068_n N_X_c_1461_n 0.0249485f $X=11.725 $Y=2.09 $X2=0 $Y2=0
cc_862 N_VPWR_c_1070_n N_X_c_1461_n 0.00385303f $X=12.675 $Y=1.985 $X2=0 $Y2=0
cc_863 N_X_c_1285_n N_VGND_c_1573_n 0.0281769f $X=5.8 $Y=0.515 $X2=0 $Y2=0
cc_864 N_X_c_1285_n N_VGND_c_1574_n 0.0282477f $X=5.8 $Y=0.515 $X2=0 $Y2=0
cc_865 N_X_c_1286_n N_VGND_c_1574_n 0.00252612f $X=6.66 $Y=0.515 $X2=0 $Y2=0
cc_866 N_X_c_1286_n N_VGND_c_1575_n 0.0108429f $X=6.66 $Y=0.515 $X2=0 $Y2=0
cc_867 N_X_c_1286_n N_VGND_c_1576_n 0.00287438f $X=6.66 $Y=0.515 $X2=0 $Y2=0
cc_868 N_X_c_1287_n N_VGND_c_1576_n 0.00261701f $X=7.52 $Y=0.515 $X2=0 $Y2=0
cc_869 N_X_c_1287_n N_VGND_c_1577_n 0.0130171f $X=7.52 $Y=0.515 $X2=0 $Y2=0
cc_870 N_X_c_1287_n N_VGND_c_1578_n 0.0302985f $X=7.52 $Y=0.515 $X2=0 $Y2=0
cc_871 N_X_c_1288_n N_VGND_c_1578_n 0.0302985f $X=8.45 $Y=0.515 $X2=0 $Y2=0
cc_872 N_X_c_1288_n N_VGND_c_1579_n 0.00310872f $X=8.45 $Y=0.515 $X2=0 $Y2=0
cc_873 N_X_c_1289_n N_VGND_c_1579_n 0.0298545f $X=9.38 $Y=0.515 $X2=0 $Y2=0
cc_874 N_X_c_1289_n N_VGND_c_1580_n 0.0285298f $X=9.38 $Y=0.515 $X2=0 $Y2=0
cc_875 N_X_c_1290_n N_VGND_c_1580_n 0.0296145f $X=10.31 $Y=0.515 $X2=0 $Y2=0
cc_876 N_X_c_1290_n N_VGND_c_1581_n 0.0294122f $X=10.31 $Y=0.515 $X2=0 $Y2=0
cc_877 N_X_c_1291_n N_VGND_c_1581_n 0.00268474f $X=11.24 $Y=0.515 $X2=0 $Y2=0
cc_878 N_X_c_1291_n N_VGND_c_1582_n 0.0293792f $X=11.24 $Y=0.515 $X2=0 $Y2=0
cc_879 N_X_c_1292_n N_VGND_c_1582_n 0.0294388f $X=12.18 $Y=0.515 $X2=0 $Y2=0
cc_880 N_X_c_1292_n N_VGND_c_1584_n 0.0308109f $X=12.18 $Y=0.515 $X2=0 $Y2=0
cc_881 N_X_c_1285_n N_VGND_c_1593_n 0.0109942f $X=5.8 $Y=0.515 $X2=0 $Y2=0
cc_882 N_X_c_1291_n N_VGND_c_1595_n 0.00950426f $X=11.24 $Y=0.515 $X2=0 $Y2=0
cc_883 N_X_c_1288_n N_VGND_c_1599_n 0.0130022f $X=8.45 $Y=0.515 $X2=0 $Y2=0
cc_884 N_X_c_1289_n N_VGND_c_1600_n 0.0116636f $X=9.38 $Y=0.515 $X2=0 $Y2=0
cc_885 N_X_c_1290_n N_VGND_c_1601_n 0.0109942f $X=10.31 $Y=0.515 $X2=0 $Y2=0
cc_886 N_X_c_1292_n N_VGND_c_1602_n 0.0144922f $X=12.18 $Y=0.515 $X2=0 $Y2=0
cc_887 N_X_c_1285_n N_VGND_c_1610_n 0.00904371f $X=5.8 $Y=0.515 $X2=0 $Y2=0
cc_888 N_X_c_1286_n N_VGND_c_1610_n 0.0089748f $X=6.66 $Y=0.515 $X2=0 $Y2=0
cc_889 N_X_c_1287_n N_VGND_c_1610_n 0.0107298f $X=7.52 $Y=0.515 $X2=0 $Y2=0
cc_890 N_X_c_1288_n N_VGND_c_1610_n 0.0107057f $X=8.45 $Y=0.515 $X2=0 $Y2=0
cc_891 N_X_c_1289_n N_VGND_c_1610_n 0.00959771f $X=9.38 $Y=0.515 $X2=0 $Y2=0
cc_892 N_X_c_1290_n N_VGND_c_1610_n 0.00904371f $X=10.31 $Y=0.515 $X2=0 $Y2=0
cc_893 N_X_c_1291_n N_VGND_c_1610_n 0.0078668f $X=11.24 $Y=0.515 $X2=0 $Y2=0
cc_894 N_X_c_1292_n N_VGND_c_1610_n 0.0118826f $X=12.18 $Y=0.515 $X2=0 $Y2=0
