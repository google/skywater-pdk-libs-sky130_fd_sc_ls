* NGSPICE file created from sky130_fd_sc_ls__maj3_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__maj3_4 A B C VGND VNB VPB VPWR X
M1000 VPWR a_219_392# X VPB phighvt w=1.12e+06u l=150000u
+  ad=2.1282e+12p pd=1.677e+07u as=6.72e+11p ps=5.68e+06u
M1001 a_219_392# B a_501_392# VPB phighvt w=1e+06u l=150000u
+  ad=9.5e+11p pd=7.9e+06u as=6.5e+11p ps=5.3e+06u
M1002 a_219_392# C a_906_78# VNB nshort w=640000u l=150000u
+  ad=5.376e+11p pd=5.52e+06u as=4.45475e+11p ps=4.25e+06u
M1003 X a_219_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_906_78# A VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.2479e+12p ps=1.196e+07u
M1005 a_501_392# B a_219_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_905_392# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=6e+11p pd=5.2e+06u as=0p ps=0u
M1007 VGND C a_504_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=5.41775e+11p ps=4.6e+06u
M1008 a_906_78# C a_219_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A a_906_78# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_219_392# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_219_392# B a_119_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=6.5e+11p ps=5.3e+06u
M1012 VPWR C a_501_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A a_114_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=5.7375e+11p ps=4.61e+06u
M1014 a_119_392# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_219_392# C a_905_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_114_125# B a_219_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_504_125# C VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_905_392# C a_219_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_114_125# A VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_219_392# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.44e+11p ps=4.16e+06u
M1021 VGND a_219_392# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_119_392# B a_219_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_219_392# B a_114_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_504_125# B a_219_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 X a_219_392# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 X a_219_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_501_392# C VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR A a_905_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR A a_119_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_219_392# B a_504_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 X a_219_392# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

