* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dlrbp_1 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_823_98# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VPWR a_642_392# a_823_98# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 a_1342_74# a_823_98# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X3 VPWR a_1342_74# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X4 a_27_142# D VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X5 VPWR GATE a_226_104# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X6 a_753_508# a_823_98# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND a_823_98# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 VGND a_1342_74# Q_N VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 VPWR a_823_98# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X10 a_564_392# a_226_104# a_642_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_642_392# a_226_104# a_775_124# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_823_98# a_642_392# a_1051_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 a_27_142# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X14 a_775_124# a_823_98# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_642_392# a_353_98# a_753_508# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_571_80# a_353_98# a_642_392# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 a_353_98# a_226_104# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 VPWR a_27_142# a_564_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VGND GATE a_226_104# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X20 a_353_98# a_226_104# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 a_1051_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 a_1342_74# a_823_98# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X23 VGND a_27_142# a_571_80# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
