* File: sky130_fd_sc_ls__dlxtn_1.spice
* Created: Wed Sep  2 11:04:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dlxtn_1.pex.spice"
.subckt sky130_fd_sc_ls__dlxtn_1  VNB VPB D GATE_N VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_D_M1004_g N_A_27_115#_M1004_s VNB NSHORT L=0.15 W=0.55
+ AD=0.171896 AS=0.15675 PD=1.33876 PS=1.67 NRD=56.184 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1006 N_A_217_419#_M1006_d N_GATE_N_M1006_g N_VGND_M1004_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.231279 PD=2.05 PS=1.80124 NRD=0 NRS=41.76 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A_217_419#_M1002_g N_A_369_392#_M1002_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.251922 AS=0.2109 PD=1.53899 PS=2.05 NRD=66.48 NRS=0 M=1
+ R=4.93333 SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1015 A_655_79# N_A_27_115#_M1015_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.217878 PD=0.88 PS=1.33101 NRD=12.18 NRS=0.936 M=1 R=4.26667
+ SA=75001.1 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1016 N_A_669_392#_M1016_d N_A_217_419#_M1016_g A_655_79# VNB NSHORT L=0.15
+ W=0.64 AD=0.168211 AS=0.0768 PD=1.52151 PS=0.88 NRD=25.308 NRS=12.18 M=1
+ R=4.26667 SA=75001.4 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1005 A_871_139# N_A_369_392#_M1005_g N_A_669_392#_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.110389 PD=0.66 PS=0.998491 NRD=18.564 NRS=35.712 M=1
+ R=2.8 SA=75001.8 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_863_441#_M1013_g A_871_139# VNB NSHORT L=0.15 W=0.42
+ AD=0.0930736 AS=0.0504 PD=0.832075 PS=0.66 NRD=37.848 NRS=18.564 M=1 R=2.8
+ SA=75002.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1014 N_A_863_441#_M1014_d N_A_669_392#_M1014_g N_VGND_M1013_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.141826 PD=1.85 PS=1.26792 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75001.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_Q_M1001_d N_A_863_441#_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2146 AS=0.2109 PD=2.06 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_D_M1010_g N_A_27_115#_M1010_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.147 AS=0.2478 PD=1.19 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1011 N_A_217_419#_M1011_d N_GATE_N_M1011_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.3192 AS=0.147 PD=2.44 PS=1.19 NRD=22.261 NRS=2.3443 M=1 R=5.6
+ SA=75000.7 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A_217_419#_M1003_g N_A_369_392#_M1003_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.23294 AS=0.2478 PD=1.47457 PS=2.27 NRD=52.1262 NRS=2.3443
+ M=1 R=5.6 SA=75000.2 SB=75002 A=0.126 P=1.98 MULT=1
MM1012 A_585_392# N_A_27_115#_M1012_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.27731 PD=1.27 PS=1.75543 NRD=15.7403 NRS=21.6503 M=1 R=6.66667
+ SA=75000.8 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1008 N_A_669_392#_M1008_d N_A_369_392#_M1008_g A_585_392# VPB PHIGHVT L=0.15
+ W=1 AD=0.361127 AS=0.135 PD=2.20423 PS=1.27 NRD=19.7 NRS=15.7403 M=1 R=6.66667
+ SA=75001.2 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1000 A_812_508# N_A_217_419#_M1000_g N_A_669_392#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.151673 PD=0.69 PS=0.925775 NRD=37.5088 NRS=89.1031 M=1
+ R=2.8 SA=75001.8 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1017 N_VPWR_M1017_d N_A_863_441#_M1017_g A_812_508# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.131354 AS=0.0567 PD=0.976056 PS=0.69 NRD=7.0329 NRS=37.5088 M=1 R=2.8
+ SA=75002.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1007 N_A_863_441#_M1007_d N_A_669_392#_M1007_g N_VPWR_M1017_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.312746 PD=2.59 PS=2.32394 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75001.4 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1009 N_Q_M1009_d N_A_863_441#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX18_noxref VNB VPB NWDIODE A=13.206 P=17.92
c_72 VNB 0 4.76483e-20 $X=0 $Y=0
c_928 A_655_79# 0 3.15497e-20 $X=3.275 $Y=0.395
*
.include "sky130_fd_sc_ls__dlxtn_1.pxi.spice"
*
.ends
*
*
