* File: sky130_fd_sc_ls__bufinv_8.pxi.spice
* Created: Fri Aug 28 13:08:15 2020
* 
x_PM_SKY130_FD_SC_LS__BUFINV_8%A N_A_c_106_n N_A_M1013_g N_A_M1021_g A
+ N_A_c_108_n PM_SKY130_FD_SC_LS__BUFINV_8%A
x_PM_SKY130_FD_SC_LS__BUFINV_8%A_183_48# N_A_183_48#_M1004_d N_A_183_48#_M1012_d
+ N_A_183_48#_M1014_d N_A_183_48#_M1023_d N_A_183_48#_M1001_g
+ N_A_183_48#_c_153_n N_A_183_48#_M1000_g N_A_183_48#_M1003_g
+ N_A_183_48#_c_154_n N_A_183_48#_M1002_g N_A_183_48#_c_155_n
+ N_A_183_48#_M1006_g N_A_183_48#_M1005_g N_A_183_48#_c_156_n
+ N_A_183_48#_M1007_g N_A_183_48#_M1009_g N_A_183_48#_c_157_n
+ N_A_183_48#_M1010_g N_A_183_48#_M1011_g N_A_183_48#_c_158_n
+ N_A_183_48#_M1016_g N_A_183_48#_M1015_g N_A_183_48#_c_159_n
+ N_A_183_48#_M1019_g N_A_183_48#_M1017_g N_A_183_48#_c_160_n
+ N_A_183_48#_M1022_g N_A_183_48#_M1020_g N_A_183_48#_c_144_n
+ N_A_183_48#_c_145_n N_A_183_48#_c_146_n N_A_183_48#_c_147_n
+ N_A_183_48#_c_148_n N_A_183_48#_c_176_p N_A_183_48#_c_149_n
+ N_A_183_48#_c_150_n N_A_183_48#_c_162_n N_A_183_48#_c_163_n
+ N_A_183_48#_c_151_n N_A_183_48#_c_164_n N_A_183_48#_c_152_n
+ PM_SKY130_FD_SC_LS__BUFINV_8%A_183_48#
x_PM_SKY130_FD_SC_LS__BUFINV_8%A_27_368# N_A_27_368#_M1021_s N_A_27_368#_M1013_s
+ N_A_27_368#_c_371_n N_A_27_368#_M1014_g N_A_27_368#_M1004_g
+ N_A_27_368#_c_372_n N_A_27_368#_M1018_g N_A_27_368#_M1008_g
+ N_A_27_368#_c_373_n N_A_27_368#_M1023_g N_A_27_368#_M1012_g
+ N_A_27_368#_c_374_n N_A_27_368#_c_365_n N_A_27_368#_c_366_n
+ N_A_27_368#_c_367_n N_A_27_368#_c_388_n N_A_27_368#_c_368_n
+ N_A_27_368#_c_422_n N_A_27_368#_c_433_n N_A_27_368#_c_376_n
+ N_A_27_368#_c_377_n N_A_27_368#_c_378_n N_A_27_368#_c_457_p
+ N_A_27_368#_c_369_n N_A_27_368#_c_370_n PM_SKY130_FD_SC_LS__BUFINV_8%A_27_368#
x_PM_SKY130_FD_SC_LS__BUFINV_8%VPWR N_VPWR_M1013_d N_VPWR_M1002_s N_VPWR_M1007_s
+ N_VPWR_M1016_s N_VPWR_M1022_s N_VPWR_M1018_s N_VPWR_c_515_n N_VPWR_c_516_n
+ N_VPWR_c_517_n N_VPWR_c_518_n N_VPWR_c_519_n N_VPWR_c_520_n N_VPWR_c_521_n
+ N_VPWR_c_522_n VPWR N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_525_n
+ N_VPWR_c_526_n N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_514_n N_VPWR_c_530_n
+ N_VPWR_c_531_n N_VPWR_c_532_n N_VPWR_c_533_n N_VPWR_c_534_n
+ PM_SKY130_FD_SC_LS__BUFINV_8%VPWR
x_PM_SKY130_FD_SC_LS__BUFINV_8%Y N_Y_M1001_d N_Y_M1005_d N_Y_M1011_d N_Y_M1017_d
+ N_Y_M1000_d N_Y_M1006_d N_Y_M1010_d N_Y_M1019_d N_Y_c_613_n N_Y_c_622_n
+ N_Y_c_614_n N_Y_c_615_n N_Y_c_616_n N_Y_c_617_n N_Y_c_618_n N_Y_c_657_n
+ N_Y_c_619_n N_Y_c_620_n Y Y Y Y PM_SKY130_FD_SC_LS__BUFINV_8%Y
x_PM_SKY130_FD_SC_LS__BUFINV_8%VGND N_VGND_M1021_d N_VGND_M1003_s N_VGND_M1009_s
+ N_VGND_M1015_s N_VGND_M1020_s N_VGND_M1008_s N_VGND_c_715_n N_VGND_c_716_n
+ N_VGND_c_717_n N_VGND_c_718_n N_VGND_c_719_n N_VGND_c_720_n VGND
+ N_VGND_c_721_n N_VGND_c_722_n N_VGND_c_723_n N_VGND_c_724_n N_VGND_c_725_n
+ N_VGND_c_726_n N_VGND_c_727_n N_VGND_c_728_n N_VGND_c_729_n N_VGND_c_730_n
+ N_VGND_c_731_n N_VGND_c_732_n N_VGND_c_733_n N_VGND_c_734_n
+ PM_SKY130_FD_SC_LS__BUFINV_8%VGND
cc_1 VNB N_A_c_106_n 0.0340423f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_A_M1021_g 0.0327781f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_3 VNB N_A_c_108_n 0.0147537f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_4 VNB N_A_183_48#_M1001_g 0.0215966f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_5 VNB N_A_183_48#_M1003_g 0.0213269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_183_48#_M1005_g 0.0211937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_183_48#_M1009_g 0.0212282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_183_48#_M1011_g 0.0217898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_183_48#_M1015_g 0.0217898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_183_48#_M1017_g 0.022104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_183_48#_M1020_g 0.0231611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_183_48#_c_144_n 0.0086775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_183_48#_c_145_n 0.00197374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_183_48#_c_146_n 0.00209186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_183_48#_c_147_n 0.00496443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_183_48#_c_148_n 0.003141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_183_48#_c_149_n 0.0227723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_183_48#_c_150_n 0.0220728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_183_48#_c_151_n 0.0104445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_183_48#_c_152_n 0.22295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_368#_M1004_g 0.0216729f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_22 VNB N_A_27_368#_M1008_g 0.022431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_368#_M1012_g 0.0287448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_368#_c_365_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_368#_c_366_n 0.00538315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_368#_c_367_n 0.00909915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_368#_c_368_n 0.00862727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_368#_c_369_n 0.00269557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_368#_c_370_n 0.0801452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_514_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_613_n 0.00381057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_614_n 0.00195975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_615_n 0.00309972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_616_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_617_n 0.0053906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_618_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_619_n 0.00145912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_620_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB Y 0.00257348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_715_n 0.00571296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_716_n 0.00498656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_717_n 0.00498656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_718_n 0.00516528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_719_n 0.00500818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_720_n 0.00570743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_721_n 0.0178682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_722_n 0.0186748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_723_n 0.0150174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_724_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_725_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_726_n 0.0153775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_727_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_728_n 0.345062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_729_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_730_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_731_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_732_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_733_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_734_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VPB N_A_c_106_n 0.0355825f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_61 VPB N_A_c_108_n 0.00743971f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_62 VPB N_A_183_48#_c_153_n 0.0152291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_183_48#_c_154_n 0.0145806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_183_48#_c_155_n 0.0147204f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_183_48#_c_156_n 0.014741f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_183_48#_c_157_n 0.014741f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_183_48#_c_158_n 0.014741f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_183_48#_c_159_n 0.0156967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_183_48#_c_160_n 0.0163631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_183_48#_c_150_n 0.018854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_183_48#_c_162_n 0.0275864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_183_48#_c_163_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_183_48#_c_164_n 0.00704942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_183_48#_c_152_n 0.0519406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_27_368#_c_371_n 0.0158492f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_27_368#_c_372_n 0.0153274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_27_368#_c_373_n 0.0193831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_27_368#_c_374_n 0.0243843f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_27_368#_c_368_n 0.00331088f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_27_368#_c_376_n 0.00266721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_27_368#_c_377_n 0.00195961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_27_368#_c_378_n 0.0179584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_27_368#_c_369_n 0.0027421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_27_368#_c_370_n 0.0198344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_515_n 0.00584464f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_516_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_517_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_518_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_519_n 0.00581944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_520_n 0.00581944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_521_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_522_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_523_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_524_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_525_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_526_n 0.0218958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_527_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_528_n 0.017793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_514_n 0.111893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_530_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_531_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_532_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_533_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_534_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_Y_c_622_n 0.0121156f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 N_A_M1021_g N_A_183_48#_M1001_g 0.0228206f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_c_106_n N_A_183_48#_c_153_n 0.0324428f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A_c_106_n N_A_183_48#_c_152_n 0.0139152f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_109 N_A_c_106_n N_A_27_368#_c_374_n 0.00747601f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A_M1021_g N_A_27_368#_c_365_n 0.00159319f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A_c_106_n N_A_27_368#_c_366_n 7.7117e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_112 N_A_M1021_g N_A_27_368#_c_366_n 0.0146818f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A_c_108_n N_A_27_368#_c_366_n 0.012562f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A_c_106_n N_A_27_368#_c_367_n 0.00126636f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_115 N_A_c_108_n N_A_27_368#_c_367_n 0.0219605f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_116 N_A_c_106_n N_A_27_368#_c_388_n 0.014804f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A_c_108_n N_A_27_368#_c_388_n 0.00339179f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_118 N_A_c_106_n N_A_27_368#_c_368_n 0.00919461f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A_M1021_g N_A_27_368#_c_368_n 0.00374261f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A_c_108_n N_A_27_368#_c_368_n 0.0329132f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_121 N_A_c_106_n N_A_27_368#_c_378_n 0.0054792f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A_c_108_n N_A_27_368#_c_378_n 0.0255473f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_123 N_A_c_106_n N_VPWR_c_515_n 0.00532643f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A_c_106_n N_VPWR_c_523_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A_c_106_n N_VPWR_c_514_n 0.00860926f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A_M1021_g Y 3.41373e-19 $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A_M1021_g Y 6.75874e-19 $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A_M1021_g N_VGND_c_715_n 0.0132976f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A_M1021_g N_VGND_c_721_n 0.00383152f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_M1021_g N_VGND_c_728_n 0.00761248f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A_183_48#_c_160_n N_A_27_368#_c_371_n 0.0328539f $X=4.285 $Y=1.765
+ $X2=0 $Y2=0
cc_132 N_A_183_48#_c_163_n N_A_27_368#_c_371_n 0.0123186f $X=5.01 $Y=2.305 $X2=0
+ $Y2=0
cc_133 N_A_183_48#_M1020_g N_A_27_368#_M1004_g 0.0189988f $X=4.3 $Y=0.74 $X2=0
+ $Y2=0
cc_134 N_A_183_48#_c_144_n N_A_27_368#_M1004_g 7.44057e-19 $X=4.65 $Y=1.465
+ $X2=0 $Y2=0
cc_135 N_A_183_48#_c_145_n N_A_27_368#_M1004_g 0.00529113f $X=4.735 $Y=1.3 $X2=0
+ $Y2=0
cc_136 N_A_183_48#_c_146_n N_A_27_368#_M1004_g 4.16154e-19 $X=5.02 $Y=0.515
+ $X2=0 $Y2=0
cc_137 N_A_183_48#_c_148_n N_A_27_368#_M1004_g 0.0132227f $X=5.125 $Y=1.005
+ $X2=0 $Y2=0
cc_138 N_A_183_48#_c_176_p N_A_27_368#_c_372_n 0.0122751f $X=5.795 $Y=2.225
+ $X2=0 $Y2=0
cc_139 N_A_183_48#_c_150_n N_A_27_368#_c_372_n 9.31641e-19 $X=5.96 $Y=1.985
+ $X2=0 $Y2=0
cc_140 N_A_183_48#_c_163_n N_A_27_368#_c_372_n 0.0103638f $X=5.01 $Y=2.305 $X2=0
+ $Y2=0
cc_141 N_A_183_48#_c_145_n N_A_27_368#_M1008_g 9.46656e-19 $X=4.735 $Y=1.3 $X2=0
+ $Y2=0
cc_142 N_A_183_48#_c_146_n N_A_27_368#_M1008_g 4.16154e-19 $X=5.02 $Y=0.515
+ $X2=0 $Y2=0
cc_143 N_A_183_48#_c_147_n N_A_27_368#_M1008_g 0.0153525f $X=5.795 $Y=1.005
+ $X2=0 $Y2=0
cc_144 N_A_183_48#_c_149_n N_A_27_368#_M1008_g 5.56882e-19 $X=5.96 $Y=0.515
+ $X2=0 $Y2=0
cc_145 N_A_183_48#_c_150_n N_A_27_368#_M1008_g 8.9077e-19 $X=5.96 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A_183_48#_c_176_p N_A_27_368#_c_373_n 0.015945f $X=5.795 $Y=2.225 $X2=0
+ $Y2=0
cc_147 N_A_183_48#_c_150_n N_A_27_368#_c_373_n 0.0066695f $X=5.96 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A_183_48#_c_162_n N_A_27_368#_c_373_n 9.4299e-19 $X=5.96 $Y=2.4 $X2=0
+ $Y2=0
cc_149 N_A_183_48#_c_163_n N_A_27_368#_c_373_n 6.32426e-19 $X=5.01 $Y=2.305
+ $X2=0 $Y2=0
cc_150 N_A_183_48#_c_164_n N_A_27_368#_c_373_n 0.00141023f $X=5.96 $Y=2.225
+ $X2=0 $Y2=0
cc_151 N_A_183_48#_c_147_n N_A_27_368#_M1012_g 0.0176987f $X=5.795 $Y=1.005
+ $X2=0 $Y2=0
cc_152 N_A_183_48#_c_149_n N_A_27_368#_M1012_g 0.00889319f $X=5.96 $Y=0.515
+ $X2=0 $Y2=0
cc_153 N_A_183_48#_c_150_n N_A_27_368#_M1012_g 0.00744164f $X=5.96 $Y=1.985
+ $X2=0 $Y2=0
cc_154 N_A_183_48#_c_151_n N_A_27_368#_M1012_g 9.50735e-19 $X=5.96 $Y=1.005
+ $X2=0 $Y2=0
cc_155 N_A_183_48#_M1001_g N_A_27_368#_c_366_n 0.00116372f $X=0.99 $Y=0.74 $X2=0
+ $Y2=0
cc_156 N_A_183_48#_M1001_g N_A_27_368#_c_368_n 0.00543775f $X=0.99 $Y=0.74 $X2=0
+ $Y2=0
cc_157 N_A_183_48#_c_153_n N_A_27_368#_c_368_n 0.00270815f $X=1.005 $Y=1.765
+ $X2=0 $Y2=0
cc_158 N_A_183_48#_c_153_n N_A_27_368#_c_422_n 0.0190541f $X=1.005 $Y=1.765
+ $X2=0 $Y2=0
cc_159 N_A_183_48#_c_154_n N_A_27_368#_c_422_n 0.0148716f $X=1.455 $Y=1.765
+ $X2=0 $Y2=0
cc_160 N_A_183_48#_c_155_n N_A_27_368#_c_422_n 0.0148856f $X=1.905 $Y=1.765
+ $X2=0 $Y2=0
cc_161 N_A_183_48#_c_156_n N_A_27_368#_c_422_n 0.0148856f $X=2.355 $Y=1.765
+ $X2=0 $Y2=0
cc_162 N_A_183_48#_c_157_n N_A_27_368#_c_422_n 0.0148856f $X=2.805 $Y=1.765
+ $X2=0 $Y2=0
cc_163 N_A_183_48#_c_158_n N_A_27_368#_c_422_n 0.0148856f $X=3.255 $Y=1.765
+ $X2=0 $Y2=0
cc_164 N_A_183_48#_c_159_n N_A_27_368#_c_422_n 0.0155265f $X=3.705 $Y=1.765
+ $X2=0 $Y2=0
cc_165 N_A_183_48#_c_160_n N_A_27_368#_c_422_n 0.016981f $X=4.285 $Y=1.765 $X2=0
+ $Y2=0
cc_166 N_A_183_48#_c_144_n N_A_27_368#_c_422_n 0.00388353f $X=4.65 $Y=1.465
+ $X2=0 $Y2=0
cc_167 N_A_183_48#_c_163_n N_A_27_368#_c_422_n 0.00976109f $X=5.01 $Y=2.305
+ $X2=0 $Y2=0
cc_168 N_A_183_48#_c_152_n N_A_27_368#_c_422_n 6.90209e-19 $X=4.285 $Y=1.532
+ $X2=0 $Y2=0
cc_169 N_A_183_48#_c_163_n N_A_27_368#_c_433_n 0.00531806f $X=5.01 $Y=2.305
+ $X2=0 $Y2=0
cc_170 N_A_183_48#_M1014_d N_A_27_368#_c_376_n 0.00108773f $X=4.86 $Y=1.84 $X2=0
+ $Y2=0
cc_171 N_A_183_48#_c_144_n N_A_27_368#_c_376_n 0.0198373f $X=4.65 $Y=1.465 $X2=0
+ $Y2=0
cc_172 N_A_183_48#_c_148_n N_A_27_368#_c_376_n 0.00468499f $X=5.125 $Y=1.005
+ $X2=0 $Y2=0
cc_173 N_A_183_48#_c_163_n N_A_27_368#_c_376_n 0.00703968f $X=5.01 $Y=2.305
+ $X2=0 $Y2=0
cc_174 N_A_183_48#_c_160_n N_A_27_368#_c_377_n 0.00108028f $X=4.285 $Y=1.765
+ $X2=0 $Y2=0
cc_175 N_A_183_48#_c_144_n N_A_27_368#_c_377_n 0.01491f $X=4.65 $Y=1.465 $X2=0
+ $Y2=0
cc_176 N_A_183_48#_c_153_n N_A_27_368#_c_378_n 9.07821e-19 $X=1.005 $Y=1.765
+ $X2=0 $Y2=0
cc_177 N_A_183_48#_M1014_d N_A_27_368#_c_369_n 0.00154606f $X=4.86 $Y=1.84 $X2=0
+ $Y2=0
cc_178 N_A_183_48#_c_144_n N_A_27_368#_c_369_n 0.0259125f $X=4.65 $Y=1.465 $X2=0
+ $Y2=0
cc_179 N_A_183_48#_c_148_n N_A_27_368#_c_369_n 0.0455162f $X=5.125 $Y=1.005
+ $X2=0 $Y2=0
cc_180 N_A_183_48#_c_176_p N_A_27_368#_c_369_n 0.0293407f $X=5.795 $Y=2.225
+ $X2=0 $Y2=0
cc_181 N_A_183_48#_c_150_n N_A_27_368#_c_369_n 0.0427207f $X=5.96 $Y=1.985 $X2=0
+ $Y2=0
cc_182 N_A_183_48#_c_163_n N_A_27_368#_c_369_n 0.0112875f $X=5.01 $Y=2.305 $X2=0
+ $Y2=0
cc_183 N_A_183_48#_c_152_n N_A_27_368#_c_369_n 2.29472e-19 $X=4.285 $Y=1.532
+ $X2=0 $Y2=0
cc_184 N_A_183_48#_c_144_n N_A_27_368#_c_370_n 0.0135218f $X=4.65 $Y=1.465 $X2=0
+ $Y2=0
cc_185 N_A_183_48#_c_147_n N_A_27_368#_c_370_n 0.0012067f $X=5.795 $Y=1.005
+ $X2=0 $Y2=0
cc_186 N_A_183_48#_c_148_n N_A_27_368#_c_370_n 0.00135251f $X=5.125 $Y=1.005
+ $X2=0 $Y2=0
cc_187 N_A_183_48#_c_176_p N_A_27_368#_c_370_n 9.27004e-19 $X=5.795 $Y=2.225
+ $X2=0 $Y2=0
cc_188 N_A_183_48#_c_150_n N_A_27_368#_c_370_n 0.0166242f $X=5.96 $Y=1.985 $X2=0
+ $Y2=0
cc_189 N_A_183_48#_c_163_n N_A_27_368#_c_370_n 6.80003e-19 $X=5.01 $Y=2.305
+ $X2=0 $Y2=0
cc_190 N_A_183_48#_c_152_n N_A_27_368#_c_370_n 0.0235998f $X=4.285 $Y=1.532
+ $X2=0 $Y2=0
cc_191 N_A_183_48#_c_176_p N_VPWR_M1018_s 0.00473156f $X=5.795 $Y=2.225 $X2=0
+ $Y2=0
cc_192 N_A_183_48#_c_153_n N_VPWR_c_515_n 0.0112251f $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_A_183_48#_c_154_n N_VPWR_c_515_n 0.0015077f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_194 N_A_183_48#_c_153_n N_VPWR_c_516_n 0.0015077f $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A_183_48#_c_154_n N_VPWR_c_516_n 0.0112999f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_196 N_A_183_48#_c_155_n N_VPWR_c_516_n 0.0112999f $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_A_183_48#_c_156_n N_VPWR_c_516_n 0.0015077f $X=2.355 $Y=1.765 $X2=0
+ $Y2=0
cc_198 N_A_183_48#_c_155_n N_VPWR_c_517_n 0.0015077f $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_199 N_A_183_48#_c_156_n N_VPWR_c_517_n 0.0112999f $X=2.355 $Y=1.765 $X2=0
+ $Y2=0
cc_200 N_A_183_48#_c_157_n N_VPWR_c_517_n 0.0112999f $X=2.805 $Y=1.765 $X2=0
+ $Y2=0
cc_201 N_A_183_48#_c_158_n N_VPWR_c_517_n 0.0015077f $X=3.255 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_A_183_48#_c_157_n N_VPWR_c_518_n 0.0015077f $X=2.805 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_A_183_48#_c_158_n N_VPWR_c_518_n 0.0112999f $X=3.255 $Y=1.765 $X2=0
+ $Y2=0
cc_204 N_A_183_48#_c_159_n N_VPWR_c_518_n 0.0124787f $X=3.705 $Y=1.765 $X2=0
+ $Y2=0
cc_205 N_A_183_48#_c_160_n N_VPWR_c_518_n 0.00228588f $X=4.285 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_A_183_48#_c_159_n N_VPWR_c_519_n 0.00228588f $X=3.705 $Y=1.765 $X2=0
+ $Y2=0
cc_207 N_A_183_48#_c_160_n N_VPWR_c_519_n 0.0124039f $X=4.285 $Y=1.765 $X2=0
+ $Y2=0
cc_208 N_A_183_48#_c_163_n N_VPWR_c_519_n 0.0157994f $X=5.01 $Y=2.305 $X2=0
+ $Y2=0
cc_209 N_A_183_48#_c_176_p N_VPWR_c_520_n 0.0202249f $X=5.795 $Y=2.225 $X2=0
+ $Y2=0
cc_210 N_A_183_48#_c_162_n N_VPWR_c_520_n 0.0195323f $X=5.96 $Y=2.4 $X2=0 $Y2=0
cc_211 N_A_183_48#_c_163_n N_VPWR_c_520_n 0.0195517f $X=5.01 $Y=2.305 $X2=0
+ $Y2=0
cc_212 N_A_183_48#_c_157_n N_VPWR_c_521_n 0.00413917f $X=2.805 $Y=1.765 $X2=0
+ $Y2=0
cc_213 N_A_183_48#_c_158_n N_VPWR_c_521_n 0.00413917f $X=3.255 $Y=1.765 $X2=0
+ $Y2=0
cc_214 N_A_183_48#_c_153_n N_VPWR_c_524_n 0.00413917f $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_215 N_A_183_48#_c_154_n N_VPWR_c_524_n 0.00413917f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_216 N_A_183_48#_c_155_n N_VPWR_c_525_n 0.00413917f $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_217 N_A_183_48#_c_156_n N_VPWR_c_525_n 0.00413917f $X=2.355 $Y=1.765 $X2=0
+ $Y2=0
cc_218 N_A_183_48#_c_159_n N_VPWR_c_526_n 0.00413917f $X=3.705 $Y=1.765 $X2=0
+ $Y2=0
cc_219 N_A_183_48#_c_160_n N_VPWR_c_526_n 0.00413917f $X=4.285 $Y=1.765 $X2=0
+ $Y2=0
cc_220 N_A_183_48#_c_163_n N_VPWR_c_527_n 0.014552f $X=5.01 $Y=2.305 $X2=0 $Y2=0
cc_221 N_A_183_48#_c_162_n N_VPWR_c_528_n 0.0124046f $X=5.96 $Y=2.4 $X2=0 $Y2=0
cc_222 N_A_183_48#_c_153_n N_VPWR_c_514_n 0.00817726f $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_223 N_A_183_48#_c_154_n N_VPWR_c_514_n 0.00817726f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_224 N_A_183_48#_c_155_n N_VPWR_c_514_n 0.00817726f $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_225 N_A_183_48#_c_156_n N_VPWR_c_514_n 0.00817726f $X=2.355 $Y=1.765 $X2=0
+ $Y2=0
cc_226 N_A_183_48#_c_157_n N_VPWR_c_514_n 0.00817726f $X=2.805 $Y=1.765 $X2=0
+ $Y2=0
cc_227 N_A_183_48#_c_158_n N_VPWR_c_514_n 0.00817726f $X=3.255 $Y=1.765 $X2=0
+ $Y2=0
cc_228 N_A_183_48#_c_159_n N_VPWR_c_514_n 0.00818839f $X=3.705 $Y=1.765 $X2=0
+ $Y2=0
cc_229 N_A_183_48#_c_160_n N_VPWR_c_514_n 0.00818839f $X=4.285 $Y=1.765 $X2=0
+ $Y2=0
cc_230 N_A_183_48#_c_162_n N_VPWR_c_514_n 0.0102675f $X=5.96 $Y=2.4 $X2=0 $Y2=0
cc_231 N_A_183_48#_c_163_n N_VPWR_c_514_n 0.0119791f $X=5.01 $Y=2.305 $X2=0
+ $Y2=0
cc_232 N_A_183_48#_M1003_g N_Y_c_613_n 0.0154892f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A_183_48#_M1005_g N_Y_c_613_n 0.0152302f $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A_183_48#_c_144_n N_Y_c_613_n 0.0299541f $X=4.65 $Y=1.465 $X2=0 $Y2=0
cc_235 N_A_183_48#_c_152_n N_Y_c_613_n 0.00416906f $X=4.285 $Y=1.532 $X2=0 $Y2=0
cc_236 N_A_183_48#_c_154_n N_Y_c_622_n 0.0127934f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A_183_48#_c_155_n N_Y_c_622_n 0.0118134f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A_183_48#_c_156_n N_Y_c_622_n 0.0118134f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A_183_48#_c_157_n N_Y_c_622_n 0.0118134f $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_240 N_A_183_48#_c_158_n N_Y_c_622_n 0.0118134f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A_183_48#_c_159_n N_Y_c_622_n 0.0157826f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A_183_48#_c_160_n N_Y_c_622_n 0.00741334f $X=4.285 $Y=1.765 $X2=0 $Y2=0
cc_243 N_A_183_48#_c_144_n N_Y_c_622_n 0.196358f $X=4.65 $Y=1.465 $X2=0 $Y2=0
cc_244 N_A_183_48#_c_152_n N_Y_c_622_n 0.0495179f $X=4.285 $Y=1.532 $X2=0 $Y2=0
cc_245 N_A_183_48#_M1005_g N_Y_c_614_n 3.99083e-19 $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A_183_48#_M1009_g N_Y_c_614_n 3.99083e-19 $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A_183_48#_M1009_g N_Y_c_615_n 0.0152302f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A_183_48#_M1011_g N_Y_c_615_n 0.01369f $X=2.87 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A_183_48#_c_144_n N_Y_c_615_n 0.0507189f $X=4.65 $Y=1.465 $X2=0 $Y2=0
cc_250 N_A_183_48#_c_152_n N_Y_c_615_n 0.00384615f $X=4.285 $Y=1.532 $X2=0 $Y2=0
cc_251 N_A_183_48#_M1009_g N_Y_c_616_n 5.56882e-19 $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_183_48#_M1011_g N_Y_c_616_n 0.0082419f $X=2.87 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_183_48#_M1015_g N_Y_c_616_n 0.00746139f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_183_48#_M1017_g N_Y_c_616_n 3.52398e-19 $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_183_48#_M1015_g N_Y_c_617_n 0.0115433f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A_183_48#_M1017_g N_Y_c_617_n 0.0151263f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A_183_48#_M1020_g N_Y_c_617_n 0.00323816f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A_183_48#_c_144_n N_Y_c_617_n 0.0769774f $X=4.65 $Y=1.465 $X2=0 $Y2=0
cc_259 N_A_183_48#_c_148_n N_Y_c_617_n 0.00764154f $X=5.125 $Y=1.005 $X2=0 $Y2=0
cc_260 N_A_183_48#_c_152_n N_Y_c_617_n 0.00781614f $X=4.285 $Y=1.532 $X2=0 $Y2=0
cc_261 N_A_183_48#_M1017_g N_Y_c_618_n 0.00324276f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_183_48#_M1020_g N_Y_c_618_n 0.00946516f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_183_48#_c_148_n N_Y_c_618_n 0.00335458f $X=5.125 $Y=1.005 $X2=0 $Y2=0
cc_264 N_A_183_48#_c_153_n N_Y_c_657_n 0.00343694f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_265 N_A_183_48#_c_154_n N_Y_c_657_n 8.42227e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_266 N_A_183_48#_c_144_n N_Y_c_619_n 0.0160251f $X=4.65 $Y=1.465 $X2=0 $Y2=0
cc_267 N_A_183_48#_c_152_n N_Y_c_619_n 0.00232957f $X=4.285 $Y=1.532 $X2=0 $Y2=0
cc_268 N_A_183_48#_M1011_g N_Y_c_620_n 0.00115621f $X=2.87 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_183_48#_M1015_g N_Y_c_620_n 0.00257766f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_270 N_A_183_48#_M1017_g N_Y_c_620_n 2.50354e-19 $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A_183_48#_c_144_n N_Y_c_620_n 0.0276081f $X=4.65 $Y=1.465 $X2=0 $Y2=0
cc_272 N_A_183_48#_c_152_n N_Y_c_620_n 0.00232957f $X=4.285 $Y=1.532 $X2=0 $Y2=0
cc_273 N_A_183_48#_M1001_g Y 0.00600697f $X=0.99 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A_183_48#_M1003_g Y 0.00829833f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_275 N_A_183_48#_M1005_g Y 5.00623e-19 $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A_183_48#_M1001_g Y 0.00377972f $X=0.99 $Y=0.74 $X2=0 $Y2=0
cc_277 N_A_183_48#_M1003_g Y 8.07377e-19 $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_278 N_A_183_48#_M1001_g Y 0.00361253f $X=0.99 $Y=0.74 $X2=0 $Y2=0
cc_279 N_A_183_48#_c_153_n Y 7.4672e-19 $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_280 N_A_183_48#_M1003_g Y 0.00538497f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_281 N_A_183_48#_c_154_n Y 9.96548e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_282 N_A_183_48#_M1005_g Y 7.96256e-19 $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A_183_48#_c_144_n Y 0.0177955f $X=4.65 $Y=1.465 $X2=0 $Y2=0
cc_284 N_A_183_48#_c_152_n Y 0.0363429f $X=4.285 $Y=1.532 $X2=0 $Y2=0
cc_285 N_A_183_48#_c_148_n N_VGND_M1020_s 0.00318074f $X=5.125 $Y=1.005 $X2=0
+ $Y2=0
cc_286 N_A_183_48#_c_147_n N_VGND_M1008_s 0.00253871f $X=5.795 $Y=1.005 $X2=0
+ $Y2=0
cc_287 N_A_183_48#_M1001_g N_VGND_c_715_n 0.00233397f $X=0.99 $Y=0.74 $X2=0
+ $Y2=0
cc_288 N_A_183_48#_M1003_g N_VGND_c_716_n 0.00365073f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_289 N_A_183_48#_M1005_g N_VGND_c_716_n 0.00799341f $X=1.94 $Y=0.74 $X2=0
+ $Y2=0
cc_290 N_A_183_48#_M1009_g N_VGND_c_716_n 4.27258e-19 $X=2.37 $Y=0.74 $X2=0
+ $Y2=0
cc_291 N_A_183_48#_M1005_g N_VGND_c_717_n 4.27258e-19 $X=1.94 $Y=0.74 $X2=0
+ $Y2=0
cc_292 N_A_183_48#_M1009_g N_VGND_c_717_n 0.00792092f $X=2.37 $Y=0.74 $X2=0
+ $Y2=0
cc_293 N_A_183_48#_M1011_g N_VGND_c_717_n 0.00365073f $X=2.87 $Y=0.74 $X2=0
+ $Y2=0
cc_294 N_A_183_48#_M1015_g N_VGND_c_718_n 0.00406778f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_295 N_A_183_48#_M1017_g N_VGND_c_718_n 0.00979254f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_296 N_A_183_48#_M1020_g N_VGND_c_718_n 4.87331e-19 $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_297 N_A_183_48#_M1020_g N_VGND_c_719_n 0.00365073f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_298 N_A_183_48#_c_144_n N_VGND_c_719_n 0.00785549f $X=4.65 $Y=1.465 $X2=0
+ $Y2=0
cc_299 N_A_183_48#_c_146_n N_VGND_c_719_n 0.0142435f $X=5.02 $Y=0.515 $X2=0
+ $Y2=0
cc_300 N_A_183_48#_c_148_n N_VGND_c_719_n 0.00333948f $X=5.125 $Y=1.005 $X2=0
+ $Y2=0
cc_301 N_A_183_48#_c_146_n N_VGND_c_720_n 0.0142435f $X=5.02 $Y=0.515 $X2=0
+ $Y2=0
cc_302 N_A_183_48#_c_147_n N_VGND_c_720_n 0.0215485f $X=5.795 $Y=1.005 $X2=0
+ $Y2=0
cc_303 N_A_183_48#_c_149_n N_VGND_c_720_n 0.0142986f $X=5.96 $Y=0.515 $X2=0
+ $Y2=0
cc_304 N_A_183_48#_M1001_g N_VGND_c_722_n 0.00456932f $X=0.99 $Y=0.74 $X2=0
+ $Y2=0
cc_305 N_A_183_48#_M1003_g N_VGND_c_722_n 0.00434272f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_306 N_A_183_48#_M1005_g N_VGND_c_723_n 0.00383152f $X=1.94 $Y=0.74 $X2=0
+ $Y2=0
cc_307 N_A_183_48#_M1009_g N_VGND_c_723_n 0.00383152f $X=2.37 $Y=0.74 $X2=0
+ $Y2=0
cc_308 N_A_183_48#_M1011_g N_VGND_c_724_n 0.00434272f $X=2.87 $Y=0.74 $X2=0
+ $Y2=0
cc_309 N_A_183_48#_M1015_g N_VGND_c_724_n 0.00434272f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_310 N_A_183_48#_M1017_g N_VGND_c_725_n 0.00383152f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_311 N_A_183_48#_M1020_g N_VGND_c_725_n 0.00434272f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A_183_48#_c_146_n N_VGND_c_726_n 0.00889602f $X=5.02 $Y=0.515 $X2=0
+ $Y2=0
cc_313 N_A_183_48#_c_149_n N_VGND_c_727_n 0.0145639f $X=5.96 $Y=0.515 $X2=0
+ $Y2=0
cc_314 N_A_183_48#_M1001_g N_VGND_c_728_n 0.00889942f $X=0.99 $Y=0.74 $X2=0
+ $Y2=0
cc_315 N_A_183_48#_M1003_g N_VGND_c_728_n 0.00820916f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_316 N_A_183_48#_M1005_g N_VGND_c_728_n 0.0075754f $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A_183_48#_M1009_g N_VGND_c_728_n 0.0075754f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A_183_48#_M1011_g N_VGND_c_728_n 0.00820718f $X=2.87 $Y=0.74 $X2=0
+ $Y2=0
cc_319 N_A_183_48#_M1015_g N_VGND_c_728_n 0.00820718f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A_183_48#_M1017_g N_VGND_c_728_n 0.00758198f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_321 N_A_183_48#_M1020_g N_VGND_c_728_n 0.0082143f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_322 N_A_183_48#_c_146_n N_VGND_c_728_n 0.00743504f $X=5.02 $Y=0.515 $X2=0
+ $Y2=0
cc_323 N_A_183_48#_c_149_n N_VGND_c_728_n 0.0119984f $X=5.96 $Y=0.515 $X2=0
+ $Y2=0
cc_324 N_A_27_368#_c_388_n N_VPWR_M1013_d 0.00400043f $X=0.72 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_325 N_A_27_368#_c_368_n N_VPWR_M1013_d 0.00553081f $X=0.805 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_326 N_A_27_368#_c_457_p N_VPWR_M1013_d 0.00168207f $X=0.805 $Y=2.325
+ $X2=-0.19 $Y2=-0.245
cc_327 N_A_27_368#_c_422_n N_VPWR_M1002_s 0.00379409f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_328 N_A_27_368#_c_422_n N_VPWR_M1007_s 0.00379409f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_329 N_A_27_368#_c_422_n N_VPWR_M1016_s 0.00379409f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_330 N_A_27_368#_c_422_n N_VPWR_M1022_s 0.00366644f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_331 N_A_27_368#_c_433_n N_VPWR_M1022_s 0.00361524f $X=4.48 $Y=2.24 $X2=0
+ $Y2=0
cc_332 N_A_27_368#_c_376_n N_VPWR_M1022_s 0.00174574f $X=4.99 $Y=1.885 $X2=0
+ $Y2=0
cc_333 N_A_27_368#_c_377_n N_VPWR_M1022_s 8.13096e-19 $X=4.565 $Y=1.885 $X2=0
+ $Y2=0
cc_334 N_A_27_368#_c_369_n N_VPWR_M1018_s 0.00328409f $X=5.475 $Y=1.485 $X2=0
+ $Y2=0
cc_335 N_A_27_368#_c_374_n N_VPWR_c_515_n 0.0157994f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_336 N_A_27_368#_c_388_n N_VPWR_c_515_n 0.00671628f $X=0.72 $Y=2.325 $X2=0
+ $Y2=0
cc_337 N_A_27_368#_c_422_n N_VPWR_c_515_n 0.00102433f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_338 N_A_27_368#_c_457_p N_VPWR_c_515_n 0.0137497f $X=0.805 $Y=2.325 $X2=0
+ $Y2=0
cc_339 N_A_27_368#_c_422_n N_VPWR_c_516_n 0.0171814f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_340 N_A_27_368#_c_422_n N_VPWR_c_517_n 0.0171814f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_341 N_A_27_368#_c_422_n N_VPWR_c_518_n 0.0171814f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_342 N_A_27_368#_c_371_n N_VPWR_c_519_n 0.00393828f $X=4.785 $Y=1.765 $X2=0
+ $Y2=0
cc_343 N_A_27_368#_c_422_n N_VPWR_c_519_n 0.0142616f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_344 N_A_27_368#_c_376_n N_VPWR_c_519_n 0.00272979f $X=4.99 $Y=1.885 $X2=0
+ $Y2=0
cc_345 N_A_27_368#_c_372_n N_VPWR_c_520_n 0.0044704f $X=5.235 $Y=1.765 $X2=0
+ $Y2=0
cc_346 N_A_27_368#_c_373_n N_VPWR_c_520_n 0.0130894f $X=5.735 $Y=1.765 $X2=0
+ $Y2=0
cc_347 N_A_27_368#_c_374_n N_VPWR_c_523_n 0.0145938f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_348 N_A_27_368#_c_371_n N_VPWR_c_527_n 0.00445602f $X=4.785 $Y=1.765 $X2=0
+ $Y2=0
cc_349 N_A_27_368#_c_372_n N_VPWR_c_527_n 0.00445602f $X=5.235 $Y=1.765 $X2=0
+ $Y2=0
cc_350 N_A_27_368#_c_373_n N_VPWR_c_528_n 0.00413917f $X=5.735 $Y=1.765 $X2=0
+ $Y2=0
cc_351 N_A_27_368#_c_371_n N_VPWR_c_514_n 0.00857432f $X=4.785 $Y=1.765 $X2=0
+ $Y2=0
cc_352 N_A_27_368#_c_372_n N_VPWR_c_514_n 0.00857378f $X=5.235 $Y=1.765 $X2=0
+ $Y2=0
cc_353 N_A_27_368#_c_373_n N_VPWR_c_514_n 0.00821221f $X=5.735 $Y=1.765 $X2=0
+ $Y2=0
cc_354 N_A_27_368#_c_374_n N_VPWR_c_514_n 0.0120466f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_355 N_A_27_368#_c_422_n N_Y_M1000_d 0.00890962f $X=4.395 $Y=2.325 $X2=0 $Y2=0
cc_356 N_A_27_368#_c_422_n N_Y_M1006_d 0.00891381f $X=4.395 $Y=2.325 $X2=0 $Y2=0
cc_357 N_A_27_368#_c_422_n N_Y_M1010_d 0.00891381f $X=4.395 $Y=2.325 $X2=0 $Y2=0
cc_358 N_A_27_368#_c_422_n N_Y_M1019_d 0.0157948f $X=4.395 $Y=2.325 $X2=0 $Y2=0
cc_359 N_A_27_368#_c_422_n N_Y_c_622_n 0.157165f $X=4.395 $Y=2.325 $X2=0 $Y2=0
cc_360 N_A_27_368#_c_377_n N_Y_c_622_n 0.00889663f $X=4.565 $Y=1.885 $X2=0 $Y2=0
cc_361 N_A_27_368#_M1004_g N_Y_c_618_n 6.39165e-19 $X=4.8 $Y=0.74 $X2=0 $Y2=0
cc_362 N_A_27_368#_c_368_n N_Y_c_657_n 0.012847f $X=0.805 $Y=2.24 $X2=0 $Y2=0
cc_363 N_A_27_368#_c_422_n N_Y_c_657_n 0.0172495f $X=4.395 $Y=2.325 $X2=0 $Y2=0
cc_364 N_A_27_368#_c_366_n Y 0.00596854f $X=0.72 $Y=1.095 $X2=0 $Y2=0
cc_365 N_A_27_368#_c_366_n Y 0.00417827f $X=0.72 $Y=1.095 $X2=0 $Y2=0
cc_366 N_A_27_368#_c_368_n Y 0.0464398f $X=0.805 $Y=2.24 $X2=0 $Y2=0
cc_367 N_A_27_368#_c_366_n N_VGND_M1021_d 0.00286042f $X=0.72 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_368 N_A_27_368#_c_365_n N_VGND_c_715_n 0.0182902f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_369 N_A_27_368#_c_366_n N_VGND_c_715_n 0.02058f $X=0.72 $Y=1.095 $X2=0 $Y2=0
cc_370 N_A_27_368#_M1004_g N_VGND_c_719_n 0.00796521f $X=4.8 $Y=0.74 $X2=0 $Y2=0
cc_371 N_A_27_368#_M1008_g N_VGND_c_719_n 4.26797e-19 $X=5.245 $Y=0.74 $X2=0
+ $Y2=0
cc_372 N_A_27_368#_M1004_g N_VGND_c_720_n 4.26797e-19 $X=4.8 $Y=0.74 $X2=0 $Y2=0
cc_373 N_A_27_368#_M1008_g N_VGND_c_720_n 0.00796521f $X=5.245 $Y=0.74 $X2=0
+ $Y2=0
cc_374 N_A_27_368#_M1012_g N_VGND_c_720_n 0.00503266f $X=5.745 $Y=0.74 $X2=0
+ $Y2=0
cc_375 N_A_27_368#_c_365_n N_VGND_c_721_n 0.011066f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_376 N_A_27_368#_M1004_g N_VGND_c_726_n 0.00383152f $X=4.8 $Y=0.74 $X2=0 $Y2=0
cc_377 N_A_27_368#_M1008_g N_VGND_c_726_n 0.00383152f $X=5.245 $Y=0.74 $X2=0
+ $Y2=0
cc_378 N_A_27_368#_M1012_g N_VGND_c_727_n 0.00434272f $X=5.745 $Y=0.74 $X2=0
+ $Y2=0
cc_379 N_A_27_368#_M1004_g N_VGND_c_728_n 0.00757689f $X=4.8 $Y=0.74 $X2=0 $Y2=0
cc_380 N_A_27_368#_M1008_g N_VGND_c_728_n 0.00757689f $X=5.245 $Y=0.74 $X2=0
+ $Y2=0
cc_381 N_A_27_368#_M1012_g N_VGND_c_728_n 0.00824376f $X=5.745 $Y=0.74 $X2=0
+ $Y2=0
cc_382 N_A_27_368#_c_365_n N_VGND_c_728_n 0.00915947f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_383 N_VPWR_M1002_s N_Y_c_622_n 0.00201049f $X=1.53 $Y=1.84 $X2=0 $Y2=0
cc_384 N_VPWR_M1007_s N_Y_c_622_n 0.00201049f $X=2.43 $Y=1.84 $X2=0 $Y2=0
cc_385 N_VPWR_M1016_s N_Y_c_622_n 0.00201049f $X=3.33 $Y=1.84 $X2=0 $Y2=0
cc_386 N_Y_c_613_n N_VGND_M1003_s 0.00253871f $X=2.06 $Y=1.005 $X2=0 $Y2=0
cc_387 N_Y_c_615_n N_VGND_M1009_s 0.00253871f $X=2.92 $Y=1.005 $X2=0 $Y2=0
cc_388 N_Y_c_617_n N_VGND_M1015_s 0.00250873f $X=3.92 $Y=1.045 $X2=0 $Y2=0
cc_389 Y N_VGND_c_715_n 0.0191764f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_390 N_Y_c_613_n N_VGND_c_716_n 0.0215485f $X=2.06 $Y=1.005 $X2=0 $Y2=0
cc_391 N_Y_c_614_n N_VGND_c_716_n 0.0142351f $X=2.155 $Y=0.515 $X2=0 $Y2=0
cc_392 Y N_VGND_c_716_n 0.0142986f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_393 N_Y_c_614_n N_VGND_c_717_n 0.0142351f $X=2.155 $Y=0.515 $X2=0 $Y2=0
cc_394 N_Y_c_615_n N_VGND_c_717_n 0.0215485f $X=2.92 $Y=1.005 $X2=0 $Y2=0
cc_395 N_Y_c_616_n N_VGND_c_717_n 0.0142986f $X=3.085 $Y=0.515 $X2=0 $Y2=0
cc_396 N_Y_c_616_n N_VGND_c_718_n 0.0173003f $X=3.085 $Y=0.515 $X2=0 $Y2=0
cc_397 N_Y_c_617_n N_VGND_c_718_n 0.0209867f $X=3.92 $Y=1.045 $X2=0 $Y2=0
cc_398 N_Y_c_618_n N_VGND_c_718_n 0.0173003f $X=4.085 $Y=0.515 $X2=0 $Y2=0
cc_399 N_Y_c_618_n N_VGND_c_719_n 0.0142986f $X=4.085 $Y=0.515 $X2=0 $Y2=0
cc_400 Y N_VGND_c_722_n 0.014552f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_401 N_Y_c_614_n N_VGND_c_723_n 0.00838873f $X=2.155 $Y=0.515 $X2=0 $Y2=0
cc_402 N_Y_c_616_n N_VGND_c_724_n 0.0144922f $X=3.085 $Y=0.515 $X2=0 $Y2=0
cc_403 N_Y_c_618_n N_VGND_c_725_n 0.0145639f $X=4.085 $Y=0.515 $X2=0 $Y2=0
cc_404 N_Y_c_614_n N_VGND_c_728_n 0.00694347f $X=2.155 $Y=0.515 $X2=0 $Y2=0
cc_405 N_Y_c_616_n N_VGND_c_728_n 0.0118826f $X=3.085 $Y=0.515 $X2=0 $Y2=0
cc_406 N_Y_c_618_n N_VGND_c_728_n 0.0119984f $X=4.085 $Y=0.515 $X2=0 $Y2=0
cc_407 Y N_VGND_c_728_n 0.0119791f $X=1.115 $Y=0.47 $X2=0 $Y2=0
