* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__nor3_4 A B C VGND VNB VPB VPWR Y
M1000 VPWR A a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=1.652e+12p ps=1.415e+07u
M1001 Y C VGND VNB nshort w=740000u l=150000u
+  ad=6.29e+11p pd=6.14e+06u as=1.22935e+12p ps=9.25e+06u
M1002 VGND A Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND C Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y C a_295_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=1.0458e+12p pd=6.56e+06u as=1.9762e+12p ps=1.303e+07u
M1007 a_295_368# C Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_368# B a_295_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_295_368# C Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_295_368# B a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_368# B a_295_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_295_368# B a_27_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y C a_295_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
