* File: sky130_fd_sc_ls__or2b_2.spice
* Created: Fri Aug 28 13:57:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__or2b_2.pex.spice"
.subckt sky130_fd_sc_ls__or2b_2  VNB VPB B_N A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_B_N_M1001_g N_A_27_368#_M1001_s VNB NSHORT L=0.15 W=0.55
+ AD=0.107506 AS=0.15675 PD=0.937984 PS=1.67 NRD=17.448 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1003 N_X_M1003_d N_A_187_48#_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.74
+ AD=0.10545 AS=0.144644 PD=1.025 PS=1.26202 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1004 N_X_M1003_d N_A_187_48#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.10545 AS=0.251922 PD=1.025 PS=1.53899 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75001 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1002 N_A_187_48#_M1002_d N_A_M1002_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1104 AS=0.217878 PD=0.985 PS=1.33101 NRD=12.18 NRS=0.936 M=1 R=4.26667
+ SA=75001.8 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1005_d N_A_27_368#_M1005_g N_A_187_48#_M1002_d VNB NSHORT L=0.15
+ W=0.64 AD=0.2336 AS=0.1104 PD=2.01 PS=0.985 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.3 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1006_d N_B_N_M1006_g N_A_27_368#_M1006_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.174 AS=0.2478 PD=1.29 PS=2.27 NRD=35.6767 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75002.5 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1006_d N_A_187_48#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.232 AS=0.2884 PD=1.72 PS=1.635 NRD=1.7533 NRS=20.2122 M=1 R=7.46667
+ SA=75000.6 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1008_d N_A_187_48#_M1008_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.240589 AS=0.2884 PD=1.62717 PS=1.635 NRD=1.7533 NRS=21.0987 M=1 R=7.46667
+ SA=75001.3 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1009 A_470_368# N_A_M1009_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.214811 PD=1.27 PS=1.45283 NRD=15.7403 NRS=26.5753 M=1 R=6.66667
+ SA=75001.9 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1007 N_A_187_48#_M1007_d N_A_27_368#_M1007_g A_470_368# VPB PHIGHVT L=0.15 W=1
+ AD=0.415 AS=0.135 PD=2.83 PS=1.27 NRD=25.5903 NRS=15.7403 M=1 R=6.66667
+ SA=75002.3 SB=75000.3 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ls__or2b_2.pxi.spice"
*
.ends
*
*
