# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__dfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__dfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.700000 2.025000 2.080000 2.355000 ;
        RECT 1.910000 1.125000 2.270000 1.780000 ;
        RECT 1.910000 1.780000 2.080000 2.025000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.530100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.640000 0.350000 8.070000 1.130000 ;
        RECT 7.665000 2.030000 8.070000 2.980000 ;
        RECT 7.900000 1.130000 8.070000 2.030000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.535700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.140000 0.350000 9.515000 1.130000 ;
        RECT 9.160000 1.820000 9.515000 2.980000 ;
        RECT 9.345000 1.130000 9.515000 1.820000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.500000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.600000 0.085000 ;
        RECT 0.625000  0.085000 1.005000 0.560000 ;
        RECT 1.855000  0.085000 2.205000 0.560000 ;
        RECT 3.980000  0.085000 4.310000 0.410000 ;
        RECT 6.080000  0.085000 6.410000 1.040000 ;
        RECT 7.140000  0.085000 7.470000 0.680000 ;
        RECT 8.710000  0.085000 8.960000 1.130000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 9.600000 3.415000 ;
        RECT 0.560000 2.060000 0.810000 3.245000 ;
        RECT 1.555000 2.885000 1.885000 3.245000 ;
        RECT 3.740000 2.925000 4.130000 3.245000 ;
        RECT 6.165000 2.390000 6.495000 3.245000 ;
        RECT 7.240000 2.030000 7.490000 3.245000 ;
        RECT 8.655000 1.820000 8.985000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.110000 1.720000 0.840000 1.890000 ;
      RECT 0.110000 1.890000 0.360000 2.980000 ;
      RECT 0.115000 0.350000 0.445000 0.730000 ;
      RECT 0.115000 0.730000 2.545000 0.900000 ;
      RECT 0.115000 0.900000 0.445000 1.010000 ;
      RECT 0.670000 0.900000 1.090000 1.550000 ;
      RECT 0.670000 1.550000 0.840000 1.720000 ;
      RECT 1.010000 1.815000 1.435000 2.545000 ;
      RECT 1.010000 2.545000 2.225000 2.715000 ;
      RECT 1.010000 2.715000 1.340000 2.980000 ;
      RECT 1.265000 1.070000 1.595000 1.485000 ;
      RECT 1.265000 1.485000 1.740000 1.815000 ;
      RECT 2.055000 2.715000 4.470000 2.755000 ;
      RECT 2.055000 2.755000 3.290000 2.885000 ;
      RECT 2.250000 2.045000 2.610000 2.375000 ;
      RECT 2.375000 0.255000 3.655000 0.425000 ;
      RECT 2.375000 0.425000 2.545000 0.730000 ;
      RECT 2.440000 1.070000 2.885000 1.240000 ;
      RECT 2.440000 1.240000 2.610000 2.045000 ;
      RECT 2.715000 0.595000 2.885000 1.070000 ;
      RECT 2.780000 1.410000 3.315000 1.580000 ;
      RECT 2.780000 1.580000 2.950000 2.245000 ;
      RECT 2.780000 2.245000 4.280000 2.415000 ;
      RECT 2.780000 2.415000 2.950000 2.545000 ;
      RECT 3.065000 0.595000 3.315000 1.410000 ;
      RECT 3.120000 1.750000 3.655000 2.075000 ;
      RECT 3.120000 2.585000 4.470000 2.715000 ;
      RECT 3.485000 0.425000 3.655000 0.580000 ;
      RECT 3.485000 0.580000 5.715000 0.620000 ;
      RECT 3.485000 0.620000 4.650000 0.750000 ;
      RECT 3.485000 0.750000 3.655000 1.750000 ;
      RECT 3.825000 1.015000 4.900000 1.185000 ;
      RECT 3.825000 1.185000 4.620000 1.370000 ;
      RECT 4.020000 1.630000 4.280000 2.245000 ;
      RECT 4.300000 2.755000 4.470000 2.800000 ;
      RECT 4.300000 2.800000 5.150000 2.905000 ;
      RECT 4.300000 2.905000 5.990000 3.075000 ;
      RECT 4.450000 1.370000 4.620000 1.855000 ;
      RECT 4.450000 1.855000 4.810000 2.025000 ;
      RECT 4.480000 0.290000 5.715000 0.580000 ;
      RECT 4.570000 0.920000 4.900000 1.015000 ;
      RECT 4.640000 2.025000 4.810000 2.615000 ;
      RECT 4.790000 1.355000 5.150000 1.685000 ;
      RECT 4.980000 1.685000 5.150000 2.800000 ;
      RECT 5.125000 0.790000 5.590000 1.120000 ;
      RECT 5.320000 1.120000 5.590000 1.210000 ;
      RECT 5.320000 1.210000 7.130000 1.380000 ;
      RECT 5.320000 1.380000 5.490000 2.115000 ;
      RECT 5.320000 2.115000 5.570000 2.735000 ;
      RECT 5.660000 1.615000 5.990000 1.945000 ;
      RECT 5.820000 1.945000 5.990000 2.905000 ;
      RECT 6.230000 1.550000 6.560000 1.690000 ;
      RECT 6.230000 1.690000 7.730000 1.860000 ;
      RECT 6.230000 1.860000 7.040000 2.220000 ;
      RECT 6.640000 0.440000 6.970000 0.850000 ;
      RECT 6.640000 0.850000 7.470000 1.020000 ;
      RECT 6.710000 2.220000 7.040000 2.860000 ;
      RECT 6.800000 1.190000 7.130000 1.210000 ;
      RECT 6.800000 1.380000 7.130000 1.520000 ;
      RECT 7.300000 1.020000 7.470000 1.350000 ;
      RECT 7.300000 1.350000 7.730000 1.690000 ;
      RECT 8.280000 0.625000 8.530000 1.300000 ;
      RECT 8.280000 1.300000 9.175000 1.630000 ;
      RECT 8.280000 1.630000 8.455000 2.700000 ;
  END
END sky130_fd_sc_ls__dfxbp_1
