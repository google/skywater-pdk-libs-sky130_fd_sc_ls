* File: sky130_fd_sc_ls__o311ai_4.pxi.spice
* Created: Wed Sep  2 11:21:50 2020
* 
x_PM_SKY130_FD_SC_LS__O311AI_4%C1 N_C1_c_146_n N_C1_M1003_g N_C1_c_153_n
+ N_C1_M1011_g N_C1_c_147_n N_C1_M1018_g N_C1_c_154_n N_C1_M1022_g N_C1_c_148_n
+ N_C1_M1019_g N_C1_c_149_n N_C1_c_150_n N_C1_c_151_n N_C1_M1029_g C1 C1
+ N_C1_c_152_n PM_SKY130_FD_SC_LS__O311AI_4%C1
x_PM_SKY130_FD_SC_LS__O311AI_4%B1 N_B1_c_220_n N_B1_M1020_g N_B1_c_212_n
+ N_B1_c_213_n N_B1_c_223_n N_B1_M1028_g N_B1_M1002_g N_B1_M1014_g N_B1_M1015_g
+ N_B1_M1027_g B1 B1 B1 B1 N_B1_c_219_n PM_SKY130_FD_SC_LS__O311AI_4%B1
x_PM_SKY130_FD_SC_LS__O311AI_4%A3 N_A3_c_284_n N_A3_M1000_g N_A3_M1008_g
+ N_A3_c_285_n N_A3_M1009_g N_A3_M1010_g N_A3_c_286_n N_A3_M1030_g N_A3_M1024_g
+ N_A3_c_287_n N_A3_M1032_g N_A3_M1031_g A3 A3 N_A3_c_288_n N_A3_c_282_n
+ N_A3_c_290_n N_A3_c_283_n A3 PM_SKY130_FD_SC_LS__O311AI_4%A3
x_PM_SKY130_FD_SC_LS__O311AI_4%A2 N_A2_c_381_n N_A2_M1006_g N_A2_M1001_g
+ N_A2_c_382_n N_A2_M1021_g N_A2_M1004_g N_A2_c_383_n N_A2_M1026_g N_A2_c_378_n
+ N_A2_M1016_g N_A2_c_384_n N_A2_M1033_g N_A2_c_379_n N_A2_M1025_g A2 A2
+ N_A2_c_385_n N_A2_c_380_n PM_SKY130_FD_SC_LS__O311AI_4%A2
x_PM_SKY130_FD_SC_LS__O311AI_4%A1 N_A1_M1005_g N_A1_c_466_n N_A1_c_467_n
+ N_A1_M1012_g N_A1_c_474_n N_A1_M1007_g N_A1_c_475_n N_A1_M1013_g N_A1_c_476_n
+ N_A1_M1017_g N_A1_c_469_n N_A1_M1034_g N_A1_c_477_n N_A1_M1023_g N_A1_c_470_n
+ N_A1_M1035_g A1 A1 A1 N_A1_c_478_n N_A1_c_471_n
+ PM_SKY130_FD_SC_LS__O311AI_4%A1
x_PM_SKY130_FD_SC_LS__O311AI_4%VPWR N_VPWR_M1011_d N_VPWR_M1022_d N_VPWR_M1028_s
+ N_VPWR_M1007_d N_VPWR_M1013_d N_VPWR_M1023_d N_VPWR_c_547_n N_VPWR_c_548_n
+ N_VPWR_c_549_n N_VPWR_c_550_n N_VPWR_c_551_n N_VPWR_c_552_n N_VPWR_c_553_n
+ N_VPWR_c_554_n N_VPWR_c_555_n VPWR N_VPWR_c_556_n N_VPWR_c_557_n
+ N_VPWR_c_558_n N_VPWR_c_559_n N_VPWR_c_560_n N_VPWR_c_561_n N_VPWR_c_562_n
+ N_VPWR_c_546_n PM_SKY130_FD_SC_LS__O311AI_4%VPWR
x_PM_SKY130_FD_SC_LS__O311AI_4%Y N_Y_M1003_d N_Y_M1019_d N_Y_M1011_s N_Y_M1020_d
+ N_Y_M1000_s N_Y_M1030_s N_Y_c_668_n N_Y_c_662_n N_Y_c_673_n N_Y_c_659_n
+ N_Y_c_663_n N_Y_c_664_n N_Y_c_719_n N_Y_c_721_n N_Y_c_726_n N_Y_c_680_n
+ N_Y_c_685_n N_Y_c_665_n N_Y_c_666_n N_Y_c_734_n Y Y N_Y_c_660_n Y
+ PM_SKY130_FD_SC_LS__O311AI_4%Y
x_PM_SKY130_FD_SC_LS__O311AI_4%A_841_368# N_A_841_368#_M1000_d
+ N_A_841_368#_M1009_d N_A_841_368#_M1032_d N_A_841_368#_M1021_d
+ N_A_841_368#_M1033_d N_A_841_368#_c_796_n N_A_841_368#_c_797_n
+ N_A_841_368#_c_798_n N_A_841_368#_c_854_n N_A_841_368#_c_799_n
+ N_A_841_368#_c_813_n N_A_841_368#_c_800_n N_A_841_368#_c_862_p
+ N_A_841_368#_c_801_n N_A_841_368#_c_802_n N_A_841_368#_c_803_n
+ N_A_841_368#_c_804_n N_A_841_368#_c_805_n
+ PM_SKY130_FD_SC_LS__O311AI_4%A_841_368#
x_PM_SKY130_FD_SC_LS__O311AI_4%A_1350_368# N_A_1350_368#_M1006_s
+ N_A_1350_368#_M1026_s N_A_1350_368#_M1007_s N_A_1350_368#_M1017_s
+ N_A_1350_368#_c_870_n N_A_1350_368#_c_874_n N_A_1350_368#_c_867_n
+ N_A_1350_368#_c_868_n N_A_1350_368#_c_888_n N_A_1350_368#_c_892_n
+ N_A_1350_368#_c_869_n N_A_1350_368#_c_877_n N_A_1350_368#_c_881_n
+ N_A_1350_368#_c_897_n PM_SKY130_FD_SC_LS__O311AI_4%A_1350_368#
x_PM_SKY130_FD_SC_LS__O311AI_4%A_27_74# N_A_27_74#_M1003_s N_A_27_74#_M1018_s
+ N_A_27_74#_M1029_s N_A_27_74#_M1014_s N_A_27_74#_M1027_s N_A_27_74#_c_923_n
+ N_A_27_74#_c_924_n N_A_27_74#_c_925_n N_A_27_74#_c_948_n N_A_27_74#_c_926_n
+ PM_SKY130_FD_SC_LS__O311AI_4%A_27_74#
x_PM_SKY130_FD_SC_LS__O311AI_4%A_459_74# N_A_459_74#_M1002_d N_A_459_74#_M1015_d
+ N_A_459_74#_M1008_s N_A_459_74#_M1024_s N_A_459_74#_M1001_s
+ N_A_459_74#_M1016_s N_A_459_74#_M1005_s N_A_459_74#_M1034_s
+ N_A_459_74#_c_963_n N_A_459_74#_c_964_n N_A_459_74#_c_965_n
+ N_A_459_74#_c_966_n N_A_459_74#_c_967_n N_A_459_74#_c_991_n
+ N_A_459_74#_c_968_n N_A_459_74#_c_996_n N_A_459_74#_c_969_n
+ N_A_459_74#_c_970_n N_A_459_74#_c_971_n N_A_459_74#_c_972_n
+ N_A_459_74#_c_973_n N_A_459_74#_c_974_n N_A_459_74#_c_975_n
+ N_A_459_74#_c_976_n N_A_459_74#_c_998_n N_A_459_74#_c_999_n
+ N_A_459_74#_c_977_n N_A_459_74#_c_978_n N_A_459_74#_c_1039_n
+ PM_SKY130_FD_SC_LS__O311AI_4%A_459_74#
x_PM_SKY130_FD_SC_LS__O311AI_4%VGND N_VGND_M1008_d N_VGND_M1010_d N_VGND_M1031_d
+ N_VGND_M1004_d N_VGND_M1025_d N_VGND_M1012_d N_VGND_M1035_d N_VGND_c_1112_n
+ N_VGND_c_1113_n N_VGND_c_1114_n N_VGND_c_1115_n N_VGND_c_1116_n
+ N_VGND_c_1117_n N_VGND_c_1118_n VGND N_VGND_c_1119_n N_VGND_c_1120_n
+ N_VGND_c_1121_n N_VGND_c_1122_n N_VGND_c_1123_n N_VGND_c_1124_n
+ N_VGND_c_1125_n N_VGND_c_1126_n N_VGND_c_1127_n N_VGND_c_1128_n
+ N_VGND_c_1129_n N_VGND_c_1130_n N_VGND_c_1131_n N_VGND_c_1132_n
+ PM_SKY130_FD_SC_LS__O311AI_4%VGND
cc_1 VNB N_C1_c_146_n 0.0204707f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_2 VNB N_C1_c_147_n 0.0152712f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.185
cc_3 VNB N_C1_c_148_n 0.0149102f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.185
cc_4 VNB N_C1_c_149_n 0.0223569f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=1.26
cc_5 VNB N_C1_c_150_n 0.121207f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=1.26
cc_6 VNB N_C1_c_151_n 0.0147616f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.185
cc_7 VNB N_C1_c_152_n 0.0156012f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.465
cc_8 VNB N_B1_c_212_n 0.00834596f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_9 VNB N_B1_c_213_n 0.00672099f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_10 VNB N_B1_M1002_g 0.023123f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=2.4
cc_11 VNB N_B1_M1014_g 0.0221713f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=0.74
cc_12 VNB N_B1_M1015_g 0.0223226f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=0.74
cc_13 VNB N_B1_M1027_g 0.0304926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB B1 0.0110294f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.475
cc_15 VNB N_B1_c_219_n 0.0823936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A3_M1008_g 0.0287422f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_17 VNB N_A3_M1010_g 0.0244469f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.185
cc_18 VNB N_A3_M1024_g 0.0244287f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=0.74
cc_19 VNB N_A3_M1031_g 0.0247143f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.465
cc_20 VNB N_A3_c_282_n 0.0939197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A3_c_283_n 0.0023959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_M1001_g 0.0258894f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_23 VNB N_A2_M1004_g 0.0230723f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.185
cc_24 VNB N_A2_c_378_n 0.016486f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.185
cc_25 VNB N_A2_c_379_n 0.0161012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_c_380_n 0.106649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A1_M1005_g 0.0315883f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_28 VNB N_A1_c_466_n 0.00596486f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_29 VNB N_A1_c_467_n 0.00495433f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_30 VNB N_A1_M1012_g 0.0316257f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.74
cc_31 VNB N_A1_c_469_n 0.0189372f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=0.74
cc_32 VNB N_A1_c_470_n 0.0198259f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.465
cc_33 VNB N_A1_c_471_n 0.11825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_546_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_659_n 0.0471346f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.475
cc_36 VNB N_Y_c_660_n 0.00164207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB Y 0.00406123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_74#_c_923_n 0.012589f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=1.26
cc_39 VNB N_A_27_74#_c_924_n 0.0218403f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.185
cc_40 VNB N_A_27_74#_c_925_n 0.00963967f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=0.74
cc_41 VNB N_A_27_74#_c_926_n 0.00205354f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.465
cc_42 VNB N_A_459_74#_c_963_n 0.0207409f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.475
cc_43 VNB N_A_459_74#_c_964_n 0.00525772f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.465
cc_44 VNB N_A_459_74#_c_965_n 0.00638704f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.465
cc_45 VNB N_A_459_74#_c_966_n 0.00387414f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=1.475
cc_46 VNB N_A_459_74#_c_967_n 0.00206045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_459_74#_c_968_n 0.00239415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_459_74#_c_969_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_459_74#_c_970_n 0.00672511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_459_74#_c_971_n 0.00181921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_459_74#_c_972_n 0.012969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_459_74#_c_973_n 0.00206647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_459_74#_c_974_n 0.00159982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_459_74#_c_975_n 0.0106354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_459_74#_c_976_n 0.00220643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_459_74#_c_977_n 0.00190558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_459_74#_c_978_n 0.0010144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1112_n 0.0105224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1113_n 0.00794664f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.475
cc_60 VNB N_VGND_c_1114_n 0.00801909f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.465
cc_61 VNB N_VGND_c_1115_n 0.00512538f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_62 VNB N_VGND_c_1116_n 0.00647008f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.54
cc_63 VNB N_VGND_c_1117_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.54
cc_64 VNB N_VGND_c_1118_n 0.0505272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1119_n 0.109865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1120_n 0.0159624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1121_n 0.0180412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1122_n 0.0166074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1123_n 0.0189911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1124_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1125_n 0.00613127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1126_n 0.00632082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1127_n 0.00651315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1128_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1129_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1130_n 0.0172515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1131_n 0.0262931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1132_n 0.564514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VPB N_C1_c_153_n 0.0203833f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_80 VPB N_C1_c_154_n 0.0171086f $X=-0.19 $Y=1.66 $X2=1.18 $Y2=1.765
cc_81 VPB N_C1_c_150_n 0.0151029f $X=-0.19 $Y=1.66 $X2=1.435 $Y2=1.26
cc_82 VPB N_C1_c_152_n 0.0173437f $X=-0.19 $Y=1.66 $X2=1.075 $Y2=1.465
cc_83 VPB N_B1_c_220_n 0.0161908f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.185
cc_84 VPB N_B1_c_212_n 0.00761466f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_85 VPB N_B1_c_213_n 0.00557822f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_86 VPB N_B1_c_223_n 0.0178223f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_87 VPB B1 0.0220575f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.475
cc_88 VPB N_B1_c_219_n 0.0548315f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A3_c_284_n 0.0188518f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.185
cc_90 VPB N_A3_c_285_n 0.0155751f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=0.74
cc_91 VPB N_A3_c_286_n 0.0163916f $X=-0.19 $Y=1.66 $X2=1.36 $Y2=0.74
cc_92 VPB N_A3_c_287_n 0.0160381f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_93 VPB N_A3_c_288_n 0.00445883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A3_c_282_n 0.0591735f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A3_c_290_n 0.00416634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A2_c_381_n 0.0152626f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.185
cc_97 VPB N_A2_c_382_n 0.0157714f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=0.74
cc_98 VPB N_A2_c_383_n 0.0154462f $X=-0.19 $Y=1.66 $X2=1.36 $Y2=0.74
cc_99 VPB N_A2_c_384_n 0.0187612f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_100 VPB N_A2_c_385_n 0.00752098f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.54
cc_101 VPB N_A2_c_380_n 0.0476822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A1_c_466_n 0.00794688f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_103 VPB N_A1_c_467_n 0.00495506f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_104 VPB N_A1_c_474_n 0.0190573f $X=-0.19 $Y=1.66 $X2=1.18 $Y2=2.4
cc_105 VPB N_A1_c_475_n 0.0149966f $X=-0.19 $Y=1.66 $X2=1.36 $Y2=0.74
cc_106 VPB N_A1_c_476_n 0.0149989f $X=-0.19 $Y=1.66 $X2=1.435 $Y2=1.26
cc_107 VPB N_A1_c_477_n 0.0177521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A1_c_478_n 0.00921801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A1_c_471_n 0.0547331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_547_n 0.0120106f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=0.74
cc_111 VPB N_VPWR_c_548_n 0.0489067f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_112 VPB N_VPWR_c_549_n 0.00581763f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.465
cc_113 VPB N_VPWR_c_550_n 0.0115963f $X=-0.19 $Y=1.66 $X2=1.075 $Y2=1.475
cc_114 VPB N_VPWR_c_551_n 0.00271781f $X=-0.19 $Y=1.66 $X2=1.36 $Y2=1.185
cc_115 VPB N_VPWR_c_552_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_553_n 0.0639451f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.54
cc_117 VPB N_VPWR_c_554_n 0.0223565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_555_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_556_n 0.113171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_557_n 0.0159778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_558_n 0.0182909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_559_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_560_n 0.0614903f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_561_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_562_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_546_n 0.116297f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_Y_c_662_n 0.00330637f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.475
cc_128 VPB N_Y_c_663_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.075 $Y2=1.465
cc_129 VPB N_Y_c_664_n 0.0148222f $X=-0.19 $Y=1.66 $X2=1.36 $Y2=1.185
cc_130 VPB N_Y_c_665_n 0.00237222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_Y_c_666_n 0.00212753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB Y 0.00203304f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_841_368#_c_796_n 0.00748204f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=1.185
cc_134 VPB N_A_841_368#_c_797_n 0.00273412f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=0.74
cc_135 VPB N_A_841_368#_c_798_n 0.00483682f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_136 VPB N_A_841_368#_c_799_n 0.00392363f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.465
cc_137 VPB N_A_841_368#_c_800_n 0.00273412f $X=-0.19 $Y=1.66 $X2=1.075 $Y2=1.465
cc_138 VPB N_A_841_368#_c_801_n 0.00669267f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_841_368#_c_802_n 0.00528239f $X=-0.19 $Y=1.66 $X2=1.075 $Y2=1.54
cc_140 VPB N_A_841_368#_c_803_n 0.00244483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_841_368#_c_804_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_841_368#_c_805_n 0.00257243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_1350_368#_c_867_n 0.0132311f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_144 VPB N_A_1350_368#_c_868_n 0.00233217f $X=-0.19 $Y=1.66 $X2=0.395
+ $Y2=1.475
cc_145 VPB N_A_1350_368#_c_869_n 0.00243101f $X=-0.19 $Y=1.66 $X2=1.075
+ $Y2=1.475
cc_146 N_C1_c_154_n N_B1_c_220_n 0.0297694f $X=1.18 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_147 N_C1_c_149_n N_B1_c_213_n 0.0162438f $X=1.715 $Y=1.26 $X2=0 $Y2=0
cc_148 N_C1_c_150_n N_B1_c_213_n 0.00848653f $X=1.435 $Y=1.26 $X2=0 $Y2=0
cc_149 N_C1_c_152_n N_B1_c_213_n 0.00125707f $X=1.075 $Y=1.465 $X2=0 $Y2=0
cc_150 N_C1_c_151_n N_B1_M1002_g 0.0324285f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_151 N_C1_c_153_n N_VPWR_c_548_n 0.01858f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_152 N_C1_c_154_n N_VPWR_c_548_n 8.11309e-19 $X=1.18 $Y=1.765 $X2=0 $Y2=0
cc_153 N_C1_c_150_n N_VPWR_c_548_n 9.23094e-19 $X=1.435 $Y=1.26 $X2=0 $Y2=0
cc_154 N_C1_c_152_n N_VPWR_c_548_n 0.0257495f $X=1.075 $Y=1.465 $X2=0 $Y2=0
cc_155 N_C1_c_153_n N_VPWR_c_549_n 5.77739e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_156 N_C1_c_154_n N_VPWR_c_549_n 0.0111057f $X=1.18 $Y=1.765 $X2=0 $Y2=0
cc_157 N_C1_c_153_n N_VPWR_c_554_n 0.00413917f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_158 N_C1_c_154_n N_VPWR_c_554_n 0.00413917f $X=1.18 $Y=1.765 $X2=0 $Y2=0
cc_159 N_C1_c_153_n N_VPWR_c_546_n 0.00819493f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_160 N_C1_c_154_n N_VPWR_c_546_n 0.00819493f $X=1.18 $Y=1.765 $X2=0 $Y2=0
cc_161 N_C1_c_153_n N_Y_c_668_n 0.0018637f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_162 N_C1_c_150_n N_Y_c_668_n 0.00175566f $X=1.435 $Y=1.26 $X2=0 $Y2=0
cc_163 N_C1_c_152_n N_Y_c_668_n 0.0284242f $X=1.075 $Y=1.465 $X2=0 $Y2=0
cc_164 N_C1_c_153_n N_Y_c_662_n 0.00869413f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_165 N_C1_c_154_n N_Y_c_662_n 0.00643865f $X=1.18 $Y=1.765 $X2=0 $Y2=0
cc_166 N_C1_c_154_n N_Y_c_673_n 0.0160448f $X=1.18 $Y=1.765 $X2=0 $Y2=0
cc_167 N_C1_c_149_n N_Y_c_673_n 4.9691e-19 $X=1.715 $Y=1.26 $X2=0 $Y2=0
cc_168 N_C1_c_150_n N_Y_c_673_n 0.00716273f $X=1.435 $Y=1.26 $X2=0 $Y2=0
cc_169 N_C1_c_152_n N_Y_c_673_n 0.0114816f $X=1.075 $Y=1.465 $X2=0 $Y2=0
cc_170 N_C1_c_149_n N_Y_c_659_n 0.00350562f $X=1.715 $Y=1.26 $X2=0 $Y2=0
cc_171 N_C1_c_151_n N_Y_c_659_n 0.00520798f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_172 N_C1_c_154_n N_Y_c_663_n 6.21762e-19 $X=1.18 $Y=1.765 $X2=0 $Y2=0
cc_173 N_C1_c_146_n N_Y_c_680_n 0.00429752f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_174 N_C1_c_147_n N_Y_c_680_n 0.0128945f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_175 N_C1_c_148_n N_Y_c_680_n 0.0147571f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_176 N_C1_c_150_n N_Y_c_680_n 0.00585463f $X=1.435 $Y=1.26 $X2=0 $Y2=0
cc_177 N_C1_c_152_n N_Y_c_680_n 0.0419281f $X=1.075 $Y=1.465 $X2=0 $Y2=0
cc_178 N_C1_c_147_n N_Y_c_685_n 4.05917e-19 $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_179 N_C1_c_148_n N_Y_c_685_n 0.0036256f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_180 N_C1_c_149_n N_Y_c_685_n 0.0130927f $X=1.715 $Y=1.26 $X2=0 $Y2=0
cc_181 N_C1_c_150_n N_Y_c_685_n 0.00507672f $X=1.435 $Y=1.26 $X2=0 $Y2=0
cc_182 N_C1_c_151_n N_Y_c_685_n 0.00632997f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_183 N_C1_c_154_n N_Y_c_665_n 6.04745e-19 $X=1.18 $Y=1.765 $X2=0 $Y2=0
cc_184 N_C1_c_146_n N_A_27_74#_c_924_n 0.00194058f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_185 N_C1_c_150_n N_A_27_74#_c_924_n 0.00381029f $X=1.435 $Y=1.26 $X2=0 $Y2=0
cc_186 N_C1_c_152_n N_A_27_74#_c_924_n 0.0211412f $X=1.075 $Y=1.465 $X2=0 $Y2=0
cc_187 N_C1_c_146_n N_A_27_74#_c_925_n 0.0144205f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_188 N_C1_c_147_n N_A_27_74#_c_925_n 0.0102631f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_189 N_C1_c_148_n N_A_27_74#_c_925_n 0.0101492f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_190 N_C1_c_149_n N_A_27_74#_c_925_n 3.14401e-19 $X=1.715 $Y=1.26 $X2=0 $Y2=0
cc_191 N_C1_c_151_n N_A_27_74#_c_925_n 0.0121821f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_192 N_C1_c_151_n N_A_459_74#_c_963_n 2.00992e-19 $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_193 N_C1_c_146_n N_VGND_c_1119_n 0.00291649f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_194 N_C1_c_147_n N_VGND_c_1119_n 0.00291649f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_195 N_C1_c_148_n N_VGND_c_1119_n 0.00291649f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_196 N_C1_c_151_n N_VGND_c_1119_n 0.00291649f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_197 N_C1_c_146_n N_VGND_c_1132_n 0.00362829f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_198 N_C1_c_147_n N_VGND_c_1132_n 0.00359171f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_199 N_C1_c_148_n N_VGND_c_1132_n 0.00359121f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_200 N_C1_c_151_n N_VGND_c_1132_n 0.00359219f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_201 B1 N_A3_c_284_n 4.83587e-19 $X=3.995 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_202 B1 N_A3_c_282_n 0.00640001f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_203 B1 N_A3_c_283_n 0.0124194f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_204 N_B1_c_220_n N_VPWR_c_549_n 0.00548019f $X=1.68 $Y=1.765 $X2=0 $Y2=0
cc_205 N_B1_c_220_n N_VPWR_c_559_n 0.00445602f $X=1.68 $Y=1.765 $X2=0 $Y2=0
cc_206 N_B1_c_223_n N_VPWR_c_559_n 0.00445602f $X=2.13 $Y=1.765 $X2=0 $Y2=0
cc_207 N_B1_c_223_n N_VPWR_c_560_n 0.00400188f $X=2.13 $Y=1.765 $X2=0 $Y2=0
cc_208 N_B1_c_220_n N_VPWR_c_546_n 0.00857432f $X=1.68 $Y=1.765 $X2=0 $Y2=0
cc_209 N_B1_c_223_n N_VPWR_c_546_n 0.00861697f $X=2.13 $Y=1.765 $X2=0 $Y2=0
cc_210 N_B1_c_220_n N_Y_c_673_n 0.0129388f $X=1.68 $Y=1.765 $X2=0 $Y2=0
cc_211 N_B1_c_212_n N_Y_c_659_n 0.00738449f $X=2.04 $Y=1.65 $X2=0 $Y2=0
cc_212 N_B1_M1002_g N_Y_c_659_n 0.0133957f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_213 N_B1_M1014_g N_Y_c_659_n 0.0104926f $X=2.65 $Y=0.74 $X2=0 $Y2=0
cc_214 N_B1_M1015_g N_Y_c_659_n 0.0105534f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_215 N_B1_M1027_g N_Y_c_659_n 0.0125939f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_216 B1 N_Y_c_659_n 0.147849f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_217 N_B1_c_219_n N_Y_c_659_n 0.00784304f $X=3.43 $Y=1.515 $X2=0 $Y2=0
cc_218 N_B1_c_220_n N_Y_c_663_n 0.0108556f $X=1.68 $Y=1.765 $X2=0 $Y2=0
cc_219 N_B1_c_223_n N_Y_c_663_n 0.0150947f $X=2.13 $Y=1.765 $X2=0 $Y2=0
cc_220 N_B1_c_223_n N_Y_c_664_n 0.0161429f $X=2.13 $Y=1.765 $X2=0 $Y2=0
cc_221 B1 N_Y_c_664_n 0.152506f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_222 N_B1_c_219_n N_Y_c_664_n 0.00808202f $X=3.43 $Y=1.515 $X2=0 $Y2=0
cc_223 N_B1_c_213_n N_Y_c_685_n 6.83304e-19 $X=1.77 $Y=1.65 $X2=0 $Y2=0
cc_224 N_B1_M1002_g N_Y_c_685_n 9.07448e-19 $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_225 N_B1_c_220_n N_Y_c_665_n 0.00316685f $X=1.68 $Y=1.765 $X2=0 $Y2=0
cc_226 N_B1_c_212_n N_Y_c_665_n 0.00760533f $X=2.04 $Y=1.65 $X2=0 $Y2=0
cc_227 N_B1_c_213_n N_Y_c_665_n 4.64856e-19 $X=1.77 $Y=1.65 $X2=0 $Y2=0
cc_228 N_B1_c_223_n N_Y_c_665_n 0.00631593f $X=2.13 $Y=1.765 $X2=0 $Y2=0
cc_229 N_B1_c_219_n N_Y_c_665_n 4.64856e-19 $X=3.43 $Y=1.515 $X2=0 $Y2=0
cc_230 N_B1_M1002_g N_A_27_74#_c_925_n 4.56461e-19 $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_231 N_B1_M1002_g N_A_27_74#_c_926_n 0.0106751f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_232 N_B1_M1014_g N_A_27_74#_c_926_n 0.00838518f $X=2.65 $Y=0.74 $X2=0 $Y2=0
cc_233 N_B1_M1015_g N_A_27_74#_c_926_n 0.00849254f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_234 N_B1_M1027_g N_A_27_74#_c_926_n 0.00849254f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_235 N_B1_M1002_g N_A_459_74#_c_963_n 0.00375385f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_236 N_B1_M1014_g N_A_459_74#_c_963_n 0.0103107f $X=2.65 $Y=0.74 $X2=0 $Y2=0
cc_237 N_B1_M1015_g N_A_459_74#_c_963_n 0.0103245f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_238 N_B1_M1027_g N_A_459_74#_c_963_n 0.0131979f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_239 N_B1_M1027_g N_A_459_74#_c_964_n 0.00284982f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_240 N_B1_M1002_g N_VGND_c_1119_n 0.00329872f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_241 N_B1_M1014_g N_VGND_c_1119_n 0.00288916f $X=2.65 $Y=0.74 $X2=0 $Y2=0
cc_242 N_B1_M1015_g N_VGND_c_1119_n 0.00288916f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_243 N_B1_M1027_g N_VGND_c_1119_n 0.00288916f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_244 N_B1_M1002_g N_VGND_c_1132_n 0.00428036f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_245 N_B1_M1014_g N_VGND_c_1132_n 0.0035719f $X=2.65 $Y=0.74 $X2=0 $Y2=0
cc_246 N_B1_M1015_g N_VGND_c_1132_n 0.0035729f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_247 N_B1_M1027_g N_VGND_c_1132_n 0.00362289f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A3_c_287_n N_A2_c_381_n 0.0229358f $X=6.225 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_249 N_A3_M1031_g N_A2_M1001_g 0.0234798f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A3_c_288_n N_A2_c_380_n 2.44878e-19 $X=6.03 $Y=1.515 $X2=0 $Y2=0
cc_251 N_A3_c_282_n N_A2_c_380_n 0.0192109f $X=6.225 $Y=1.557 $X2=0 $Y2=0
cc_252 N_A3_c_284_n N_VPWR_c_556_n 0.00278257f $X=4.575 $Y=1.765 $X2=0 $Y2=0
cc_253 N_A3_c_285_n N_VPWR_c_556_n 0.00278271f $X=5.075 $Y=1.765 $X2=0 $Y2=0
cc_254 N_A3_c_286_n N_VPWR_c_556_n 0.00278271f $X=5.595 $Y=1.765 $X2=0 $Y2=0
cc_255 N_A3_c_287_n N_VPWR_c_556_n 0.00278257f $X=6.225 $Y=1.765 $X2=0 $Y2=0
cc_256 N_A3_c_284_n N_VPWR_c_560_n 0.00232643f $X=4.575 $Y=1.765 $X2=0 $Y2=0
cc_257 N_A3_c_284_n N_VPWR_c_546_n 0.00359084f $X=4.575 $Y=1.765 $X2=0 $Y2=0
cc_258 N_A3_c_285_n N_VPWR_c_546_n 0.00354917f $X=5.075 $Y=1.765 $X2=0 $Y2=0
cc_259 N_A3_c_286_n N_VPWR_c_546_n 0.00355928f $X=5.595 $Y=1.765 $X2=0 $Y2=0
cc_260 N_A3_c_287_n N_VPWR_c_546_n 0.00355377f $X=6.225 $Y=1.765 $X2=0 $Y2=0
cc_261 N_A3_M1008_g N_Y_c_659_n 0.0125331f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A3_M1010_g N_Y_c_659_n 0.011293f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A3_M1024_g N_Y_c_659_n 0.0112465f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A3_M1031_g N_Y_c_659_n 0.0143698f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A3_c_282_n N_Y_c_659_n 0.018496f $X=6.225 $Y=1.557 $X2=0 $Y2=0
cc_266 N_A3_c_283_n N_Y_c_659_n 0.125235f $X=5.185 $Y=1.605 $X2=0 $Y2=0
cc_267 N_A3_c_284_n N_Y_c_664_n 0.0177015f $X=4.575 $Y=1.765 $X2=0 $Y2=0
cc_268 N_A3_c_283_n N_Y_c_664_n 0.00607661f $X=5.185 $Y=1.605 $X2=0 $Y2=0
cc_269 N_A3_c_285_n N_Y_c_719_n 0.00772049f $X=5.075 $Y=1.765 $X2=0 $Y2=0
cc_270 N_A3_c_286_n N_Y_c_719_n 5.50646e-19 $X=5.595 $Y=1.765 $X2=0 $Y2=0
cc_271 N_A3_c_285_n N_Y_c_721_n 0.0130869f $X=5.075 $Y=1.765 $X2=0 $Y2=0
cc_272 N_A3_c_286_n N_Y_c_721_n 0.0134861f $X=5.595 $Y=1.765 $X2=0 $Y2=0
cc_273 N_A3_c_282_n N_Y_c_721_n 0.00161525f $X=6.225 $Y=1.557 $X2=0 $Y2=0
cc_274 N_A3_c_290_n N_Y_c_721_n 0.0346905f $X=5.535 $Y=1.605 $X2=0 $Y2=0
cc_275 N_A3_c_283_n N_Y_c_721_n 0.00646699f $X=5.185 $Y=1.605 $X2=0 $Y2=0
cc_276 N_A3_c_287_n N_Y_c_726_n 0.0186112f $X=6.225 $Y=1.765 $X2=0 $Y2=0
cc_277 N_A3_c_288_n N_Y_c_726_n 0.0116961f $X=6.03 $Y=1.515 $X2=0 $Y2=0
cc_278 N_A3_c_282_n N_Y_c_726_n 5.7246e-19 $X=6.225 $Y=1.557 $X2=0 $Y2=0
cc_279 N_A3_c_284_n N_Y_c_666_n 0.00113906f $X=4.575 $Y=1.765 $X2=0 $Y2=0
cc_280 N_A3_c_285_n N_Y_c_666_n 0.00314498f $X=5.075 $Y=1.765 $X2=0 $Y2=0
cc_281 N_A3_c_286_n N_Y_c_666_n 5.991e-19 $X=5.595 $Y=1.765 $X2=0 $Y2=0
cc_282 N_A3_c_282_n N_Y_c_666_n 0.00870061f $X=6.225 $Y=1.557 $X2=0 $Y2=0
cc_283 N_A3_c_283_n N_Y_c_666_n 0.0257919f $X=5.185 $Y=1.605 $X2=0 $Y2=0
cc_284 N_A3_c_287_n N_Y_c_734_n 0.00889247f $X=6.225 $Y=1.765 $X2=0 $Y2=0
cc_285 N_A3_c_288_n N_Y_c_734_n 0.0268461f $X=6.03 $Y=1.515 $X2=0 $Y2=0
cc_286 N_A3_c_282_n N_Y_c_734_n 0.00190833f $X=6.225 $Y=1.557 $X2=0 $Y2=0
cc_287 N_A3_c_287_n Y 0.00439011f $X=6.225 $Y=1.765 $X2=0 $Y2=0
cc_288 N_A3_M1031_g Y 0.00747751f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_289 N_A3_c_288_n Y 0.0283828f $X=6.03 $Y=1.515 $X2=0 $Y2=0
cc_290 N_A3_c_284_n N_A_841_368#_c_796_n 0.00769091f $X=4.575 $Y=1.765 $X2=0
+ $Y2=0
cc_291 N_A3_c_285_n N_A_841_368#_c_796_n 2.69714e-19 $X=5.075 $Y=1.765 $X2=0
+ $Y2=0
cc_292 N_A3_c_284_n N_A_841_368#_c_797_n 0.0111147f $X=4.575 $Y=1.765 $X2=0
+ $Y2=0
cc_293 N_A3_c_285_n N_A_841_368#_c_797_n 0.0142264f $X=5.075 $Y=1.765 $X2=0
+ $Y2=0
cc_294 N_A3_c_284_n N_A_841_368#_c_798_n 0.00262934f $X=4.575 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A3_c_286_n N_A_841_368#_c_799_n 0.0143474f $X=5.595 $Y=1.765 $X2=0
+ $Y2=0
cc_296 N_A3_c_287_n N_A_841_368#_c_799_n 0.011675f $X=6.225 $Y=1.765 $X2=0 $Y2=0
cc_297 N_A3_c_286_n N_A_841_368#_c_813_n 7.79236e-19 $X=5.595 $Y=1.765 $X2=0
+ $Y2=0
cc_298 N_A3_c_287_n N_A_841_368#_c_813_n 0.00905158f $X=6.225 $Y=1.765 $X2=0
+ $Y2=0
cc_299 N_A3_c_287_n N_A_841_368#_c_804_n 0.00171731f $X=6.225 $Y=1.765 $X2=0
+ $Y2=0
cc_300 N_A3_M1008_g N_A_459_74#_c_963_n 5.29638e-19 $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_301 N_A3_M1008_g N_A_459_74#_c_964_n 0.00284982f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_302 N_A3_M1008_g N_A_459_74#_c_965_n 0.0128625f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_303 N_A3_M1008_g N_A_459_74#_c_967_n 4.39567e-19 $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_304 N_A3_M1010_g N_A_459_74#_c_967_n 0.00688453f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_305 N_A3_M1024_g N_A_459_74#_c_967_n 8.14332e-19 $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_306 N_A3_M1010_g N_A_459_74#_c_991_n 0.0095689f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A3_M1024_g N_A_459_74#_c_991_n 0.0095689f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_308 N_A3_M1010_g N_A_459_74#_c_968_n 8.11586e-19 $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A3_M1024_g N_A_459_74#_c_968_n 0.00724443f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_310 N_A3_M1031_g N_A_459_74#_c_968_n 0.0072728f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_311 N_A3_M1031_g N_A_459_74#_c_996_n 0.00947961f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A3_M1031_g N_A_459_74#_c_969_n 8.13633e-19 $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_313 N_A3_M1010_g N_A_459_74#_c_998_n 0.00181289f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A3_M1024_g N_A_459_74#_c_999_n 0.00181289f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A3_M1031_g N_A_459_74#_c_999_n 0.00181289f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A3_M1031_g N_A_459_74#_c_977_n 9.18816e-19 $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A3_M1008_g N_VGND_c_1112_n 0.0078527f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A3_M1010_g N_VGND_c_1112_n 4.46147e-19 $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_319 N_A3_M1010_g N_VGND_c_1113_n 0.00320743f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A3_M1024_g N_VGND_c_1113_n 0.00465809f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_321 N_A3_M1031_g N_VGND_c_1114_n 0.00471422f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_322 N_A3_M1008_g N_VGND_c_1120_n 0.00281141f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_323 N_A3_M1010_g N_VGND_c_1120_n 0.00331438f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_324 N_A3_M1024_g N_VGND_c_1121_n 0.00331438f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_325 N_A3_M1031_g N_VGND_c_1121_n 0.00331438f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_326 N_A3_M1008_g N_VGND_c_1132_n 0.00365066f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_327 N_A3_M1010_g N_VGND_c_1132_n 0.00427695f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_328 N_A3_M1024_g N_VGND_c_1132_n 0.00427695f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_329 N_A3_M1031_g N_VGND_c_1132_n 0.00427774f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_330 N_A2_c_379_n N_A1_M1005_g 0.0181944f $X=8.245 $Y=1.2 $X2=0 $Y2=0
cc_331 N_A2_c_380_n N_A1_M1005_g 0.0152468f $X=8.175 $Y=1.482 $X2=0 $Y2=0
cc_332 N_A2_c_384_n N_VPWR_c_550_n 0.0018633f $X=8.175 $Y=1.765 $X2=0 $Y2=0
cc_333 N_A2_c_381_n N_VPWR_c_556_n 0.00278257f $X=6.675 $Y=1.765 $X2=0 $Y2=0
cc_334 N_A2_c_382_n N_VPWR_c_556_n 0.00278271f $X=7.175 $Y=1.765 $X2=0 $Y2=0
cc_335 N_A2_c_383_n N_VPWR_c_556_n 0.00278271f $X=7.725 $Y=1.765 $X2=0 $Y2=0
cc_336 N_A2_c_384_n N_VPWR_c_556_n 0.00278257f $X=8.175 $Y=1.765 $X2=0 $Y2=0
cc_337 N_A2_c_381_n N_VPWR_c_546_n 0.00354366f $X=6.675 $Y=1.765 $X2=0 $Y2=0
cc_338 N_A2_c_382_n N_VPWR_c_546_n 0.00355164f $X=7.175 $Y=1.765 $X2=0 $Y2=0
cc_339 N_A2_c_383_n N_VPWR_c_546_n 0.00354703f $X=7.725 $Y=1.765 $X2=0 $Y2=0
cc_340 N_A2_c_384_n N_VPWR_c_546_n 0.00358623f $X=8.175 $Y=1.765 $X2=0 $Y2=0
cc_341 N_A2_M1001_g N_Y_c_660_n 0.00324583f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_342 N_A2_c_381_n Y 0.00229578f $X=6.675 $Y=1.765 $X2=0 $Y2=0
cc_343 N_A2_M1001_g Y 0.00210281f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_344 N_A2_c_385_n Y 0.0334136f $X=7.61 $Y=1.515 $X2=0 $Y2=0
cc_345 N_A2_c_380_n Y 0.0100548f $X=8.175 $Y=1.482 $X2=0 $Y2=0
cc_346 N_A2_c_381_n N_A_841_368#_c_813_n 0.00817736f $X=6.675 $Y=1.765 $X2=0
+ $Y2=0
cc_347 N_A2_c_382_n N_A_841_368#_c_813_n 5.85804e-19 $X=7.175 $Y=1.765 $X2=0
+ $Y2=0
cc_348 N_A2_c_381_n N_A_841_368#_c_800_n 0.0111147f $X=6.675 $Y=1.765 $X2=0
+ $Y2=0
cc_349 N_A2_c_382_n N_A_841_368#_c_800_n 0.0143659f $X=7.175 $Y=1.765 $X2=0
+ $Y2=0
cc_350 N_A2_c_383_n N_A_841_368#_c_801_n 0.0140926f $X=7.725 $Y=1.765 $X2=0
+ $Y2=0
cc_351 N_A2_c_384_n N_A_841_368#_c_801_n 0.0134708f $X=8.175 $Y=1.765 $X2=0
+ $Y2=0
cc_352 N_A2_c_383_n N_A_841_368#_c_802_n 5.71076e-19 $X=7.725 $Y=1.765 $X2=0
+ $Y2=0
cc_353 N_A2_c_384_n N_A_841_368#_c_802_n 0.00731604f $X=8.175 $Y=1.765 $X2=0
+ $Y2=0
cc_354 N_A2_c_381_n N_A_841_368#_c_804_n 0.00171731f $X=6.675 $Y=1.765 $X2=0
+ $Y2=0
cc_355 N_A2_c_382_n N_A_1350_368#_c_870_n 0.0125195f $X=7.175 $Y=1.765 $X2=0
+ $Y2=0
cc_356 N_A2_c_383_n N_A_1350_368#_c_870_n 0.0127944f $X=7.725 $Y=1.765 $X2=0
+ $Y2=0
cc_357 N_A2_c_385_n N_A_1350_368#_c_870_n 0.0466568f $X=7.61 $Y=1.515 $X2=0
+ $Y2=0
cc_358 N_A2_c_380_n N_A_1350_368#_c_870_n 0.00184966f $X=8.175 $Y=1.482 $X2=0
+ $Y2=0
cc_359 N_A2_c_382_n N_A_1350_368#_c_874_n 5.2199e-19 $X=7.175 $Y=1.765 $X2=0
+ $Y2=0
cc_360 N_A2_c_383_n N_A_1350_368#_c_874_n 0.00868111f $X=7.725 $Y=1.765 $X2=0
+ $Y2=0
cc_361 N_A2_c_384_n N_A_1350_368#_c_867_n 0.0174411f $X=8.175 $Y=1.765 $X2=0
+ $Y2=0
cc_362 N_A2_c_382_n N_A_1350_368#_c_877_n 0.0089318f $X=7.175 $Y=1.765 $X2=0
+ $Y2=0
cc_363 N_A2_c_383_n N_A_1350_368#_c_877_n 6.13607e-19 $X=7.725 $Y=1.765 $X2=0
+ $Y2=0
cc_364 N_A2_c_385_n N_A_1350_368#_c_877_n 0.025478f $X=7.61 $Y=1.515 $X2=0 $Y2=0
cc_365 N_A2_c_380_n N_A_1350_368#_c_877_n 0.00167317f $X=8.175 $Y=1.482 $X2=0
+ $Y2=0
cc_366 N_A2_c_383_n N_A_1350_368#_c_881_n 0.00153983f $X=7.725 $Y=1.765 $X2=0
+ $Y2=0
cc_367 N_A2_c_380_n N_A_1350_368#_c_881_n 0.00727992f $X=8.175 $Y=1.482 $X2=0
+ $Y2=0
cc_368 N_A2_M1001_g N_A_459_74#_c_968_n 8.06429e-19 $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_369 N_A2_M1001_g N_A_459_74#_c_996_n 0.0114917f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_370 N_A2_c_385_n N_A_459_74#_c_996_n 0.00430774f $X=7.61 $Y=1.515 $X2=0 $Y2=0
cc_371 N_A2_c_380_n N_A_459_74#_c_996_n 0.00462064f $X=8.175 $Y=1.482 $X2=0
+ $Y2=0
cc_372 N_A2_M1001_g N_A_459_74#_c_969_n 0.00661943f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_373 N_A2_M1004_g N_A_459_74#_c_969_n 3.97481e-19 $X=7.27 $Y=0.74 $X2=0 $Y2=0
cc_374 N_A2_M1004_g N_A_459_74#_c_970_n 0.0127949f $X=7.27 $Y=0.74 $X2=0 $Y2=0
cc_375 N_A2_c_378_n N_A_459_74#_c_970_n 0.015874f $X=7.74 $Y=1.2 $X2=0 $Y2=0
cc_376 N_A2_c_385_n N_A_459_74#_c_970_n 0.0477395f $X=7.61 $Y=1.515 $X2=0 $Y2=0
cc_377 N_A2_c_380_n N_A_459_74#_c_970_n 0.00497406f $X=8.175 $Y=1.482 $X2=0
+ $Y2=0
cc_378 N_A2_c_378_n N_A_459_74#_c_971_n 0.00814722f $X=7.74 $Y=1.2 $X2=0 $Y2=0
cc_379 N_A2_c_379_n N_A_459_74#_c_971_n 0.00156085f $X=8.245 $Y=1.2 $X2=0 $Y2=0
cc_380 N_A2_c_380_n N_A_459_74#_c_972_n 0.0183445f $X=8.175 $Y=1.482 $X2=0 $Y2=0
cc_381 N_A2_c_379_n N_A_459_74#_c_973_n 2.1934e-19 $X=8.245 $Y=1.2 $X2=0 $Y2=0
cc_382 N_A2_c_379_n N_A_459_74#_c_974_n 6.00311e-19 $X=8.245 $Y=1.2 $X2=0 $Y2=0
cc_383 N_A2_M1001_g N_A_459_74#_c_977_n 0.00668147f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_384 N_A2_c_385_n N_A_459_74#_c_977_n 0.0211953f $X=7.61 $Y=1.515 $X2=0 $Y2=0
cc_385 N_A2_c_380_n N_A_459_74#_c_977_n 0.00236559f $X=8.175 $Y=1.482 $X2=0
+ $Y2=0
cc_386 N_A2_M1004_g N_A_459_74#_c_978_n 5.55763e-19 $X=7.27 $Y=0.74 $X2=0 $Y2=0
cc_387 N_A2_c_378_n N_A_459_74#_c_978_n 7.16428e-19 $X=7.74 $Y=1.2 $X2=0 $Y2=0
cc_388 N_A2_c_385_n N_A_459_74#_c_978_n 0.00906486f $X=7.61 $Y=1.515 $X2=0 $Y2=0
cc_389 N_A2_c_380_n N_A_459_74#_c_978_n 0.01739f $X=8.175 $Y=1.482 $X2=0 $Y2=0
cc_390 N_A2_M1001_g N_VGND_c_1114_n 0.00325376f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_391 N_A2_M1001_g N_VGND_c_1115_n 5.16425e-19 $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_392 N_A2_M1004_g N_VGND_c_1115_n 0.0103635f $X=7.27 $Y=0.74 $X2=0 $Y2=0
cc_393 N_A2_c_378_n N_VGND_c_1115_n 0.00243974f $X=7.74 $Y=1.2 $X2=0 $Y2=0
cc_394 N_A2_c_378_n N_VGND_c_1116_n 5.07467e-19 $X=7.74 $Y=1.2 $X2=0 $Y2=0
cc_395 N_A2_c_379_n N_VGND_c_1116_n 0.0130384f $X=8.245 $Y=1.2 $X2=0 $Y2=0
cc_396 N_A2_M1001_g N_VGND_c_1122_n 0.00331438f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_397 N_A2_M1004_g N_VGND_c_1122_n 0.00383152f $X=7.27 $Y=0.74 $X2=0 $Y2=0
cc_398 N_A2_c_378_n N_VGND_c_1123_n 0.00461464f $X=7.74 $Y=1.2 $X2=0 $Y2=0
cc_399 N_A2_c_379_n N_VGND_c_1123_n 0.00383152f $X=8.245 $Y=1.2 $X2=0 $Y2=0
cc_400 N_A2_M1001_g N_VGND_c_1132_n 0.00427774f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_401 N_A2_M1004_g N_VGND_c_1132_n 0.0075754f $X=7.27 $Y=0.74 $X2=0 $Y2=0
cc_402 N_A2_c_378_n N_VGND_c_1132_n 0.00908525f $X=7.74 $Y=1.2 $X2=0 $Y2=0
cc_403 N_A2_c_379_n N_VGND_c_1132_n 0.00758242f $X=8.245 $Y=1.2 $X2=0 $Y2=0
cc_404 N_A1_c_474_n N_VPWR_c_550_n 0.0113689f $X=9.185 $Y=1.765 $X2=0 $Y2=0
cc_405 N_A1_c_475_n N_VPWR_c_550_n 4.96035e-19 $X=9.635 $Y=1.765 $X2=0 $Y2=0
cc_406 N_A1_c_474_n N_VPWR_c_551_n 4.96035e-19 $X=9.185 $Y=1.765 $X2=0 $Y2=0
cc_407 N_A1_c_475_n N_VPWR_c_551_n 0.0103012f $X=9.635 $Y=1.765 $X2=0 $Y2=0
cc_408 N_A1_c_476_n N_VPWR_c_551_n 0.0104324f $X=10.085 $Y=1.765 $X2=0 $Y2=0
cc_409 N_A1_c_477_n N_VPWR_c_551_n 5.15164e-19 $X=10.535 $Y=1.765 $X2=0 $Y2=0
cc_410 N_A1_c_477_n N_VPWR_c_553_n 0.011094f $X=10.535 $Y=1.765 $X2=0 $Y2=0
cc_411 N_A1_c_474_n N_VPWR_c_557_n 0.00413917f $X=9.185 $Y=1.765 $X2=0 $Y2=0
cc_412 N_A1_c_475_n N_VPWR_c_557_n 0.00413917f $X=9.635 $Y=1.765 $X2=0 $Y2=0
cc_413 N_A1_c_476_n N_VPWR_c_558_n 0.00413917f $X=10.085 $Y=1.765 $X2=0 $Y2=0
cc_414 N_A1_c_477_n N_VPWR_c_558_n 0.00445602f $X=10.535 $Y=1.765 $X2=0 $Y2=0
cc_415 N_A1_c_474_n N_VPWR_c_546_n 0.00817726f $X=9.185 $Y=1.765 $X2=0 $Y2=0
cc_416 N_A1_c_475_n N_VPWR_c_546_n 0.00817726f $X=9.635 $Y=1.765 $X2=0 $Y2=0
cc_417 N_A1_c_476_n N_VPWR_c_546_n 0.00817726f $X=10.085 $Y=1.765 $X2=0 $Y2=0
cc_418 N_A1_c_477_n N_VPWR_c_546_n 0.00861084f $X=10.535 $Y=1.765 $X2=0 $Y2=0
cc_419 N_A1_c_474_n N_A_841_368#_c_801_n 5.94256e-19 $X=9.185 $Y=1.765 $X2=0
+ $Y2=0
cc_420 N_A1_c_474_n N_A_841_368#_c_802_n 0.00100131f $X=9.185 $Y=1.765 $X2=0
+ $Y2=0
cc_421 N_A1_c_467_n N_A_1350_368#_c_867_n 0.0130812f $X=8.75 $Y=1.605 $X2=0
+ $Y2=0
cc_422 N_A1_c_474_n N_A_1350_368#_c_867_n 0.0176052f $X=9.185 $Y=1.765 $X2=0
+ $Y2=0
cc_423 N_A1_c_478_n N_A_1350_368#_c_867_n 0.00849498f $X=10.35 $Y=1.515 $X2=0
+ $Y2=0
cc_424 N_A1_c_474_n N_A_1350_368#_c_868_n 2.92088e-19 $X=9.185 $Y=1.765 $X2=0
+ $Y2=0
cc_425 N_A1_c_475_n N_A_1350_368#_c_868_n 2.92088e-19 $X=9.635 $Y=1.765 $X2=0
+ $Y2=0
cc_426 N_A1_c_475_n N_A_1350_368#_c_888_n 0.0136211f $X=9.635 $Y=1.765 $X2=0
+ $Y2=0
cc_427 N_A1_c_476_n N_A_1350_368#_c_888_n 0.0136211f $X=10.085 $Y=1.765 $X2=0
+ $Y2=0
cc_428 N_A1_c_478_n N_A_1350_368#_c_888_n 0.0450321f $X=10.35 $Y=1.515 $X2=0
+ $Y2=0
cc_429 N_A1_c_471_n N_A_1350_368#_c_888_n 0.00132918f $X=10.535 $Y=1.482 $X2=0
+ $Y2=0
cc_430 N_A1_c_477_n N_A_1350_368#_c_892_n 0.00288396f $X=10.535 $Y=1.765 $X2=0
+ $Y2=0
cc_431 N_A1_c_478_n N_A_1350_368#_c_892_n 0.0187917f $X=10.35 $Y=1.515 $X2=0
+ $Y2=0
cc_432 N_A1_c_471_n N_A_1350_368#_c_892_n 0.00133119f $X=10.535 $Y=1.482 $X2=0
+ $Y2=0
cc_433 N_A1_c_476_n N_A_1350_368#_c_869_n 2.94821e-19 $X=10.085 $Y=1.765 $X2=0
+ $Y2=0
cc_434 N_A1_c_477_n N_A_1350_368#_c_869_n 0.00955117f $X=10.535 $Y=1.765 $X2=0
+ $Y2=0
cc_435 N_A1_c_478_n N_A_1350_368#_c_897_n 0.0183565f $X=10.35 $Y=1.515 $X2=0
+ $Y2=0
cc_436 N_A1_c_471_n N_A_1350_368#_c_897_n 0.0013074f $X=10.535 $Y=1.482 $X2=0
+ $Y2=0
cc_437 N_A1_M1005_g N_A_459_74#_c_972_n 0.0142591f $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_438 N_A1_c_466_n N_A_459_74#_c_972_n 0.00285025f $X=9.03 $Y=1.605 $X2=0 $Y2=0
cc_439 N_A1_M1012_g N_A_459_74#_c_972_n 0.0028354f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_440 N_A1_c_478_n N_A_459_74#_c_972_n 0.00974864f $X=10.35 $Y=1.515 $X2=0
+ $Y2=0
cc_441 N_A1_M1005_g N_A_459_74#_c_973_n 0.00725305f $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_442 N_A1_M1012_g N_A_459_74#_c_973_n 3.97173e-19 $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_443 N_A1_M1005_g N_A_459_74#_c_974_n 0.00467801f $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_444 N_A1_M1012_g N_A_459_74#_c_974_n 0.00432461f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_445 N_A1_M1012_g N_A_459_74#_c_975_n 0.0184943f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_446 N_A1_c_469_n N_A_459_74#_c_975_n 0.0150704f $X=10.1 $Y=1.2 $X2=0 $Y2=0
cc_447 N_A1_c_478_n N_A_459_74#_c_975_n 0.0802473f $X=10.35 $Y=1.515 $X2=0 $Y2=0
cc_448 N_A1_c_471_n N_A_459_74#_c_975_n 0.0183904f $X=10.535 $Y=1.482 $X2=0
+ $Y2=0
cc_449 N_A1_c_469_n N_A_459_74#_c_976_n 0.0120086f $X=10.1 $Y=1.2 $X2=0 $Y2=0
cc_450 N_A1_c_470_n N_A_459_74#_c_976_n 4.13268e-19 $X=10.545 $Y=1.2 $X2=0 $Y2=0
cc_451 N_A1_M1005_g N_A_459_74#_c_978_n 3.35826e-19 $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_452 N_A1_M1005_g N_A_459_74#_c_1039_n 0.00199342f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_453 N_A1_M1005_g N_VGND_c_1116_n 0.0019818f $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_454 N_A1_c_469_n N_VGND_c_1118_n 6.05373e-19 $X=10.1 $Y=1.2 $X2=0 $Y2=0
cc_455 N_A1_c_470_n N_VGND_c_1118_n 0.0160304f $X=10.545 $Y=1.2 $X2=0 $Y2=0
cc_456 N_A1_c_471_n N_VGND_c_1118_n 2.15716e-19 $X=10.535 $Y=1.482 $X2=0 $Y2=0
cc_457 N_A1_c_469_n N_VGND_c_1124_n 0.00451267f $X=10.1 $Y=1.2 $X2=0 $Y2=0
cc_458 N_A1_c_470_n N_VGND_c_1124_n 0.00383152f $X=10.545 $Y=1.2 $X2=0 $Y2=0
cc_459 N_A1_M1005_g N_VGND_c_1130_n 0.00434272f $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_460 N_A1_M1012_g N_VGND_c_1130_n 0.00383152f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_461 N_A1_M1005_g N_VGND_c_1131_n 5.00706e-19 $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_462 N_A1_M1012_g N_VGND_c_1131_n 0.0120529f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_463 N_A1_c_469_n N_VGND_c_1131_n 0.00510378f $X=10.1 $Y=1.2 $X2=0 $Y2=0
cc_464 N_A1_M1005_g N_VGND_c_1132_n 0.00820382f $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_465 N_A1_M1012_g N_VGND_c_1132_n 0.00752925f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_466 N_A1_c_469_n N_VGND_c_1132_n 0.00879879f $X=10.1 $Y=1.2 $X2=0 $Y2=0
cc_467 N_A1_c_470_n N_VGND_c_1132_n 0.00757689f $X=10.545 $Y=1.2 $X2=0 $Y2=0
cc_468 N_VPWR_c_548_n N_Y_c_668_n 0.00919225f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_469 N_VPWR_c_548_n N_Y_c_662_n 0.043762f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_470 N_VPWR_c_549_n N_Y_c_662_n 0.0266809f $X=1.405 $Y=2.455 $X2=0 $Y2=0
cc_471 N_VPWR_c_554_n N_Y_c_662_n 0.0146357f $X=1.24 $Y=3.33 $X2=0 $Y2=0
cc_472 N_VPWR_c_546_n N_Y_c_662_n 0.0121141f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_473 N_VPWR_M1022_d N_Y_c_673_n 0.00651362f $X=1.255 $Y=1.84 $X2=0 $Y2=0
cc_474 N_VPWR_c_549_n N_Y_c_673_n 0.0202249f $X=1.405 $Y=2.455 $X2=0 $Y2=0
cc_475 N_VPWR_c_549_n N_Y_c_663_n 0.0266809f $X=1.405 $Y=2.455 $X2=0 $Y2=0
cc_476 N_VPWR_c_559_n N_Y_c_663_n 0.014552f $X=2.24 $Y=2.852 $X2=0 $Y2=0
cc_477 N_VPWR_c_560_n N_Y_c_663_n 0.0268614f $X=3.905 $Y=2.852 $X2=0 $Y2=0
cc_478 N_VPWR_c_546_n N_Y_c_663_n 0.0119791f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_479 N_VPWR_M1028_s N_Y_c_664_n 0.0461734f $X=2.205 $Y=1.84 $X2=0 $Y2=0
cc_480 N_VPWR_c_560_n N_Y_c_664_n 0.133101f $X=3.905 $Y=2.852 $X2=0 $Y2=0
cc_481 N_VPWR_c_560_n N_A_841_368#_c_796_n 0.0383128f $X=3.905 $Y=2.852 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_556_n N_A_841_368#_c_797_n 0.0422753f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_546_n N_A_841_368#_c_797_n 0.0238861f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_484 N_VPWR_c_556_n N_A_841_368#_c_798_n 0.0236039f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_560_n N_A_841_368#_c_798_n 0.0112249f $X=3.905 $Y=2.852 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_546_n N_A_841_368#_c_798_n 0.012761f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_487 N_VPWR_c_556_n N_A_841_368#_c_799_n 0.0487171f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_546_n N_A_841_368#_c_799_n 0.0276459f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_556_n N_A_841_368#_c_800_n 0.0422753f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_546_n N_A_841_368#_c_800_n 0.0238861f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_550_n N_A_841_368#_c_801_n 0.0121617f $X=8.96 $Y=2.415 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_556_n N_A_841_368#_c_801_n 0.0626582f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_546_n N_A_841_368#_c_801_n 0.0347672f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_550_n N_A_841_368#_c_802_n 0.038732f $X=8.96 $Y=2.415 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_556_n N_A_841_368#_c_803_n 0.0236566f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_546_n N_A_841_368#_c_803_n 0.0128296f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_556_n N_A_841_368#_c_804_n 0.0235512f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_546_n N_A_841_368#_c_804_n 0.0126924f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_556_n N_A_841_368#_c_805_n 0.0236566f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_546_n N_A_841_368#_c_805_n 0.0128296f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_501 N_VPWR_M1007_d N_A_1350_368#_c_867_n 0.00703016f $X=8.815 $Y=1.84 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_550_n N_A_1350_368#_c_867_n 0.0213061f $X=8.96 $Y=2.415 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_550_n N_A_1350_368#_c_868_n 0.025138f $X=8.96 $Y=2.415 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_551_n N_A_1350_368#_c_868_n 0.025138f $X=9.86 $Y=2.415 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_557_n N_A_1350_368#_c_868_n 0.0101736f $X=9.695 $Y=3.33 $X2=0
+ $Y2=0
cc_506 N_VPWR_c_546_n N_A_1350_368#_c_868_n 0.0084208f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_507 N_VPWR_M1013_d N_A_1350_368#_c_888_n 0.00366f $X=9.71 $Y=1.84 $X2=0 $Y2=0
cc_508 N_VPWR_c_551_n N_A_1350_368#_c_888_n 0.0166391f $X=9.86 $Y=2.415 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_553_n N_A_1350_368#_c_892_n 0.0142382f $X=10.76 $Y=1.985 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_551_n N_A_1350_368#_c_869_n 0.0251606f $X=9.86 $Y=2.415 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_553_n N_A_1350_368#_c_869_n 0.0549702f $X=10.76 $Y=1.985 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_558_n N_A_1350_368#_c_869_n 0.0123628f $X=10.675 $Y=3.33 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_546_n N_A_1350_368#_c_869_n 0.0101999f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_514 N_Y_c_664_n N_A_841_368#_M1000_d 0.0126804f $X=4.685 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_515 N_Y_c_721_n N_A_841_368#_M1009_d 0.00503909f $X=5.685 $Y=2.035 $X2=0
+ $Y2=0
cc_516 N_Y_c_726_n N_A_841_368#_M1032_d 0.00285816f $X=6.365 $Y=2.035 $X2=0
+ $Y2=0
cc_517 Y N_A_841_368#_M1032_d 0.00125935f $X=6.48 $Y=1.295 $X2=0 $Y2=0
cc_518 N_Y_c_664_n N_A_841_368#_c_796_n 0.0219924f $X=4.685 $Y=2.035 $X2=0 $Y2=0
cc_519 N_Y_M1000_s N_A_841_368#_c_797_n 0.00250873f $X=4.65 $Y=1.84 $X2=0 $Y2=0
cc_520 N_Y_c_719_n N_A_841_368#_c_797_n 0.018923f $X=4.85 $Y=2.31 $X2=0 $Y2=0
cc_521 N_Y_c_721_n N_A_841_368#_c_854_n 0.0208278f $X=5.685 $Y=2.035 $X2=0 $Y2=0
cc_522 N_Y_M1030_s N_A_841_368#_c_799_n 0.00642382f $X=5.67 $Y=1.84 $X2=0 $Y2=0
cc_523 N_Y_c_734_n N_A_841_368#_c_799_n 0.0218444f $X=5.85 $Y=2.115 $X2=0 $Y2=0
cc_524 N_Y_c_726_n N_A_841_368#_c_813_n 0.0176424f $X=6.365 $Y=2.035 $X2=0 $Y2=0
cc_525 N_Y_c_734_n N_A_841_368#_c_813_n 0.0242295f $X=5.85 $Y=2.115 $X2=0 $Y2=0
cc_526 N_Y_c_680_n N_A_27_74#_M1018_s 0.00342755f $X=1.41 $Y=1.015 $X2=0 $Y2=0
cc_527 N_Y_c_659_n N_A_27_74#_M1029_s 0.00176461f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_528 N_Y_c_659_n N_A_27_74#_M1014_s 0.00176891f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_529 N_Y_c_659_n N_A_27_74#_M1027_s 0.00213024f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_530 N_Y_M1003_d N_A_27_74#_c_925_n 0.00174304f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_531 N_Y_M1019_d N_A_27_74#_c_925_n 0.00169393f $X=1.435 $Y=0.37 $X2=0 $Y2=0
cc_532 N_Y_c_659_n N_A_27_74#_c_925_n 0.0036578f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_533 N_Y_c_680_n N_A_27_74#_c_925_n 0.0633287f $X=1.41 $Y=1.015 $X2=0 $Y2=0
cc_534 N_Y_c_659_n N_A_27_74#_c_948_n 0.0133131f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_535 N_Y_c_659_n N_A_27_74#_c_926_n 0.0955773f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_536 N_Y_c_659_n N_A_459_74#_M1002_d 0.00176891f $X=6.365 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_537 N_Y_c_659_n N_A_459_74#_M1015_d 0.00187547f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_538 N_Y_c_659_n N_A_459_74#_M1008_s 0.00176461f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_539 N_Y_c_659_n N_A_459_74#_M1024_s 0.00176461f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_540 N_Y_c_659_n N_A_459_74#_c_963_n 0.0061464f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_541 N_Y_c_659_n N_A_459_74#_c_965_n 0.0410903f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_542 N_Y_c_659_n N_A_459_74#_c_966_n 0.0141908f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_543 N_Y_c_659_n N_A_459_74#_c_991_n 0.0405558f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_544 N_Y_c_659_n N_A_459_74#_c_996_n 0.00843866f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_545 N_Y_c_660_n N_A_459_74#_c_996_n 0.018143f $X=6.48 $Y=1.26 $X2=0 $Y2=0
cc_546 N_Y_c_659_n N_A_459_74#_c_998_n 0.0151907f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_547 N_Y_c_659_n N_A_459_74#_c_999_n 0.0170682f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_548 N_Y_c_660_n N_A_459_74#_c_977_n 0.00490592f $X=6.48 $Y=1.26 $X2=0 $Y2=0
cc_549 N_Y_c_659_n N_VGND_M1008_d 0.00213024f $X=6.365 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_550 N_Y_c_659_n N_VGND_M1010_d 0.00355802f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_551 N_Y_c_660_n N_VGND_M1031_d 0.002798f $X=6.48 $Y=1.26 $X2=0 $Y2=0
cc_552 N_A_841_368#_c_800_n N_A_1350_368#_M1006_s 0.00250873f $X=7.285 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_553 N_A_841_368#_c_801_n N_A_1350_368#_M1026_s 0.00197722f $X=8.235 $Y=2.99
+ $X2=0 $Y2=0
cc_554 N_A_841_368#_M1021_d N_A_1350_368#_c_870_n 0.00589767f $X=7.25 $Y=1.84
+ $X2=0 $Y2=0
cc_555 N_A_841_368#_c_862_p N_A_1350_368#_c_870_n 0.0232685f $X=7.45 $Y=2.455
+ $X2=0 $Y2=0
cc_556 N_A_841_368#_c_801_n N_A_1350_368#_c_874_n 0.0151173f $X=8.235 $Y=2.99
+ $X2=0 $Y2=0
cc_557 N_A_841_368#_M1033_d N_A_1350_368#_c_867_n 0.00806595f $X=8.25 $Y=1.84
+ $X2=0 $Y2=0
cc_558 N_A_841_368#_c_802_n N_A_1350_368#_c_867_n 0.0213061f $X=8.4 $Y=2.415
+ $X2=0 $Y2=0
cc_559 N_A_841_368#_c_800_n N_A_1350_368#_c_877_n 0.018923f $X=7.285 $Y=2.99
+ $X2=0 $Y2=0
cc_560 N_A_1350_368#_c_867_n N_A_459_74#_c_972_n 0.0296443f $X=9.295 $Y=2.05
+ $X2=0 $Y2=0
cc_561 N_A_1350_368#_c_867_n N_A_459_74#_c_978_n 0.00107938f $X=9.295 $Y=2.05
+ $X2=0 $Y2=0
cc_562 N_A_1350_368#_c_881_n N_A_459_74#_c_978_n 0.0041686f $X=7.95 $Y=2.035
+ $X2=0 $Y2=0
cc_563 N_A_27_74#_c_926_n N_A_459_74#_M1002_d 0.00335829f $X=3.735 $Y=0.835
+ $X2=-0.19 $Y2=-0.245
cc_564 N_A_27_74#_c_926_n N_A_459_74#_M1015_d 0.003555f $X=3.735 $Y=0.835 $X2=0
+ $Y2=0
cc_565 N_A_27_74#_M1014_s N_A_459_74#_c_963_n 0.00179007f $X=2.725 $Y=0.37 $X2=0
+ $Y2=0
cc_566 N_A_27_74#_M1027_s N_A_459_74#_c_963_n 0.002891f $X=3.595 $Y=0.37 $X2=0
+ $Y2=0
cc_567 N_A_27_74#_c_925_n N_A_459_74#_c_963_n 0.0101071f $X=1.92 $Y=0.475 $X2=0
+ $Y2=0
cc_568 N_A_27_74#_c_926_n N_A_459_74#_c_963_n 0.0865605f $X=3.735 $Y=0.835 $X2=0
+ $Y2=0
cc_569 N_A_27_74#_c_926_n N_A_459_74#_c_966_n 0.015741f $X=3.735 $Y=0.835 $X2=0
+ $Y2=0
cc_570 N_A_27_74#_c_923_n N_VGND_c_1119_n 0.0111552f $X=0.24 $Y=0.6 $X2=0 $Y2=0
cc_571 N_A_27_74#_c_925_n N_VGND_c_1119_n 0.0702753f $X=1.92 $Y=0.475 $X2=0
+ $Y2=0
cc_572 N_A_27_74#_c_926_n N_VGND_c_1119_n 0.00197884f $X=3.735 $Y=0.835 $X2=0
+ $Y2=0
cc_573 N_A_27_74#_c_923_n N_VGND_c_1132_n 0.00923333f $X=0.24 $Y=0.6 $X2=0 $Y2=0
cc_574 N_A_27_74#_c_925_n N_VGND_c_1132_n 0.0589522f $X=1.92 $Y=0.475 $X2=0
+ $Y2=0
cc_575 N_A_27_74#_c_926_n N_VGND_c_1132_n 0.00654682f $X=3.735 $Y=0.835 $X2=0
+ $Y2=0
cc_576 N_A_459_74#_c_965_n N_VGND_M1008_d 0.00447087f $X=4.92 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_577 N_A_459_74#_c_991_n N_VGND_M1010_d 0.00724158f $X=5.86 $Y=0.835 $X2=0
+ $Y2=0
cc_578 N_A_459_74#_c_996_n N_VGND_M1031_d 0.00831277f $X=6.89 $Y=0.835 $X2=0
+ $Y2=0
cc_579 N_A_459_74#_c_970_n N_VGND_M1004_d 0.0022694f $X=7.945 $Y=1.095 $X2=0
+ $Y2=0
cc_580 N_A_459_74#_c_975_n N_VGND_M1012_d 0.0117895f $X=10.165 $Y=1.045 $X2=0
+ $Y2=0
cc_581 N_A_459_74#_c_963_n N_VGND_c_1112_n 0.0221151f $X=4.07 $Y=0.455 $X2=0
+ $Y2=0
cc_582 N_A_459_74#_c_965_n N_VGND_c_1112_n 0.0212697f $X=4.92 $Y=0.835 $X2=0
+ $Y2=0
cc_583 N_A_459_74#_c_967_n N_VGND_c_1112_n 0.00897147f $X=5.005 $Y=0.635 $X2=0
+ $Y2=0
cc_584 N_A_459_74#_c_967_n N_VGND_c_1113_n 0.00865936f $X=5.005 $Y=0.635 $X2=0
+ $Y2=0
cc_585 N_A_459_74#_c_991_n N_VGND_c_1113_n 0.0256608f $X=5.86 $Y=0.835 $X2=0
+ $Y2=0
cc_586 N_A_459_74#_c_968_n N_VGND_c_1113_n 0.00900273f $X=6.025 $Y=0.635 $X2=0
+ $Y2=0
cc_587 N_A_459_74#_c_968_n N_VGND_c_1114_n 0.00900616f $X=6.025 $Y=0.635 $X2=0
+ $Y2=0
cc_588 N_A_459_74#_c_996_n N_VGND_c_1114_n 0.0264479f $X=6.89 $Y=0.835 $X2=0
+ $Y2=0
cc_589 N_A_459_74#_c_969_n N_VGND_c_1114_n 0.0086628f $X=7.055 $Y=0.515 $X2=0
+ $Y2=0
cc_590 N_A_459_74#_c_969_n N_VGND_c_1115_n 0.0177526f $X=7.055 $Y=0.515 $X2=0
+ $Y2=0
cc_591 N_A_459_74#_c_970_n N_VGND_c_1115_n 0.017402f $X=7.945 $Y=1.095 $X2=0
+ $Y2=0
cc_592 N_A_459_74#_c_971_n N_VGND_c_1115_n 0.0120634f $X=8.03 $Y=0.515 $X2=0
+ $Y2=0
cc_593 N_A_459_74#_c_971_n N_VGND_c_1116_n 0.0281649f $X=8.03 $Y=0.515 $X2=0
+ $Y2=0
cc_594 N_A_459_74#_c_972_n N_VGND_c_1116_n 0.0207473f $X=8.725 $Y=1.385 $X2=0
+ $Y2=0
cc_595 N_A_459_74#_c_973_n N_VGND_c_1116_n 0.0216462f $X=8.89 $Y=0.515 $X2=0
+ $Y2=0
cc_596 N_A_459_74#_c_1039_n N_VGND_c_1116_n 0.00756924f $X=8.85 $Y=1.045 $X2=0
+ $Y2=0
cc_597 N_A_459_74#_c_975_n N_VGND_c_1118_n 0.00697079f $X=10.165 $Y=1.045 $X2=0
+ $Y2=0
cc_598 N_A_459_74#_c_976_n N_VGND_c_1118_n 0.0225912f $X=10.33 $Y=0.515 $X2=0
+ $Y2=0
cc_599 N_A_459_74#_c_963_n N_VGND_c_1119_n 0.0878111f $X=4.07 $Y=0.455 $X2=0
+ $Y2=0
cc_600 N_A_459_74#_c_965_n N_VGND_c_1119_n 0.0024506f $X=4.92 $Y=0.835 $X2=0
+ $Y2=0
cc_601 N_A_459_74#_c_965_n N_VGND_c_1120_n 0.00197156f $X=4.92 $Y=0.835 $X2=0
+ $Y2=0
cc_602 N_A_459_74#_c_967_n N_VGND_c_1120_n 0.0108551f $X=5.005 $Y=0.635 $X2=0
+ $Y2=0
cc_603 N_A_459_74#_c_991_n N_VGND_c_1120_n 0.00197156f $X=5.86 $Y=0.835 $X2=0
+ $Y2=0
cc_604 N_A_459_74#_c_991_n N_VGND_c_1121_n 0.00197156f $X=5.86 $Y=0.835 $X2=0
+ $Y2=0
cc_605 N_A_459_74#_c_968_n N_VGND_c_1121_n 0.0143093f $X=6.025 $Y=0.635 $X2=0
+ $Y2=0
cc_606 N_A_459_74#_c_996_n N_VGND_c_1121_n 0.00197156f $X=6.89 $Y=0.835 $X2=0
+ $Y2=0
cc_607 N_A_459_74#_c_996_n N_VGND_c_1122_n 0.00197695f $X=6.89 $Y=0.835 $X2=0
+ $Y2=0
cc_608 N_A_459_74#_c_969_n N_VGND_c_1122_n 0.0109942f $X=7.055 $Y=0.515 $X2=0
+ $Y2=0
cc_609 N_A_459_74#_c_971_n N_VGND_c_1123_n 0.00749631f $X=8.03 $Y=0.515 $X2=0
+ $Y2=0
cc_610 N_A_459_74#_c_976_n N_VGND_c_1124_n 0.0110391f $X=10.33 $Y=0.515 $X2=0
+ $Y2=0
cc_611 N_A_459_74#_c_973_n N_VGND_c_1130_n 0.0109942f $X=8.89 $Y=0.515 $X2=0
+ $Y2=0
cc_612 N_A_459_74#_c_973_n N_VGND_c_1131_n 0.01839f $X=8.89 $Y=0.515 $X2=0 $Y2=0
cc_613 N_A_459_74#_c_975_n N_VGND_c_1131_n 0.0610657f $X=10.165 $Y=1.045 $X2=0
+ $Y2=0
cc_614 N_A_459_74#_c_976_n N_VGND_c_1131_n 0.0167469f $X=10.33 $Y=0.515 $X2=0
+ $Y2=0
cc_615 N_A_459_74#_c_963_n N_VGND_c_1132_n 0.0692687f $X=4.07 $Y=0.455 $X2=0
+ $Y2=0
cc_616 N_A_459_74#_c_965_n N_VGND_c_1132_n 0.00976958f $X=4.92 $Y=0.835 $X2=0
+ $Y2=0
cc_617 N_A_459_74#_c_967_n N_VGND_c_1132_n 0.00898945f $X=5.005 $Y=0.635 $X2=0
+ $Y2=0
cc_618 N_A_459_74#_c_991_n N_VGND_c_1132_n 0.00943478f $X=5.86 $Y=0.835 $X2=0
+ $Y2=0
cc_619 N_A_459_74#_c_968_n N_VGND_c_1132_n 0.0118109f $X=6.025 $Y=0.635 $X2=0
+ $Y2=0
cc_620 N_A_459_74#_c_996_n N_VGND_c_1132_n 0.00947592f $X=6.89 $Y=0.835 $X2=0
+ $Y2=0
cc_621 N_A_459_74#_c_969_n N_VGND_c_1132_n 0.00904371f $X=7.055 $Y=0.515 $X2=0
+ $Y2=0
cc_622 N_A_459_74#_c_971_n N_VGND_c_1132_n 0.0062048f $X=8.03 $Y=0.515 $X2=0
+ $Y2=0
cc_623 N_A_459_74#_c_973_n N_VGND_c_1132_n 0.00904371f $X=8.89 $Y=0.515 $X2=0
+ $Y2=0
cc_624 N_A_459_74#_c_976_n N_VGND_c_1132_n 0.00911606f $X=10.33 $Y=0.515 $X2=0
+ $Y2=0
