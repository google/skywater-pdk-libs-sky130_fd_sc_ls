* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__or3b_4 A B C_N VGND VNB VPB VPWR X
M1000 X a_409_392# VGND VNB nshort w=740000u l=150000u
+  ad=4.329e+11p pd=4.13e+06u as=1.64125e+12p ps=1.215e+07u
M1001 X a_409_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=1.407e+12p ps=1.133e+07u
M1002 VPWR a_409_392# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_409_392# B VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1004 VGND a_409_392# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_27_392# a_409_392# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_307_392# a_27_392# a_409_392# VPB phighvt w=1e+06u l=150000u
+  ad=6.6e+11p pd=5.32e+06u as=3.25e+11p ps=2.65e+06u
M1007 a_217_392# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=6.6e+11p pd=5.32e+06u as=0p ps=0u
M1008 X a_409_392# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A a_409_392# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND C_N a_27_392# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1011 a_217_392# B a_307_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A a_217_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR C_N a_27_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1014 VGND a_409_392# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_307_392# B a_217_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_409_392# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_409_392# a_27_392# a_307_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_409_392# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
