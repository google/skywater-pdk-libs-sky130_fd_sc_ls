* NGSPICE file created from sky130_fd_sc_ls__a21o_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
M1000 X a_91_48# VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=1.011e+12p ps=9.9e+06u
M1001 a_503_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=1.15e+12p pd=1.03e+07u as=1.552e+12p ps=1.362e+07u
M1002 VPWR a_91_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.72e+11p ps=5.68e+06u
M1003 VPWR A2 a_503_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_91_48# B1 a_503_392# VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1005 a_503_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_700_74# A1 a_91_48# VNB nshort w=640000u l=150000u
+  ad=5.184e+11p pd=5.46e+06u as=3.584e+11p ps=3.68e+06u
M1007 X a_91_48# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_91_48# B1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_503_392# B1 a_91_48# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_91_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_91_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_91_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_91_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A2 a_700_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_91_48# A1 a_700_74# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A1 a_503_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND B1 a_91_48# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_700_74# A2 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_91_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

