* NGSPICE file created from sky130_fd_sc_ls__nor4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
M1000 Y C VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=8.594e+11p ps=6.85e+06u
M1001 Y a_57_368# a_446_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=4.648e+11p pd=3.07e+06u as=4.704e+11p ps=3.08e+06u
M1002 a_344_368# B a_260_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=4.032e+11p pd=2.96e+06u as=3.024e+11p ps=2.78e+06u
M1003 a_446_368# C a_344_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_57_368# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND B Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_260_368# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=4.354e+11p ps=3.08e+06u
M1007 VGND D_N a_57_368# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1008 VPWR D_N a_57_368# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1009 Y A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

