* File: sky130_fd_sc_ls__decap_8.pxi.spice
* Created: Fri Aug 28 13:11:43 2020
* 
x_PM_SKY130_FD_SC_LS__DECAP_8%VGND N_VGND_M1000_s N_VGND_M1002_g N_VGND_M1003_g
+ N_VGND_c_34_n N_VGND_c_35_n N_VGND_c_36_n N_VGND_c_37_n N_VGND_c_38_n
+ N_VGND_c_39_n N_VGND_c_40_n N_VGND_c_70_p N_VGND_c_41_n N_VGND_c_42_n
+ N_VGND_c_72_p VGND N_VGND_c_43_n N_VGND_c_44_n N_VGND_c_45_n N_VGND_c_46_n
+ N_VGND_c_47_n N_VGND_c_48_n PM_SKY130_FD_SC_LS__DECAP_8%VGND
x_PM_SKY130_FD_SC_LS__DECAP_8%VPWR N_VPWR_M1002_s N_VPWR_c_83_n N_VPWR_c_80_n
+ N_VPWR_c_81_n N_VPWR_c_85_n N_VPWR_c_86_n VPWR N_VPWR_M1000_g N_VPWR_M1001_g
+ N_VPWR_c_87_n N_VPWR_c_88_n N_VPWR_c_89_n N_VPWR_c_82_n N_VPWR_c_91_n
+ N_VPWR_c_92_n N_VPWR_c_93_n PM_SKY130_FD_SC_LS__DECAP_8%VPWR
cc_1 VNB N_VGND_c_34_n 0.0111177f $X=-0.19 $Y=-0.245 $X2=0.847 $Y2=0.528
cc_2 VNB N_VGND_c_35_n 0.0103054f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.42
cc_3 VNB N_VGND_c_36_n 0.0472714f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.42
cc_4 VNB N_VGND_c_37_n 0.0026191f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=0.64
cc_5 VNB N_VGND_c_38_n 0.0111278f $X=-0.19 $Y=-0.245 $X2=2.98 $Y2=0.5
cc_6 VNB N_VGND_c_39_n 0.0214492f $X=-0.19 $Y=-0.245 $X2=2.91 $Y2=1.42
cc_7 VNB N_VGND_c_40_n 0.0457426f $X=-0.19 $Y=-0.245 $X2=2.91 $Y2=1.42
cc_8 VNB N_VGND_c_41_n 0.0197615f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0
cc_9 VNB N_VGND_c_42_n 0.0059813f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=0
cc_10 VNB N_VGND_c_43_n 0.0201227f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0
cc_11 VNB N_VGND_c_44_n 0.0178522f $X=-0.19 $Y=-0.245 $X2=2.67 $Y2=0
cc_12 VNB N_VGND_c_45_n 0.0196454f $X=-0.19 $Y=-0.245 $X2=3.6 $Y2=0
cc_13 VNB N_VGND_c_46_n 0.245687f $X=-0.19 $Y=-0.245 $X2=3.6 $Y2=0
cc_14 VNB N_VGND_c_47_n 0.0102906f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0
cc_15 VNB N_VGND_c_48_n 0.0112875f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=0
cc_16 VNB N_VPWR_c_80_n 0.00204928f $X=-0.19 $Y=-0.245 $X2=2.575 $Y2=2.46
cc_17 VNB N_VPWR_c_81_n 0.326439f $X=-0.19 $Y=-0.245 $X2=2.575 $Y2=2.46
cc_18 VNB N_VPWR_c_82_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.42
cc_19 VPB N_VGND_M1002_g 0.0960913f $X=-0.19 $Y=1.66 $X2=1.3 $Y2=2.46
cc_20 VPB N_VGND_M1003_g 0.0949548f $X=-0.19 $Y=1.66 $X2=2.575 $Y2=2.46
cc_21 VPB N_VGND_c_36_n 0.0191045f $X=-0.19 $Y=1.66 $X2=0.965 $Y2=1.42
cc_22 VPB N_VGND_c_40_n 0.0191739f $X=-0.19 $Y=1.66 $X2=2.91 $Y2=1.42
cc_23 VPB N_VPWR_c_83_n 0.00851514f $X=-0.19 $Y=1.66 $X2=1.3 $Y2=2.46
cc_24 VPB N_VPWR_c_80_n 0.00727663f $X=-0.19 $Y=1.66 $X2=2.575 $Y2=2.46
cc_25 VPB N_VPWR_c_85_n 0.0204638f $X=-0.19 $Y=1.66 $X2=0.965 $Y2=1.42
cc_26 VPB N_VPWR_c_86_n 0.00842162f $X=-0.19 $Y=1.66 $X2=1.93 $Y2=0.085
cc_27 VPB N_VPWR_c_87_n 0.0201227f $X=-0.19 $Y=1.66 $X2=2.91 $Y2=1.42
cc_28 VPB N_VPWR_c_88_n 0.0201455f $X=-0.19 $Y=1.66 $X2=2.095 $Y2=0
cc_29 VPB N_VPWR_c_89_n 0.0193272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_82_n 0.0815913f $X=-0.19 $Y=1.66 $X2=0.965 $Y2=1.42
cc_31 VPB N_VPWR_c_91_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_92_n 0.017094f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0
cc_33 VPB N_VPWR_c_93_n 0.00459324f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=0
cc_34 N_VGND_M1002_g N_VPWR_c_83_n 0.026778f $X=1.3 $Y=2.46 $X2=0 $Y2=0
cc_35 N_VGND_M1002_g N_VPWR_c_80_n 0.0988648f $X=1.3 $Y=2.46 $X2=0 $Y2=0
cc_36 N_VGND_M1003_g N_VPWR_c_80_n 0.097201f $X=2.575 $Y=2.46 $X2=0 $Y2=0
cc_37 N_VGND_c_35_n N_VPWR_c_80_n 0.0156896f $X=0.965 $Y=1.42 $X2=0 $Y2=0
cc_38 N_VGND_c_36_n N_VPWR_c_80_n 0.010579f $X=0.965 $Y=1.42 $X2=0 $Y2=0
cc_39 N_VGND_c_37_n N_VPWR_c_80_n 0.0108665f $X=1.93 $Y=0.64 $X2=0 $Y2=0
cc_40 N_VGND_c_39_n N_VPWR_c_80_n 0.0198789f $X=2.91 $Y=1.42 $X2=0 $Y2=0
cc_41 N_VGND_c_40_n N_VPWR_c_80_n 0.00936628f $X=2.91 $Y=1.42 $X2=0 $Y2=0
cc_42 N_VGND_M1002_g N_VPWR_c_81_n 0.0179422f $X=1.3 $Y=2.46 $X2=0 $Y2=0
cc_43 N_VGND_M1003_g N_VPWR_c_81_n 0.0168878f $X=2.575 $Y=2.46 $X2=0 $Y2=0
cc_44 N_VGND_c_34_n N_VPWR_c_81_n 0.0281714f $X=0.847 $Y=0.528 $X2=0 $Y2=0
cc_45 N_VGND_c_35_n N_VPWR_c_81_n 0.0391218f $X=0.965 $Y=1.42 $X2=0 $Y2=0
cc_46 N_VGND_c_36_n N_VPWR_c_81_n 0.0337139f $X=0.965 $Y=1.42 $X2=0 $Y2=0
cc_47 N_VGND_c_37_n N_VPWR_c_81_n 0.0425313f $X=1.93 $Y=0.64 $X2=0 $Y2=0
cc_48 N_VGND_c_38_n N_VPWR_c_81_n 0.0286001f $X=2.98 $Y=0.5 $X2=0 $Y2=0
cc_49 N_VGND_c_39_n N_VPWR_c_81_n 0.0377586f $X=2.91 $Y=1.42 $X2=0 $Y2=0
cc_50 N_VGND_c_40_n N_VPWR_c_81_n 0.032126f $X=2.91 $Y=1.42 $X2=0 $Y2=0
cc_51 N_VGND_c_70_p N_VPWR_c_81_n 0.0172776f $X=0.65 $Y=0.64 $X2=0 $Y2=0
cc_52 N_VGND_c_41_n N_VPWR_c_81_n 0.0196799f $X=1.765 $Y=0 $X2=0 $Y2=0
cc_53 N_VGND_c_72_p N_VPWR_c_81_n 0.0196629f $X=3.205 $Y=0.64 $X2=0 $Y2=0
cc_54 N_VGND_c_44_n N_VPWR_c_81_n 0.0178177f $X=2.67 $Y=0 $X2=0 $Y2=0
cc_55 N_VGND_c_46_n N_VPWR_c_81_n 0.0731019f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_56 N_VGND_M1003_g N_VPWR_c_85_n 0.0201226f $X=2.575 $Y=2.46 $X2=0 $Y2=0
cc_57 N_VGND_M1003_g N_VPWR_c_86_n 0.028128f $X=2.575 $Y=2.46 $X2=0 $Y2=0
cc_58 N_VGND_M1002_g N_VPWR_c_88_n 0.0198149f $X=1.3 $Y=2.46 $X2=0 $Y2=0
cc_59 N_VGND_M1002_g N_VPWR_c_82_n 0.0388855f $X=1.3 $Y=2.46 $X2=0 $Y2=0
cc_60 N_VGND_M1003_g N_VPWR_c_82_n 0.0394876f $X=2.575 $Y=2.46 $X2=0 $Y2=0
