# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ls__nand4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__nand4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.735000 1.350000 8.085000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 6.160000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 4.195000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 2.275000 1.780000 ;
    END
  END D
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 8.640000 0.245000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 8.830000 3.520000 ;
    END
  END VPB
  PIN Y
    ANTENNADIFFAREA  3.321600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.820000 1.950000 8.515000 2.120000 ;
        RECT 1.820000 2.120000 2.150000 2.980000 ;
        RECT 2.820000 2.120000 3.430000 2.980000 ;
        RECT 4.670000 2.120000 5.280000 2.980000 ;
        RECT 6.745000 0.880000 8.515000 1.130000 ;
        RECT 6.815000 0.800000 7.005000 0.880000 ;
        RECT 7.320000 2.120000 8.010000 2.980000 ;
        RECT 7.755000 0.800000 7.945000 0.880000 ;
        RECT 8.285000 1.130000 8.515000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 2.575000 1.180000 ;
      RECT 0.115000  1.950000 1.650000 3.245000 ;
      RECT 0.615000  0.085000 0.945000 0.840000 ;
      RECT 1.115000  0.350000 1.445000 1.010000 ;
      RECT 1.615000  0.085000 1.945000 0.840000 ;
      RECT 2.245000  0.350000 4.365000 0.680000 ;
      RECT 2.245000  0.680000 2.575000 1.010000 ;
      RECT 2.320000  2.290000 2.650000 3.245000 ;
      RECT 2.745000  0.850000 3.935000 0.880000 ;
      RECT 2.745000  0.880000 6.215000 1.130000 ;
      RECT 3.600000  2.290000 4.500000 3.245000 ;
      RECT 4.595000  0.350000 8.525000 0.520000 ;
      RECT 4.595000  0.520000 4.925000 0.710000 ;
      RECT 5.095000  0.800000 5.285000 0.880000 ;
      RECT 5.450000  2.290000 7.140000 3.245000 ;
      RECT 5.455000  0.520000 5.785000 0.710000 ;
      RECT 5.955000  0.800000 6.145000 0.880000 ;
      RECT 6.315000  0.520000 6.645000 0.710000 ;
      RECT 7.175000  0.520000 7.505000 0.710000 ;
      RECT 8.190000  2.290000 8.520000 3.245000 ;
      RECT 8.195000  0.520000 8.525000 0.710000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_ls__nand4_4
END LIBRARY
