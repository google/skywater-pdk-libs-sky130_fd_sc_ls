* File: sky130_fd_sc_ls__inv_16.pxi.spice
* Created: Fri Aug 28 13:27:55 2020
* 
x_PM_SKY130_FD_SC_LS__INV_16%A N_A_c_161_n N_A_M1000_g N_A_M1002_g N_A_c_162_n
+ N_A_M1001_g N_A_M1003_g N_A_c_163_n N_A_M1004_g N_A_M1005_g N_A_c_164_n
+ N_A_M1006_g N_A_M1008_g N_A_c_165_n N_A_M1007_g N_A_M1009_g N_A_M1011_g
+ N_A_c_166_n N_A_M1010_g N_A_M1012_g N_A_c_167_n N_A_M1016_g N_A_M1013_g
+ N_A_c_168_n N_A_M1017_g N_A_M1014_g N_A_c_169_n N_A_M1020_g N_A_M1015_g
+ N_A_c_170_n N_A_M1021_g N_A_M1018_g N_A_c_171_n N_A_M1022_g N_A_M1019_g
+ N_A_c_172_n N_A_M1024_g N_A_M1023_g N_A_c_173_n N_A_M1025_g N_A_M1027_g
+ N_A_c_174_n N_A_M1026_g N_A_M1029_g N_A_c_175_n N_A_M1028_g N_A_M1031_g
+ N_A_c_176_n N_A_M1030_g N_A_c_151_n N_A_c_152_n A N_A_c_153_n N_A_c_154_n
+ N_A_c_155_n N_A_c_156_n N_A_c_157_n N_A_c_158_n N_A_c_159_n N_A_c_160_n
+ N_A_c_187_n A PM_SKY130_FD_SC_LS__INV_16%A
x_PM_SKY130_FD_SC_LS__INV_16%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_M1006_d
+ N_VPWR_M1010_d N_VPWR_M1017_d N_VPWR_M1021_d N_VPWR_M1024_d N_VPWR_M1026_d
+ N_VPWR_M1030_d N_VPWR_c_468_n N_VPWR_c_469_n N_VPWR_c_470_n N_VPWR_c_471_n
+ N_VPWR_c_472_n N_VPWR_c_473_n N_VPWR_c_474_n N_VPWR_c_475_n N_VPWR_c_476_n
+ N_VPWR_c_477_n N_VPWR_c_478_n N_VPWR_c_479_n N_VPWR_c_480_n N_VPWR_c_481_n
+ N_VPWR_c_482_n VPWR N_VPWR_c_483_n N_VPWR_c_484_n N_VPWR_c_485_n
+ N_VPWR_c_486_n N_VPWR_c_487_n N_VPWR_c_488_n N_VPWR_c_489_n N_VPWR_c_490_n
+ N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_467_n
+ PM_SKY130_FD_SC_LS__INV_16%VPWR
x_PM_SKY130_FD_SC_LS__INV_16%Y N_Y_M1002_d N_Y_M1005_d N_Y_M1009_d N_Y_M1012_d
+ N_Y_M1014_d N_Y_M1018_d N_Y_M1023_d N_Y_M1029_d N_Y_M1000_s N_Y_M1004_s
+ N_Y_M1007_s N_Y_M1016_s N_Y_M1020_s N_Y_M1022_s N_Y_M1025_s N_Y_M1028_s
+ N_Y_c_613_n N_Y_c_627_n N_Y_c_614_n N_Y_c_629_n N_Y_c_615_n N_Y_c_616_n
+ N_Y_c_632_n N_Y_c_617_n N_Y_c_618_n N_Y_c_619_n N_Y_c_620_n N_Y_c_621_n
+ N_Y_c_695_n N_Y_c_622_n N_Y_c_623_n N_Y_c_624_n Y N_Y_c_633_n N_Y_c_625_n
+ N_Y_c_635_n N_Y_c_636_n N_Y_c_626_n N_Y_c_741_n N_Y_c_765_n N_Y_c_769_n
+ N_Y_c_772_n PM_SKY130_FD_SC_LS__INV_16%Y
x_PM_SKY130_FD_SC_LS__INV_16%VGND N_VGND_M1002_s N_VGND_M1003_s N_VGND_M1008_s
+ N_VGND_M1011_s N_VGND_M1013_s N_VGND_M1015_s N_VGND_M1019_s N_VGND_M1027_s
+ N_VGND_M1031_s N_VGND_c_858_n N_VGND_c_859_n N_VGND_c_860_n N_VGND_c_861_n
+ N_VGND_c_862_n N_VGND_c_863_n N_VGND_c_864_n N_VGND_c_865_n N_VGND_c_866_n
+ N_VGND_c_867_n N_VGND_c_868_n N_VGND_c_869_n N_VGND_c_870_n N_VGND_c_871_n
+ N_VGND_c_872_n N_VGND_c_873_n N_VGND_c_874_n VGND N_VGND_c_875_n
+ N_VGND_c_876_n N_VGND_c_877_n N_VGND_c_878_n N_VGND_c_879_n N_VGND_c_880_n
+ N_VGND_c_881_n N_VGND_c_882_n N_VGND_c_883_n N_VGND_c_884_n
+ PM_SKY130_FD_SC_LS__INV_16%VGND
cc_1 VNB N_A_M1002_g 0.0298158f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_2 VNB N_A_M1003_g 0.0244831f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_A_M1005_g 0.0236443f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.74
cc_4 VNB N_A_M1008_g 0.0246673f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_5 VNB N_A_M1009_g 0.0236422f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=0.74
cc_6 VNB N_A_M1011_g 0.0236401f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=0.74
cc_7 VNB N_A_M1012_g 0.023639f $X=-0.19 $Y=-0.245 $X2=3.355 $Y2=0.74
cc_8 VNB N_A_M1013_g 0.0236474f $X=-0.19 $Y=-0.245 $X2=3.785 $Y2=0.74
cc_9 VNB N_A_M1014_g 0.0230083f $X=-0.19 $Y=-0.245 $X2=4.215 $Y2=0.74
cc_10 VNB N_A_M1015_g 0.0236404f $X=-0.19 $Y=-0.245 $X2=4.645 $Y2=0.74
cc_11 VNB N_A_M1018_g 0.024294f $X=-0.19 $Y=-0.245 $X2=5.145 $Y2=0.74
cc_12 VNB N_A_M1019_g 0.0245364f $X=-0.19 $Y=-0.245 $X2=5.575 $Y2=0.74
cc_13 VNB N_A_M1023_g 0.0251803f $X=-0.19 $Y=-0.245 $X2=6.145 $Y2=0.74
cc_14 VNB N_A_M1027_g 0.0247749f $X=-0.19 $Y=-0.245 $X2=6.575 $Y2=0.74
cc_15 VNB N_A_M1029_g 0.0256095f $X=-0.19 $Y=-0.245 $X2=7.165 $Y2=0.74
cc_16 VNB N_A_M1031_g 0.0298291f $X=-0.19 $Y=-0.245 $X2=7.595 $Y2=0.74
cc_17 VNB N_A_c_151_n 0.0184543f $X=-0.19 $Y=-0.245 $X2=7.09 $Y2=1.515
cc_18 VNB N_A_c_152_n 0.0448453f $X=-0.19 $Y=-0.245 $X2=7.595 $Y2=1.557
cc_19 VNB N_A_c_153_n 0.277938f $X=-0.19 $Y=-0.245 $X2=6.745 $Y2=1.515
cc_20 VNB N_A_c_154_n 0.0023355f $X=-0.19 $Y=-0.245 $X2=6.925 $Y2=1.515
cc_21 VNB N_A_c_155_n 0.00173377f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.515
cc_22 VNB N_A_c_156_n 0.00173377f $X=-0.19 $Y=-0.245 $X2=2.17 $Y2=1.515
cc_23 VNB N_A_c_157_n 0.00173377f $X=-0.19 $Y=-0.245 $X2=3.11 $Y2=1.515
cc_24 VNB N_A_c_158_n 0.00101987f $X=-0.19 $Y=-0.245 $X2=4.025 $Y2=1.515
cc_25 VNB N_A_c_159_n 0.00173377f $X=-0.19 $Y=-0.245 $X2=4.935 $Y2=1.515
cc_26 VNB N_A_c_160_n 0.0022845f $X=-0.19 $Y=-0.245 $X2=5.93 $Y2=1.515
cc_27 VNB N_VPWR_c_467_n 0.342803f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.557
cc_28 VNB N_Y_c_613_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=3.785 $Y2=0.74
cc_29 VNB N_Y_c_614_n 0.00468918f $X=-0.19 $Y=-0.245 $X2=4.255 $Y2=1.765
cc_30 VNB N_Y_c_615_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=4.705 $Y2=2.4
cc_31 VNB N_Y_c_616_n 0.00417093f $X=-0.19 $Y=-0.245 $X2=5.145 $Y2=0.74
cc_32 VNB N_Y_c_617_n 0.00219079f $X=-0.19 $Y=-0.245 $X2=5.575 $Y2=0.74
cc_33 VNB N_Y_c_618_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_619_n 0.00237467f $X=-0.19 $Y=-0.245 $X2=5.655 $Y2=2.4
cc_35 VNB N_Y_c_620_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=6.145 $Y2=1.35
cc_36 VNB N_Y_c_621_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=6.205 $Y2=1.765
cc_37 VNB N_Y_c_622_n 0.00169784f $X=-0.19 $Y=-0.245 $X2=6.575 $Y2=1.35
cc_38 VNB N_Y_c_623_n 0.00142546f $X=-0.19 $Y=-0.245 $X2=6.575 $Y2=0.74
cc_39 VNB N_Y_c_624_n 0.00101819f $X=-0.19 $Y=-0.245 $X2=6.655 $Y2=2.4
cc_40 VNB N_Y_c_625_n 0.00473182f $X=-0.19 $Y=-0.245 $X2=7.595 $Y2=0.74
cc_41 VNB N_Y_c_626_n 0.00203504f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.557
cc_42 VNB N_VGND_c_858_n 0.0131032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_859_n 0.0502481f $X=-0.19 $Y=-0.245 $X2=2.405 $Y2=2.4
cc_44 VNB N_VGND_c_860_n 0.00986225f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=0.74
cc_45 VNB N_VGND_c_861_n 0.0103371f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=0.74
cc_46 VNB N_VGND_c_862_n 0.0100559f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=2.4
cc_47 VNB N_VGND_c_863_n 0.00669123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_864_n 0.0105034f $X=-0.19 $Y=-0.245 $X2=3.785 $Y2=1.35
cc_49 VNB N_VGND_c_865_n 0.012516f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.765
cc_50 VNB N_VGND_c_866_n 0.0121504f $X=-0.19 $Y=-0.245 $X2=4.215 $Y2=0.74
cc_51 VNB N_VGND_c_867_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_868_n 0.0567567f $X=-0.19 $Y=-0.245 $X2=4.255 $Y2=2.4
cc_53 VNB N_VGND_c_869_n 0.0181599f $X=-0.19 $Y=-0.245 $X2=4.645 $Y2=0.74
cc_54 VNB N_VGND_c_870_n 0.00482535f $X=-0.19 $Y=-0.245 $X2=4.645 $Y2=0.74
cc_55 VNB N_VGND_c_871_n 0.0173725f $X=-0.19 $Y=-0.245 $X2=4.705 $Y2=1.765
cc_56 VNB N_VGND_c_872_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=4.705 $Y2=2.4
cc_57 VNB N_VGND_c_873_n 0.0191493f $X=-0.19 $Y=-0.245 $X2=5.145 $Y2=1.35
cc_58 VNB N_VGND_c_874_n 0.00615512f $X=-0.19 $Y=-0.245 $X2=5.145 $Y2=0.74
cc_59 VNB N_VGND_c_875_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=5.175 $Y2=1.765
cc_60 VNB N_VGND_c_876_n 0.0183708f $X=-0.19 $Y=-0.245 $X2=5.575 $Y2=0.74
cc_61 VNB N_VGND_c_877_n 0.018851f $X=-0.19 $Y=-0.245 $X2=6.145 $Y2=1.35
cc_62 VNB N_VGND_c_878_n 0.019013f $X=-0.19 $Y=-0.245 $X2=7.165 $Y2=0.74
cc_63 VNB N_VGND_c_879_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=7.205 $Y2=2.4
cc_64 VNB N_VGND_c_880_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=7.09 $Y2=1.515
cc_65 VNB N_VGND_c_881_n 0.00538573f $X=-0.19 $Y=-0.245 $X2=7.595 $Y2=1.557
cc_66 VNB N_VGND_c_882_n 0.00519339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_883_n 0.00653982f $X=-0.19 $Y=-0.245 $X2=6.925 $Y2=1.515
cc_68 VNB N_VGND_c_884_n 0.436313f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.557
cc_69 VPB N_A_c_161_n 0.0173152f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_70 VPB N_A_c_162_n 0.0155292f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_71 VPB N_A_c_163_n 0.0157376f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_72 VPB N_A_c_164_n 0.0154932f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.765
cc_73 VPB N_A_c_165_n 0.0157372f $X=-0.19 $Y=1.66 $X2=2.405 $Y2=1.765
cc_74 VPB N_A_c_166_n 0.0154926f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=1.765
cc_75 VPB N_A_c_167_n 0.0154907f $X=-0.19 $Y=1.66 $X2=3.355 $Y2=1.765
cc_76 VPB N_A_c_168_n 0.0154576f $X=-0.19 $Y=1.66 $X2=3.805 $Y2=1.765
cc_77 VPB N_A_c_169_n 0.0154574f $X=-0.19 $Y=1.66 $X2=4.255 $Y2=1.765
cc_78 VPB N_A_c_170_n 0.0155916f $X=-0.19 $Y=1.66 $X2=4.705 $Y2=1.765
cc_79 VPB N_A_c_171_n 0.0158394f $X=-0.19 $Y=1.66 $X2=5.175 $Y2=1.765
cc_80 VPB N_A_c_172_n 0.0163606f $X=-0.19 $Y=1.66 $X2=5.655 $Y2=1.765
cc_81 VPB N_A_c_173_n 0.0158334f $X=-0.19 $Y=1.66 $X2=6.205 $Y2=1.765
cc_82 VPB N_A_c_174_n 0.0158329f $X=-0.19 $Y=1.66 $X2=6.655 $Y2=1.765
cc_83 VPB N_A_c_175_n 0.0159293f $X=-0.19 $Y=1.66 $X2=7.205 $Y2=1.765
cc_84 VPB N_A_c_176_n 0.017726f $X=-0.19 $Y=1.66 $X2=7.655 $Y2=1.765
cc_85 VPB N_A_c_151_n 0.0106624f $X=-0.19 $Y=1.66 $X2=7.09 $Y2=1.515
cc_86 VPB N_A_c_152_n 0.0250468f $X=-0.19 $Y=1.66 $X2=7.595 $Y2=1.557
cc_87 VPB N_A_c_153_n 0.196749f $X=-0.19 $Y=1.66 $X2=6.745 $Y2=1.515
cc_88 VPB N_A_c_154_n 0.00200166f $X=-0.19 $Y=1.66 $X2=6.925 $Y2=1.515
cc_89 VPB N_A_c_155_n 0.00198992f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.515
cc_90 VPB N_A_c_156_n 0.00198947f $X=-0.19 $Y=1.66 $X2=2.17 $Y2=1.515
cc_91 VPB N_A_c_157_n 0.00178763f $X=-0.19 $Y=1.66 $X2=3.11 $Y2=1.515
cc_92 VPB N_A_c_158_n 0.00170434f $X=-0.19 $Y=1.66 $X2=4.025 $Y2=1.515
cc_93 VPB N_A_c_159_n 0.00165017f $X=-0.19 $Y=1.66 $X2=4.935 $Y2=1.515
cc_94 VPB N_A_c_160_n 0.00185727f $X=-0.19 $Y=1.66 $X2=5.93 $Y2=1.515
cc_95 VPB N_A_c_187_n 0.0106995f $X=-0.19 $Y=1.66 $X2=6.925 $Y2=1.665
cc_96 VPB N_VPWR_c_468_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_469_n 0.0645244f $X=-0.19 $Y=1.66 $X2=2.405 $Y2=2.4
cc_98 VPB N_VPWR_c_470_n 0.00918066f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=1.35
cc_99 VPB N_VPWR_c_471_n 0.00886117f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=2.4
cc_100 VPB N_VPWR_c_472_n 0.0082016f $X=-0.19 $Y=1.66 $X2=3.355 $Y2=2.4
cc_101 VPB N_VPWR_c_473_n 0.00741433f $X=-0.19 $Y=1.66 $X2=3.805 $Y2=1.765
cc_102 VPB N_VPWR_c_474_n 0.00792857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_475_n 0.00836621f $X=-0.19 $Y=1.66 $X2=4.645 $Y2=0.74
cc_104 VPB N_VPWR_c_476_n 0.00824869f $X=-0.19 $Y=1.66 $X2=5.145 $Y2=0.74
cc_105 VPB N_VPWR_c_477_n 0.0118062f $X=-0.19 $Y=1.66 $X2=5.175 $Y2=2.4
cc_106 VPB N_VPWR_c_478_n 0.0679009f $X=-0.19 $Y=1.66 $X2=5.575 $Y2=1.35
cc_107 VPB N_VPWR_c_479_n 0.0189682f $X=-0.19 $Y=1.66 $X2=5.655 $Y2=2.4
cc_108 VPB N_VPWR_c_480_n 0.00449427f $X=-0.19 $Y=1.66 $X2=5.655 $Y2=2.4
cc_109 VPB N_VPWR_c_481_n 0.0186762f $X=-0.19 $Y=1.66 $X2=6.145 $Y2=0.74
cc_110 VPB N_VPWR_c_482_n 0.00545601f $X=-0.19 $Y=1.66 $X2=6.145 $Y2=0.74
cc_111 VPB N_VPWR_c_483_n 0.0193162f $X=-0.19 $Y=1.66 $X2=6.205 $Y2=2.4
cc_112 VPB N_VPWR_c_484_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_485_n 0.0196495f $X=-0.19 $Y=1.66 $X2=7.165 $Y2=0.74
cc_114 VPB N_VPWR_c_486_n 0.0187479f $X=-0.19 $Y=1.66 $X2=7.655 $Y2=2.4
cc_115 VPB N_VPWR_c_487_n 0.0186948f $X=-0.19 $Y=1.66 $X2=7.595 $Y2=1.557
cc_116 VPB N_VPWR_c_488_n 0.0180795f $X=-0.19 $Y=1.66 $X2=6.925 $Y2=1.515
cc_117 VPB N_VPWR_c_489_n 0.00555219f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.515
cc_118 VPB N_VPWR_c_490_n 0.0047828f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.557
cc_119 VPB N_VPWR_c_491_n 0.0047828f $X=-0.19 $Y=1.66 $X2=2.17 $Y2=1.515
cc_120 VPB N_VPWR_c_492_n 0.00632158f $X=-0.19 $Y=1.66 $X2=2.425 $Y2=1.557
cc_121 VPB N_VPWR_c_493_n 0.00632158f $X=-0.19 $Y=1.66 $X2=3.11 $Y2=1.515
cc_122 VPB N_VPWR_c_467_n 0.0896775f $X=-0.19 $Y=1.66 $X2=3.805 $Y2=1.557
cc_123 VPB N_Y_c_627_n 0.00257348f $X=-0.19 $Y=1.66 $X2=4.215 $Y2=1.35
cc_124 VPB N_Y_c_614_n 9.14603e-19 $X=-0.19 $Y=1.66 $X2=4.255 $Y2=1.765
cc_125 VPB N_Y_c_629_n 0.00257348f $X=-0.19 $Y=1.66 $X2=4.645 $Y2=0.74
cc_126 VPB N_Y_c_615_n 6.01664e-19 $X=-0.19 $Y=1.66 $X2=4.705 $Y2=2.4
cc_127 VPB N_Y_c_616_n 0.001512f $X=-0.19 $Y=1.66 $X2=5.145 $Y2=0.74
cc_128 VPB N_Y_c_632_n 0.00290642f $X=-0.19 $Y=1.66 $X2=5.175 $Y2=2.4
cc_129 VPB N_Y_c_633_n 0.00250852f $X=-0.19 $Y=1.66 $X2=7.165 $Y2=0.74
cc_130 VPB N_Y_c_625_n 0.00347841f $X=-0.19 $Y=1.66 $X2=7.595 $Y2=0.74
cc_131 VPB N_Y_c_635_n 0.00477967f $X=-0.19 $Y=1.66 $X2=1.085 $Y2=1.55
cc_132 VPB N_Y_c_636_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.557
cc_133 VPB N_Y_c_626_n 0.00389939f $X=-0.19 $Y=1.66 $X2=1.495 $Y2=1.557
cc_134 N_A_c_161_n N_VPWR_c_469_n 0.00982454f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A_c_162_n N_VPWR_c_470_n 0.00326696f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A_c_163_n N_VPWR_c_470_n 0.00879365f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A_c_153_n N_VPWR_c_470_n 0.00186112f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A_c_155_n N_VPWR_c_470_n 0.0191349f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_139 N_A_c_187_n N_VPWR_c_470_n 8.28135e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_140 N_A_c_164_n N_VPWR_c_471_n 0.00641233f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A_c_165_n N_VPWR_c_471_n 0.00870475f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A_c_153_n N_VPWR_c_471_n 0.00130763f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_143 N_A_c_156_n N_VPWR_c_471_n 0.0176185f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_144 N_A_c_187_n N_VPWR_c_471_n 7.92963e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_145 N_A_c_166_n N_VPWR_c_472_n 0.00641233f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A_c_167_n N_VPWR_c_472_n 0.00740094f $X=3.355 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A_c_153_n N_VPWR_c_472_n 0.00130763f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_148 N_A_c_157_n N_VPWR_c_472_n 0.0176185f $X=3.11 $Y=1.515 $X2=0 $Y2=0
cc_149 N_A_c_187_n N_VPWR_c_472_n 7.92963e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_150 N_A_c_168_n N_VPWR_c_473_n 0.00207454f $X=3.805 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A_c_169_n N_VPWR_c_473_n 0.00205852f $X=4.255 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A_c_153_n N_VPWR_c_473_n 0.00120219f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_153 N_A_c_158_n N_VPWR_c_473_n 0.016086f $X=4.025 $Y=1.515 $X2=0 $Y2=0
cc_154 N_A_c_187_n N_VPWR_c_473_n 7.45001e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_155 N_A_c_170_n N_VPWR_c_474_n 0.00213354f $X=4.705 $Y=1.765 $X2=0 $Y2=0
cc_156 N_A_c_171_n N_VPWR_c_474_n 0.00224365f $X=5.175 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A_c_153_n N_VPWR_c_474_n 0.00162144f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_158 N_A_c_159_n N_VPWR_c_474_n 0.0186433f $X=4.935 $Y=1.515 $X2=0 $Y2=0
cc_159 N_A_c_187_n N_VPWR_c_474_n 9.45027e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_160 N_A_c_172_n N_VPWR_c_475_n 0.00822207f $X=5.655 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A_c_173_n N_VPWR_c_475_n 0.00819414f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A_c_153_n N_VPWR_c_475_n 0.00179937f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_163 N_A_c_160_n N_VPWR_c_475_n 0.0227815f $X=5.93 $Y=1.515 $X2=0 $Y2=0
cc_164 N_A_c_187_n N_VPWR_c_475_n 0.00106883f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_165 N_A_c_174_n N_VPWR_c_476_n 0.00819414f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A_c_175_n N_VPWR_c_476_n 0.00815589f $X=7.205 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A_c_151_n N_VPWR_c_476_n 0.00177166f $X=7.09 $Y=1.515 $X2=0 $Y2=0
cc_168 N_A_c_154_n N_VPWR_c_476_n 0.0224748f $X=6.925 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A_c_187_n N_VPWR_c_476_n 9.92096e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_170 N_A_c_176_n N_VPWR_c_478_n 0.0053639f $X=7.655 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A_c_152_n N_VPWR_c_478_n 4.64517e-19 $X=7.595 $Y=1.557 $X2=0 $Y2=0
cc_172 N_A_c_167_n N_VPWR_c_479_n 0.00445602f $X=3.355 $Y=1.765 $X2=0 $Y2=0
cc_173 N_A_c_168_n N_VPWR_c_479_n 0.00461464f $X=3.805 $Y=1.765 $X2=0 $Y2=0
cc_174 N_A_c_169_n N_VPWR_c_481_n 0.00461464f $X=4.255 $Y=1.765 $X2=0 $Y2=0
cc_175 N_A_c_170_n N_VPWR_c_481_n 0.00461464f $X=4.705 $Y=1.765 $X2=0 $Y2=0
cc_176 N_A_c_161_n N_VPWR_c_483_n 0.00445411f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A_c_162_n N_VPWR_c_483_n 0.00456878f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A_c_163_n N_VPWR_c_484_n 0.00445602f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_179 N_A_c_164_n N_VPWR_c_484_n 0.00445602f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A_c_165_n N_VPWR_c_485_n 0.00445602f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_181 N_A_c_166_n N_VPWR_c_485_n 0.00445602f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A_c_171_n N_VPWR_c_486_n 0.00461464f $X=5.175 $Y=1.765 $X2=0 $Y2=0
cc_183 N_A_c_172_n N_VPWR_c_486_n 0.00461464f $X=5.655 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A_c_173_n N_VPWR_c_487_n 0.00445602f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_185 N_A_c_174_n N_VPWR_c_487_n 0.00445602f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A_c_175_n N_VPWR_c_488_n 0.00445602f $X=7.205 $Y=1.765 $X2=0 $Y2=0
cc_187 N_A_c_176_n N_VPWR_c_488_n 0.00461464f $X=7.655 $Y=1.765 $X2=0 $Y2=0
cc_188 N_A_c_161_n N_VPWR_c_467_n 0.00860947f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A_c_162_n N_VPWR_c_467_n 0.00890056f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A_c_163_n N_VPWR_c_467_n 0.00857378f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A_c_164_n N_VPWR_c_467_n 0.0085805f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A_c_165_n N_VPWR_c_467_n 0.00857378f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_193 N_A_c_166_n N_VPWR_c_467_n 0.0085805f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_194 N_A_c_167_n N_VPWR_c_467_n 0.00857378f $X=3.355 $Y=1.765 $X2=0 $Y2=0
cc_195 N_A_c_168_n N_VPWR_c_467_n 0.00908279f $X=3.805 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A_c_169_n N_VPWR_c_467_n 0.00908167f $X=4.255 $Y=1.765 $X2=0 $Y2=0
cc_197 N_A_c_170_n N_VPWR_c_467_n 0.00908357f $X=4.705 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A_c_171_n N_VPWR_c_467_n 0.00908078f $X=5.175 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A_c_172_n N_VPWR_c_467_n 0.00909441f $X=5.655 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A_c_173_n N_VPWR_c_467_n 0.00857797f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A_c_174_n N_VPWR_c_467_n 0.00857797f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A_c_175_n N_VPWR_c_467_n 0.00857797f $X=7.205 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A_c_176_n N_VPWR_c_467_n 0.00911101f $X=7.655 $Y=1.765 $X2=0 $Y2=0
cc_204 N_A_M1002_g N_Y_c_613_n 0.00772833f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A_M1003_g N_Y_c_613_n 0.00746162f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_c_163_n N_Y_c_627_n 0.00869437f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_207 N_A_c_164_n N_Y_c_627_n 0.00930243f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_208 N_A_M1003_g N_Y_c_614_n 8.65347e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A_c_163_n N_Y_c_614_n 0.0011501f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A_M1005_g N_Y_c_614_n 0.0151729f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A_c_164_n N_Y_c_614_n 0.00377504f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A_M1008_g N_Y_c_614_n 0.00396849f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A_c_165_n N_Y_c_614_n 8.76409e-19 $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_214 N_A_c_153_n N_Y_c_614_n 0.0280623f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_215 N_A_c_155_n N_Y_c_614_n 0.0286513f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_216 N_A_c_156_n N_Y_c_614_n 0.0285602f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_217 N_A_c_187_n N_Y_c_614_n 0.0319514f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_218 N_A_c_165_n N_Y_c_629_n 0.00920447f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A_c_166_n N_Y_c_629_n 0.00981252f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A_M1008_g N_Y_c_615_n 8.58503e-19 $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_c_165_n N_Y_c_615_n 0.00118452f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_222 N_A_M1009_g N_Y_c_615_n 0.015703f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A_M1011_g N_Y_c_615_n 0.0156374f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_c_166_n N_Y_c_615_n 0.00374802f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_225 N_A_M1012_g N_Y_c_615_n 8.54281e-19 $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A_c_167_n N_Y_c_615_n 8.72571e-19 $X=3.355 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A_c_153_n N_Y_c_615_n 0.0303703f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_228 N_A_c_156_n N_Y_c_615_n 0.0286513f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_229 N_A_c_157_n N_Y_c_615_n 0.0285726f $X=3.11 $Y=1.515 $X2=0 $Y2=0
cc_230 N_A_c_187_n N_Y_c_615_n 0.0337883f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_231 N_A_M1014_g N_Y_c_616_n 0.00354167f $X=4.215 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A_c_169_n N_Y_c_616_n 0.00187851f $X=4.255 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A_M1015_g N_Y_c_616_n 0.0154727f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A_c_170_n N_Y_c_616_n 0.00110542f $X=4.705 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A_M1018_g N_Y_c_616_n 8.71251e-19 $X=5.145 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A_c_153_n N_Y_c_616_n 0.0262298f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_237 N_A_c_158_n N_Y_c_616_n 0.0283819f $X=4.025 $Y=1.515 $X2=0 $Y2=0
cc_238 N_A_c_159_n N_Y_c_616_n 0.0284993f $X=4.935 $Y=1.515 $X2=0 $Y2=0
cc_239 N_A_c_187_n N_Y_c_616_n 0.0287175f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_240 N_A_c_170_n N_Y_c_632_n 4.16925e-19 $X=4.705 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A_M1018_g N_Y_c_617_n 0.00526964f $X=5.145 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A_M1019_g N_Y_c_617_n 0.0110561f $X=5.575 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A_M1023_g N_Y_c_617_n 9.81084e-19 $X=6.145 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_c_153_n N_Y_c_617_n 0.0078283f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_245 N_A_c_159_n N_Y_c_617_n 0.00658047f $X=4.935 $Y=1.515 $X2=0 $Y2=0
cc_246 N_A_c_160_n N_Y_c_617_n 0.00676348f $X=5.93 $Y=1.515 $X2=0 $Y2=0
cc_247 N_A_c_187_n N_Y_c_617_n 0.00205475f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_248 N_A_M1018_g N_Y_c_618_n 0.00722691f $X=5.145 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A_M1019_g N_Y_c_618_n 0.00830039f $X=5.575 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A_M1023_g N_Y_c_619_n 0.00815379f $X=6.145 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A_M1027_g N_Y_c_619_n 0.0120406f $X=6.575 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_M1029_g N_Y_c_619_n 9.51769e-19 $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_c_153_n N_Y_c_619_n 0.00842099f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_254 N_A_c_154_n N_Y_c_619_n 0.00735182f $X=6.925 $Y=1.515 $X2=0 $Y2=0
cc_255 N_A_c_160_n N_Y_c_619_n 0.00737762f $X=5.93 $Y=1.515 $X2=0 $Y2=0
cc_256 N_A_c_187_n N_Y_c_619_n 0.00280382f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_257 N_A_M1023_g N_Y_c_620_n 0.0080359f $X=6.145 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A_M1027_g N_Y_c_620_n 0.00821155f $X=6.575 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A_M1029_g N_Y_c_621_n 0.00753493f $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A_M1031_g N_Y_c_621_n 0.00772833f $X=7.595 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_M1002_g N_Y_c_695_n 0.00362234f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_c_153_n N_Y_c_695_n 0.0144997f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_263 N_A_c_155_n N_Y_c_695_n 0.0279825f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_264 N_A_M1002_g N_Y_c_622_n 0.0102796f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A_M1003_g N_Y_c_622_n 0.00319122f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_266 N_A_M1002_g N_Y_c_623_n 0.00198651f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A_M1003_g N_Y_c_623_n 0.0031608f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A_M1029_g N_Y_c_624_n 0.0031805f $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_M1031_g N_Y_c_624_n 0.00198651f $X=7.595 $Y=0.74 $X2=0 $Y2=0
cc_270 N_A_c_161_n N_Y_c_633_n 0.0169904f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_271 N_A_c_162_n N_Y_c_633_n 0.0136985f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_272 N_A_c_163_n N_Y_c_633_n 8.08789e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_273 N_A_c_153_n N_Y_c_633_n 0.0303512f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_274 N_A_c_187_n N_Y_c_633_n 0.00187673f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_275 N_A_M1011_g N_Y_c_625_n 8.44821e-19 $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A_c_166_n N_Y_c_625_n 7.72041e-19 $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_277 N_A_M1012_g N_Y_c_625_n 0.0148554f $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_278 N_A_c_167_n N_Y_c_625_n 0.0138412f $X=3.355 $Y=1.765 $X2=0 $Y2=0
cc_279 N_A_M1013_g N_Y_c_625_n 0.00398243f $X=3.785 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A_c_168_n N_Y_c_625_n 0.00189446f $X=3.805 $Y=1.765 $X2=0 $Y2=0
cc_281 N_A_c_153_n N_Y_c_625_n 0.0282849f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_282 N_A_c_157_n N_Y_c_625_n 0.0293067f $X=3.11 $Y=1.515 $X2=0 $Y2=0
cc_283 N_A_c_158_n N_Y_c_625_n 0.0285537f $X=4.025 $Y=1.515 $X2=0 $Y2=0
cc_284 N_A_c_187_n N_Y_c_625_n 0.0323804f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_285 N_A_c_171_n N_Y_c_635_n 0.00195892f $X=5.175 $Y=1.765 $X2=0 $Y2=0
cc_286 N_A_c_172_n N_Y_c_635_n 0.00247321f $X=5.655 $Y=1.765 $X2=0 $Y2=0
cc_287 N_A_c_153_n N_Y_c_635_n 0.0221324f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_288 N_A_c_159_n N_Y_c_635_n 0.021723f $X=4.935 $Y=1.515 $X2=0 $Y2=0
cc_289 N_A_c_160_n N_Y_c_635_n 0.0220842f $X=5.93 $Y=1.515 $X2=0 $Y2=0
cc_290 N_A_c_187_n N_Y_c_635_n 0.0341673f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_291 N_A_c_172_n N_Y_c_636_n 0.00109841f $X=5.655 $Y=1.765 $X2=0 $Y2=0
cc_292 N_A_c_173_n N_Y_c_636_n 0.0145129f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_293 N_A_c_174_n N_Y_c_636_n 0.0143565f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_294 N_A_c_175_n N_Y_c_636_n 8.03222e-19 $X=7.205 $Y=1.765 $X2=0 $Y2=0
cc_295 N_A_c_153_n N_Y_c_636_n 0.0227953f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_296 N_A_c_154_n N_Y_c_636_n 0.0214823f $X=6.925 $Y=1.515 $X2=0 $Y2=0
cc_297 N_A_c_160_n N_Y_c_636_n 0.0215141f $X=5.93 $Y=1.515 $X2=0 $Y2=0
cc_298 N_A_c_187_n N_Y_c_636_n 0.0351299f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_299 N_A_c_174_n N_Y_c_626_n 7.82206e-19 $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_300 N_A_M1029_g N_Y_c_626_n 0.0051716f $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_301 N_A_c_175_n N_Y_c_626_n 0.0140988f $X=7.205 $Y=1.765 $X2=0 $Y2=0
cc_302 N_A_M1031_g N_Y_c_626_n 0.0113953f $X=7.595 $Y=0.74 $X2=0 $Y2=0
cc_303 N_A_c_176_n N_Y_c_626_n 0.00238575f $X=7.655 $Y=1.765 $X2=0 $Y2=0
cc_304 N_A_c_152_n N_Y_c_626_n 0.0400179f $X=7.595 $Y=1.557 $X2=0 $Y2=0
cc_305 N_A_c_154_n N_Y_c_626_n 0.0291941f $X=6.925 $Y=1.515 $X2=0 $Y2=0
cc_306 N_A_c_187_n N_Y_c_626_n 0.00184883f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_307 N_A_c_162_n N_Y_c_741_n 0.0124768f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_308 N_A_c_163_n N_Y_c_741_n 0.00887184f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_309 N_A_c_164_n N_Y_c_741_n 0.00701605f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_310 N_A_c_165_n N_Y_c_741_n 0.00887184f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_311 N_A_c_166_n N_Y_c_741_n 0.00701605f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_312 N_A_c_167_n N_Y_c_741_n 0.00875751f $X=3.355 $Y=1.765 $X2=0 $Y2=0
cc_313 N_A_c_168_n N_Y_c_741_n 0.00774121f $X=3.805 $Y=1.765 $X2=0 $Y2=0
cc_314 N_A_c_169_n N_Y_c_741_n 0.00766908f $X=4.255 $Y=1.765 $X2=0 $Y2=0
cc_315 N_A_c_170_n N_Y_c_741_n 0.00764117f $X=4.705 $Y=1.765 $X2=0 $Y2=0
cc_316 N_A_c_171_n N_Y_c_741_n 0.00766908f $X=5.175 $Y=1.765 $X2=0 $Y2=0
cc_317 N_A_c_172_n N_Y_c_741_n 0.00962379f $X=5.655 $Y=1.765 $X2=0 $Y2=0
cc_318 N_A_c_173_n N_Y_c_741_n 0.00895015f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_319 N_A_c_174_n N_Y_c_741_n 0.00895015f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_320 N_A_c_175_n N_Y_c_741_n 0.0136053f $X=7.205 $Y=1.765 $X2=0 $Y2=0
cc_321 N_A_c_152_n N_Y_c_741_n 0.00204092f $X=7.595 $Y=1.557 $X2=0 $Y2=0
cc_322 N_A_c_153_n N_Y_c_741_n 0.00316449f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_323 N_A_c_154_n N_Y_c_741_n 0.00153204f $X=6.925 $Y=1.515 $X2=0 $Y2=0
cc_324 N_A_c_155_n N_Y_c_741_n 0.00152352f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_325 N_A_c_156_n N_Y_c_741_n 0.00112367f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_326 N_A_c_157_n N_Y_c_741_n 0.00100926f $X=3.11 $Y=1.515 $X2=0 $Y2=0
cc_327 N_A_c_158_n N_Y_c_741_n 0.0011123f $X=4.025 $Y=1.515 $X2=0 $Y2=0
cc_328 N_A_c_159_n N_Y_c_741_n 0.00128431f $X=4.935 $Y=1.515 $X2=0 $Y2=0
cc_329 N_A_c_160_n N_Y_c_741_n 0.0011424f $X=5.93 $Y=1.515 $X2=0 $Y2=0
cc_330 N_A_c_187_n N_Y_c_741_n 0.593249f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_331 N_A_c_163_n N_Y_c_765_n 0.0013431f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_332 N_A_c_164_n N_Y_c_765_n 0.00111176f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_333 N_A_c_153_n N_Y_c_765_n 5.81895e-19 $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_334 N_A_c_187_n N_Y_c_765_n 4.18633e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_335 N_A_c_165_n N_Y_c_769_n 0.0013431f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_336 N_A_c_166_n N_Y_c_769_n 0.00111176f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_337 N_A_c_187_n N_Y_c_769_n 2.74377e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_338 N_A_c_153_n N_Y_c_772_n 7.58724e-19 $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_339 N_A_c_187_n N_Y_c_772_n 2.45236e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_340 N_A_M1002_g N_VGND_c_859_n 0.00525456f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_341 N_A_c_153_n N_VGND_c_859_n 0.00128906f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_342 N_A_M1003_g N_VGND_c_860_n 0.00583652f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_343 N_A_M1005_g N_VGND_c_860_n 0.00227436f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_344 N_A_c_153_n N_VGND_c_860_n 0.00130331f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_345 N_A_c_155_n N_VGND_c_860_n 0.0167206f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_346 N_A_c_187_n N_VGND_c_860_n 0.00144887f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_347 N_A_M1008_g N_VGND_c_861_n 0.00238904f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_348 N_A_M1009_g N_VGND_c_861_n 0.00586329f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_349 N_A_c_153_n N_VGND_c_861_n 0.00130331f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_350 N_A_c_156_n N_VGND_c_861_n 0.018017f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_351 N_A_c_187_n N_VGND_c_861_n 0.00156118f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_352 N_A_M1011_g N_VGND_c_862_n 0.00230839f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_353 N_A_M1012_g N_VGND_c_862_n 0.00231837f $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_354 N_A_c_153_n N_VGND_c_862_n 0.00130331f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_355 N_A_c_157_n N_VGND_c_862_n 0.0173688f $X=3.11 $Y=1.515 $X2=0 $Y2=0
cc_356 N_A_c_187_n N_VGND_c_862_n 0.00150502f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_357 N_A_M1013_g N_VGND_c_863_n 0.00214082f $X=3.785 $Y=0.74 $X2=0 $Y2=0
cc_358 N_A_M1014_g N_VGND_c_863_n 0.0116992f $X=4.215 $Y=0.74 $X2=0 $Y2=0
cc_359 N_A_M1015_g N_VGND_c_863_n 6.07804e-19 $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_360 N_A_c_153_n N_VGND_c_863_n 7.66651e-19 $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_361 N_A_c_158_n N_VGND_c_863_n 0.0166865f $X=4.025 $Y=1.515 $X2=0 $Y2=0
cc_362 N_A_c_187_n N_VGND_c_863_n 0.00144416f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_363 N_A_M1015_g N_VGND_c_864_n 0.00214733f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_364 N_A_M1018_g N_VGND_c_864_n 0.00353535f $X=5.145 $Y=0.74 $X2=0 $Y2=0
cc_365 N_A_c_153_n N_VGND_c_864_n 0.00130331f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_366 N_A_c_159_n N_VGND_c_864_n 0.0163965f $X=4.935 $Y=1.515 $X2=0 $Y2=0
cc_367 N_A_c_187_n N_VGND_c_864_n 0.00161813f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_368 N_A_M1019_g N_VGND_c_865_n 0.00789946f $X=5.575 $Y=0.74 $X2=0 $Y2=0
cc_369 N_A_M1023_g N_VGND_c_865_n 0.00803145f $X=6.145 $Y=0.74 $X2=0 $Y2=0
cc_370 N_A_c_153_n N_VGND_c_865_n 0.00239626f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_371 N_A_c_160_n N_VGND_c_865_n 0.0173678f $X=5.93 $Y=1.515 $X2=0 $Y2=0
cc_372 N_A_c_187_n N_VGND_c_865_n 0.00347842f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_373 N_A_M1027_g N_VGND_c_866_n 0.00814162f $X=6.575 $Y=0.74 $X2=0 $Y2=0
cc_374 N_A_M1029_g N_VGND_c_866_n 0.00688674f $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_375 N_A_c_151_n N_VGND_c_866_n 0.00175563f $X=7.09 $Y=1.515 $X2=0 $Y2=0
cc_376 N_A_c_153_n N_VGND_c_866_n 0.00129147f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_377 N_A_c_154_n N_VGND_c_866_n 0.0176918f $X=6.925 $Y=1.515 $X2=0 $Y2=0
cc_378 N_A_c_187_n N_VGND_c_866_n 0.00408288f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_379 N_A_M1031_g N_VGND_c_868_n 0.00532106f $X=7.595 $Y=0.74 $X2=0 $Y2=0
cc_380 N_A_c_152_n N_VGND_c_868_n 0.00128906f $X=7.595 $Y=1.557 $X2=0 $Y2=0
cc_381 N_A_M1012_g N_VGND_c_869_n 0.00445602f $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_382 N_A_M1013_g N_VGND_c_869_n 0.00461464f $X=3.785 $Y=0.74 $X2=0 $Y2=0
cc_383 N_A_M1014_g N_VGND_c_871_n 0.00429299f $X=4.215 $Y=0.74 $X2=0 $Y2=0
cc_384 N_A_M1015_g N_VGND_c_871_n 0.00434272f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_385 N_A_M1018_g N_VGND_c_873_n 0.00456932f $X=5.145 $Y=0.74 $X2=0 $Y2=0
cc_386 N_A_M1019_g N_VGND_c_873_n 0.00434272f $X=5.575 $Y=0.74 $X2=0 $Y2=0
cc_387 N_A_M1002_g N_VGND_c_875_n 0.00434272f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_388 N_A_M1003_g N_VGND_c_875_n 0.00434272f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_389 N_A_M1005_g N_VGND_c_876_n 0.00445602f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_390 N_A_M1008_g N_VGND_c_876_n 0.00461464f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_391 N_A_M1009_g N_VGND_c_877_n 0.00445602f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_392 N_A_M1011_g N_VGND_c_877_n 0.00445602f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_393 N_A_M1023_g N_VGND_c_878_n 0.00434272f $X=6.145 $Y=0.74 $X2=0 $Y2=0
cc_394 N_A_M1027_g N_VGND_c_878_n 0.00434272f $X=6.575 $Y=0.74 $X2=0 $Y2=0
cc_395 N_A_M1029_g N_VGND_c_879_n 0.00434272f $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_396 N_A_M1031_g N_VGND_c_879_n 0.00434272f $X=7.595 $Y=0.74 $X2=0 $Y2=0
cc_397 N_A_M1002_g N_VGND_c_884_n 0.00823934f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_398 N_A_M1003_g N_VGND_c_884_n 0.00820718f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_399 N_A_M1005_g N_VGND_c_884_n 0.00857405f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_400 N_A_M1008_g N_VGND_c_884_n 0.00908319f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_401 N_A_M1009_g N_VGND_c_884_n 0.00857405f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_402 N_A_M1011_g N_VGND_c_884_n 0.00857405f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_403 N_A_M1012_g N_VGND_c_884_n 0.00857181f $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_404 N_A_M1013_g N_VGND_c_884_n 0.00907773f $X=3.785 $Y=0.74 $X2=0 $Y2=0
cc_405 N_A_M1014_g N_VGND_c_884_n 0.00847524f $X=4.215 $Y=0.74 $X2=0 $Y2=0
cc_406 N_A_M1015_g N_VGND_c_884_n 0.00820718f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_407 N_A_M1018_g N_VGND_c_884_n 0.00890307f $X=5.145 $Y=0.74 $X2=0 $Y2=0
cc_408 N_A_M1019_g N_VGND_c_884_n 0.00821518f $X=5.575 $Y=0.74 $X2=0 $Y2=0
cc_409 N_A_M1023_g N_VGND_c_884_n 0.00821294f $X=6.145 $Y=0.74 $X2=0 $Y2=0
cc_410 N_A_M1027_g N_VGND_c_884_n 0.00821668f $X=6.575 $Y=0.74 $X2=0 $Y2=0
cc_411 N_A_M1029_g N_VGND_c_884_n 0.00821444f $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_412 N_A_M1031_g N_VGND_c_884_n 0.00823934f $X=7.595 $Y=0.74 $X2=0 $Y2=0
cc_413 N_VPWR_c_484_n N_Y_c_627_n 0.014552f $X=2.045 $Y=3.33 $X2=0 $Y2=0
cc_414 N_VPWR_c_467_n N_Y_c_627_n 0.0119791f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_415 N_VPWR_c_485_n N_Y_c_629_n 0.014552f $X=2.995 $Y=3.33 $X2=0 $Y2=0
cc_416 N_VPWR_c_467_n N_Y_c_629_n 0.0119791f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_417 N_VPWR_c_481_n N_Y_c_632_n 0.0128508f $X=4.81 $Y=3.33 $X2=0 $Y2=0
cc_418 N_VPWR_c_467_n N_Y_c_632_n 0.0106368f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_419 N_VPWR_c_469_n N_Y_c_633_n 0.0769517f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_420 N_VPWR_c_470_n N_Y_c_633_n 0.0435606f $X=1.18 $Y=2.105 $X2=0 $Y2=0
cc_421 N_VPWR_c_483_n N_Y_c_633_n 0.0150415f $X=1.055 $Y=3.33 $X2=0 $Y2=0
cc_422 N_VPWR_c_467_n N_Y_c_633_n 0.0117634f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_423 N_VPWR_c_472_n N_Y_c_625_n 0.0419652f $X=3.08 $Y=2.105 $X2=0 $Y2=0
cc_424 N_VPWR_c_473_n N_Y_c_625_n 0.00758346f $X=4.03 $Y=2.105 $X2=0 $Y2=0
cc_425 N_VPWR_c_479_n N_Y_c_625_n 0.0130321f $X=3.915 $Y=3.33 $X2=0 $Y2=0
cc_426 N_VPWR_c_467_n N_Y_c_625_n 0.0107539f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_427 N_VPWR_c_474_n N_Y_c_635_n 0.00909849f $X=4.93 $Y=2.105 $X2=0 $Y2=0
cc_428 N_VPWR_c_475_n N_Y_c_635_n 0.0414821f $X=5.93 $Y=2.105 $X2=0 $Y2=0
cc_429 N_VPWR_c_486_n N_Y_c_635_n 0.0139663f $X=5.765 $Y=3.33 $X2=0 $Y2=0
cc_430 N_VPWR_c_467_n N_Y_c_635_n 0.0115601f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_431 N_VPWR_c_475_n N_Y_c_636_n 0.0425672f $X=5.93 $Y=2.105 $X2=0 $Y2=0
cc_432 N_VPWR_c_476_n N_Y_c_636_n 0.0425672f $X=6.93 $Y=2.105 $X2=0 $Y2=0
cc_433 N_VPWR_c_487_n N_Y_c_636_n 0.014552f $X=6.765 $Y=3.33 $X2=0 $Y2=0
cc_434 N_VPWR_c_467_n N_Y_c_636_n 0.0119791f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_435 N_VPWR_c_476_n N_Y_c_626_n 0.0417838f $X=6.93 $Y=2.105 $X2=0 $Y2=0
cc_436 N_VPWR_c_478_n N_Y_c_626_n 0.00656378f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_437 N_VPWR_c_488_n N_Y_c_626_n 0.0123628f $X=7.735 $Y=3.33 $X2=0 $Y2=0
cc_438 N_VPWR_c_467_n N_Y_c_626_n 0.0101999f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_439 N_VPWR_M1001_d N_Y_c_741_n 0.00432536f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_440 N_VPWR_M1006_d N_Y_c_741_n 0.00560175f $X=1.98 $Y=1.84 $X2=0 $Y2=0
cc_441 N_VPWR_M1010_d N_Y_c_741_n 0.0056392f $X=2.93 $Y=1.84 $X2=0 $Y2=0
cc_442 N_VPWR_M1017_d N_Y_c_741_n 0.00375833f $X=3.88 $Y=1.84 $X2=0 $Y2=0
cc_443 N_VPWR_M1021_d N_Y_c_741_n 0.00251667f $X=4.78 $Y=1.84 $X2=0 $Y2=0
cc_444 N_VPWR_M1024_d N_Y_c_741_n 0.00460059f $X=5.73 $Y=1.84 $X2=0 $Y2=0
cc_445 N_VPWR_M1026_d N_Y_c_741_n 0.00512092f $X=6.73 $Y=1.84 $X2=0 $Y2=0
cc_446 N_VPWR_c_469_n N_Y_c_741_n 0.00161913f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_447 N_VPWR_c_470_n N_Y_c_741_n 0.0278731f $X=1.18 $Y=2.105 $X2=0 $Y2=0
cc_448 N_VPWR_c_471_n N_Y_c_741_n 0.0245664f $X=2.13 $Y=2.105 $X2=0 $Y2=0
cc_449 N_VPWR_c_472_n N_Y_c_741_n 0.0245664f $X=3.08 $Y=2.105 $X2=0 $Y2=0
cc_450 N_VPWR_c_473_n N_Y_c_741_n 0.0236934f $X=4.03 $Y=2.105 $X2=0 $Y2=0
cc_451 N_VPWR_c_474_n N_Y_c_741_n 0.0274622f $X=4.93 $Y=2.105 $X2=0 $Y2=0
cc_452 N_VPWR_c_475_n N_Y_c_741_n 0.0311264f $X=5.93 $Y=2.105 $X2=0 $Y2=0
cc_453 N_VPWR_c_476_n N_Y_c_741_n 0.031051f $X=6.93 $Y=2.105 $X2=0 $Y2=0
cc_454 N_VPWR_c_478_n N_Y_c_741_n 0.00790106f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_455 N_VPWR_c_470_n N_Y_c_765_n 0.0425039f $X=1.18 $Y=2.105 $X2=0 $Y2=0
cc_456 N_VPWR_c_471_n N_Y_c_765_n 0.0675319f $X=2.13 $Y=2.105 $X2=0 $Y2=0
cc_457 N_VPWR_c_471_n N_Y_c_769_n 0.0424691f $X=2.13 $Y=2.105 $X2=0 $Y2=0
cc_458 N_VPWR_c_472_n N_Y_c_769_n 0.0675319f $X=3.08 $Y=2.105 $X2=0 $Y2=0
cc_459 N_VPWR_c_473_n N_Y_c_772_n 0.00811838f $X=4.03 $Y=2.105 $X2=0 $Y2=0
cc_460 N_VPWR_c_474_n N_Y_c_772_n 0.0419037f $X=4.93 $Y=2.105 $X2=0 $Y2=0
cc_461 N_Y_c_613_n N_VGND_c_859_n 0.0307549f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_462 N_Y_c_613_n N_VGND_c_860_n 0.0307549f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_463 N_Y_c_614_n N_VGND_c_860_n 0.028873f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_464 N_Y_c_614_n N_VGND_c_861_n 0.00297007f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_465 N_Y_c_615_n N_VGND_c_861_n 0.029171f $X=2.64 $Y=0.515 $X2=0 $Y2=0
cc_466 N_Y_c_615_n N_VGND_c_862_n 0.0291629f $X=2.64 $Y=0.515 $X2=0 $Y2=0
cc_467 N_Y_c_625_n N_VGND_c_862_n 0.0303029f $X=3.57 $Y=0.515 $X2=0 $Y2=0
cc_468 N_Y_c_616_n N_VGND_c_863_n 0.0272179f $X=4.43 $Y=0.515 $X2=0 $Y2=0
cc_469 N_Y_c_625_n N_VGND_c_863_n 0.0296712f $X=3.57 $Y=0.515 $X2=0 $Y2=0
cc_470 N_Y_c_616_n N_VGND_c_864_n 0.0296586f $X=4.43 $Y=0.515 $X2=0 $Y2=0
cc_471 N_Y_c_617_n N_VGND_c_864_n 0.00429585f $X=5.37 $Y=1.025 $X2=0 $Y2=0
cc_472 N_Y_c_618_n N_VGND_c_864_n 0.0236187f $X=5.36 $Y=0.515 $X2=0 $Y2=0
cc_473 N_Y_c_617_n N_VGND_c_865_n 0.00450652f $X=5.37 $Y=1.025 $X2=0 $Y2=0
cc_474 N_Y_c_618_n N_VGND_c_865_n 0.0246826f $X=5.36 $Y=0.515 $X2=0 $Y2=0
cc_475 N_Y_c_619_n N_VGND_c_865_n 0.0051297f $X=6.36 $Y=1.015 $X2=0 $Y2=0
cc_476 N_Y_c_620_n N_VGND_c_865_n 0.0257017f $X=6.36 $Y=0.515 $X2=0 $Y2=0
cc_477 N_Y_c_619_n N_VGND_c_866_n 0.00490968f $X=6.36 $Y=1.015 $X2=0 $Y2=0
cc_478 N_Y_c_620_n N_VGND_c_866_n 0.0245613f $X=6.36 $Y=0.515 $X2=0 $Y2=0
cc_479 N_Y_c_621_n N_VGND_c_866_n 0.0308181f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_480 N_Y_c_621_n N_VGND_c_868_n 0.0308109f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_481 N_Y_c_625_n N_VGND_c_869_n 0.0130321f $X=3.57 $Y=0.515 $X2=0 $Y2=0
cc_482 N_Y_c_616_n N_VGND_c_871_n 0.0112174f $X=4.43 $Y=0.515 $X2=0 $Y2=0
cc_483 N_Y_c_618_n N_VGND_c_873_n 0.0136595f $X=5.36 $Y=0.515 $X2=0 $Y2=0
cc_484 N_Y_c_613_n N_VGND_c_875_n 0.0144922f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_485 N_Y_c_614_n N_VGND_c_876_n 0.012809f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_486 N_Y_c_615_n N_VGND_c_877_n 0.0136595f $X=2.64 $Y=0.515 $X2=0 $Y2=0
cc_487 N_Y_c_620_n N_VGND_c_878_n 0.0144922f $X=6.36 $Y=0.515 $X2=0 $Y2=0
cc_488 N_Y_c_621_n N_VGND_c_879_n 0.0144922f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_489 N_Y_c_613_n N_VGND_c_884_n 0.0118826f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_490 N_Y_c_614_n N_VGND_c_884_n 0.0105693f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_491 N_Y_c_615_n N_VGND_c_884_n 0.0112404f $X=2.64 $Y=0.515 $X2=0 $Y2=0
cc_492 N_Y_c_616_n N_VGND_c_884_n 0.00922837f $X=4.43 $Y=0.515 $X2=0 $Y2=0
cc_493 N_Y_c_618_n N_VGND_c_884_n 0.0112404f $X=5.36 $Y=0.515 $X2=0 $Y2=0
cc_494 N_Y_c_620_n N_VGND_c_884_n 0.0118826f $X=6.36 $Y=0.515 $X2=0 $Y2=0
cc_495 N_Y_c_621_n N_VGND_c_884_n 0.0118826f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_496 N_Y_c_625_n N_VGND_c_884_n 0.0107539f $X=3.57 $Y=0.515 $X2=0 $Y2=0
