* File: sky130_fd_sc_ls__sdfrtp_4.pex.spice
* Created: Fri Aug 28 14:03:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%A_27_74# 1 2 7 9 11 12 14 17 20 23 27 30 32
+ 33 35 40
c82 35 0 1.02897e-20 $X=2.535 $Y=1.995
c83 9 0 3.56444e-20 $X=1.485 $Y=0.935
r84 35 38 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.54 $Y=1.995
+ $X2=2.54 $Y2=2.09
r85 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.535
+ $Y=1.995 $X2=2.535 $Y2=1.995
r86 31 33 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.09
+ $X2=0.28 $Y2=2.09
r87 30 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=2.09
+ $X2=2.54 $Y2=2.09
r88 30 31 125.914 $w=1.68e-07 $l=1.93e-06 $layer=LI1_cond $X=2.375 $Y=2.09
+ $X2=0.445 $Y2=2.09
r89 28 40 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.975 $Y=1.1 $X2=0.975
+ $Y2=1.01
r90 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.1 $X2=0.975 $Y2=1.1
r91 25 32 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.1
+ $X2=0.24 $Y2=1.1
r92 25 27 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=0.365 $Y=1.1
+ $X2=0.975 $Y2=1.1
r93 21 33 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.09
r94 21 23 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.465
r95 20 33 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.2 $Y=2.005
+ $X2=0.28 $Y2=2.09
r96 19 32 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=0.2 $Y=1.265
+ $X2=0.24 $Y2=1.1
r97 19 20 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.2 $Y=1.265 $X2=0.2
+ $Y2=2.005
r98 15 32 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=0.935
+ $X2=0.24 $Y2=1.1
r99 15 17 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=0.24 $Y=0.935
+ $X2=0.24 $Y2=0.58
r100 12 36 52.2586 $w=2.99e-07 $l=2.69258e-07 $layer=POLY_cond $X=2.495 $Y=2.245
+ $X2=2.535 $Y2=1.995
r101 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.495 $Y=2.245
+ $X2=2.495 $Y2=2.64
r102 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.485 $Y=0.935
+ $X2=1.485 $Y2=0.615
r103 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.01
+ $X2=0.975 $Y2=1.01
r104 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=1.01
+ $X2=1.485 $Y2=0.935
r105 7 8 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.41 $Y=1.01 $X2=1.14
+ $Y2=1.01
r106 2 23 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
r107 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%SCE 2 5 7 9 11 12 14 15 17 20 21 22 25 30
+ 31 32 44 53 55
c87 15 0 1.86316e-19 $X=2.785 $Y=1.05
r88 44 53 1.90404 $w=3.43e-07 $l=5.7e-08 $layer=LI1_cond $X=1.623 $Y=1.662
+ $X2=1.68 $Y2=1.662
r89 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=1.67 $X2=1.45 $Y2=1.67
r90 38 41 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=0.77 $Y=1.67
+ $X2=1.45 $Y2=1.67
r91 32 55 6.34154 $w=3.43e-07 $l=1.01e-07 $layer=LI1_cond $X=1.694 $Y=1.662
+ $X2=1.795 $Y2=1.662
r92 32 53 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=1.694 $Y=1.662
+ $X2=1.68 $Y2=1.662
r93 32 44 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=1.609 $Y=1.662
+ $X2=1.623 $Y2=1.662
r94 32 42 5.31126 $w=3.43e-07 $l=1.59e-07 $layer=LI1_cond $X=1.609 $Y=1.662
+ $X2=1.45 $Y2=1.662
r95 31 42 8.35104 $w=3.43e-07 $l=2.5e-07 $layer=LI1_cond $X=1.2 $Y=1.662
+ $X2=1.45 $Y2=1.662
r96 30 31 16.034 $w=3.43e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.662 $X2=1.2
+ $Y2=1.662
r97 30 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.67 $X2=0.77 $Y2=1.67
r98 25 28 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.57 $Y=1.425
+ $X2=2.57 $Y2=1.575
r99 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.565
+ $Y=1.425 $X2=2.565 $Y2=1.425
r100 22 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=1.575
+ $X2=2.57 $Y2=1.575
r101 22 55 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.405 $Y=1.575
+ $X2=1.795 $Y2=1.575
r102 21 41 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.535 $Y=1.67
+ $X2=1.45 $Y2=1.67
r103 19 38 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.595 $Y=1.67
+ $X2=0.77 $Y2=1.67
r104 19 20 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.595 $Y=1.67
+ $X2=0.505 $Y2=1.67
r105 15 26 72.7678 $w=2.96e-07 $l=4.45814e-07 $layer=POLY_cond $X=2.785 $Y=1.05
+ $X2=2.63 $Y2=1.425
r106 15 17 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.785 $Y=1.05
+ $X2=2.785 $Y2=0.615
r107 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.625 $Y=2.245
+ $X2=1.625 $Y2=2.64
r108 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.625 $Y=2.155
+ $X2=1.625 $Y2=2.245
r109 10 21 30.0773 $w=3.3e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.625 $Y=1.835
+ $X2=1.535 $Y2=1.67
r110 10 11 124.387 $w=1.8e-07 $l=3.2e-07 $layer=POLY_cond $X=1.625 $Y=1.835
+ $X2=1.625 $Y2=2.155
r111 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.64
r112 3 20 34.7346 $w=1.65e-07 $l=1.69926e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.505 $Y2=1.67
r113 3 5 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.495 $Y2=0.58
r114 2 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=2.155
+ $X2=0.505 $Y2=2.245
r115 1 20 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=1.67
r116 1 2 124.387 $w=1.8e-07 $l=3.2e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%D 3 5 6 8 9 12 13 14
c46 6 0 1.02897e-20 $X=2.045 $Y=2.245
r47 12 15 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.952 $Y=1.1
+ $X2=1.952 $Y2=1.265
r48 12 14 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.952 $Y=1.1
+ $X2=1.952 $Y2=0.935
r49 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.1 $X2=1.935 $Y2=1.1
r50 9 13 6.7033 $w=4.53e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.037
+ $X2=1.935 $Y2=1.037
r51 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.045 $Y=2.245
+ $X2=2.045 $Y2=2.64
r52 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.045 $Y=2.155 $X2=2.045
+ $Y2=2.245
r53 5 15 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=2.045 $Y=2.155
+ $X2=2.045 $Y2=1.265
r54 3 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2 $Y=0.615 $X2=2
+ $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%SCD 1 3 6 10 11 12 16
c43 11 0 1.86316e-19 $X=3.12 $Y=1.665
r44 11 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.11 $Y=1.605
+ $X2=3.11 $Y2=2.035
r45 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.105
+ $Y=1.605 $X2=3.105 $Y2=1.605
r46 10 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.105 $Y=1.945
+ $X2=3.105 $Y2=1.605
r47 9 16 40.0117 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.105 $Y=1.44
+ $X2=3.105 $Y2=1.605
r48 6 9 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=3.145 $Y=0.615
+ $X2=3.145 $Y2=1.44
r49 1 10 54.7727 $w=2.64e-07 $l=3.33167e-07 $layer=POLY_cond $X=3.035 $Y=2.245
+ $X2=3.105 $Y2=1.945
r50 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.035 $Y=2.245
+ $X2=3.035 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%CLK 1 3 6 10
c54 10 0 1.48635e-19 $X=4.08 $Y=1.295
c55 1 0 1.68197e-19 $X=4.605 $Y=1.41
r56 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.005
+ $Y=1.455 $X2=4.005 $Y2=1.455
r57 10 14 2.10813 $w=4.08e-07 $l=7.5e-08 $layer=LI1_cond $X=4.08 $Y=1.385
+ $X2=4.005 $Y2=1.385
r58 4 16 21.5811 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=4.645 $Y=1.8
+ $X2=4.645 $Y2=1.545
r59 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.645 $Y=1.8 $X2=4.645
+ $Y2=2.46
r60 1 16 5.75522 $w=3.35e-07 $l=4e-08 $layer=POLY_cond $X=4.605 $Y=1.545
+ $X2=4.645 $Y2=1.545
r61 1 13 86.3284 $w=3.35e-07 $l=6e-07 $layer=POLY_cond $X=4.605 $Y=1.545
+ $X2=4.005 $Y2=1.545
r62 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.605 $Y=1.41
+ $X2=4.605 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%A_1034_392# 1 2 8 9 11 12 16 18 20 21 22 23
+ 25 29 31 32 33 34 36 39 42 43 44 46 48 49 51 58 59 67 68 70
c229 70 0 1.2914e-19 $X=6.065 $Y=1.66
c230 68 0 1.40436e-19 $X=9.33 $Y=1.07
c231 67 0 1.39722e-19 $X=9.25 $Y=1.07
c232 58 0 2.21688e-19 $X=5.407 $Y=1.24
c233 31 0 7.48709e-20 $X=5.535 $Y=1.585
r234 67 76 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.25 $Y=1.07 $X2=9.25
+ $Y2=1.16
r235 66 68 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.25 $Y=1.07 $X2=9.33
+ $Y2=1.07
r236 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.25
+ $Y=1.07 $X2=9.25 $Y2=1.07
r237 63 66 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.91 $Y=1.07
+ $X2=9.25 $Y2=1.07
r238 59 61 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.14 $Y=0.415
+ $X2=7.14 $Y2=0.665
r239 57 58 13.0794 $w=4.03e-07 $l=3.2e-07 $layer=LI1_cond $X=5.407 $Y=0.92
+ $X2=5.407 $Y2=1.24
r240 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.79
+ $Y=2.215 $X2=9.79 $Y2=2.215
r241 49 51 13.7196 $w=3.13e-07 $l=3.75e-07 $layer=LI1_cond $X=9.415 $Y=2.222
+ $X2=9.79 $Y2=2.222
r242 48 49 7.64049 $w=3.15e-07 $l=1.94921e-07 $layer=LI1_cond $X=9.33 $Y=2.065
+ $X2=9.415 $Y2=2.222
r243 47 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.33 $Y=1.235
+ $X2=9.33 $Y2=1.07
r244 47 48 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=9.33 $Y=1.235
+ $X2=9.33 $Y2=2.065
r245 46 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.91 $Y=0.905
+ $X2=8.91 $Y2=1.07
r246 45 46 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=8.91 $Y=0.425
+ $X2=8.91 $Y2=0.905
r247 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.825 $Y=0.34
+ $X2=8.91 $Y2=0.425
r248 43 44 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.825 $Y=0.34
+ $X2=8.1 $Y2=0.34
r249 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.015 $Y=0.425
+ $X2=8.1 $Y2=0.34
r250 41 42 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.015 $Y=0.425
+ $X2=8.015 $Y2=0.58
r251 40 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.225 $Y=0.665
+ $X2=7.14 $Y2=0.665
r252 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.93 $Y=0.665
+ $X2=8.015 $Y2=0.58
r253 39 40 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=7.93 $Y=0.665
+ $X2=7.225 $Y2=0.665
r254 37 73 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.065 $Y=1.75
+ $X2=6.065 $Y2=1.915
r255 37 70 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.065 $Y=1.75
+ $X2=6.065 $Y2=1.66
r256 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.065
+ $Y=1.75 $X2=6.065 $Y2=1.75
r257 34 56 11.5779 $w=3.53e-07 $l=4.42691e-07 $layer=LI1_cond $X=5.655 $Y=1.75
+ $X2=5.405 $Y2=2.085
r258 34 36 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.655 $Y=1.75
+ $X2=6.065 $Y2=1.75
r259 32 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.055 $Y=0.415
+ $X2=7.14 $Y2=0.415
r260 32 33 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=7.055 $Y=0.415
+ $X2=5.62 $Y2=0.415
r261 31 34 8.99262 $w=3.53e-07 $l=2.16852e-07 $layer=LI1_cond $X=5.535 $Y=1.585
+ $X2=5.655 $Y2=1.75
r262 31 58 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.535 $Y=1.585
+ $X2=5.535 $Y2=1.24
r263 29 57 4.97969 $w=4.03e-07 $l=1.75e-07 $layer=LI1_cond $X=5.417 $Y=0.745
+ $X2=5.417 $Y2=0.92
r264 26 33 8.41448 $w=1.7e-07 $l=2.41793e-07 $layer=LI1_cond $X=5.417 $Y=0.5
+ $X2=5.62 $Y2=0.415
r265 26 29 6.97157 $w=4.03e-07 $l=2.45e-07 $layer=LI1_cond $X=5.417 $Y=0.5
+ $X2=5.417 $Y2=0.745
r266 23 52 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=9.835 $Y=2.465
+ $X2=9.79 $Y2=2.215
r267 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.835 $Y=2.465
+ $X2=9.835 $Y2=2.75
r268 21 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.085 $Y=1.16
+ $X2=9.25 $Y2=1.16
r269 21 22 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=9.085 $Y=1.16
+ $X2=8.725 $Y2=1.16
r270 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.65 $Y=1.085
+ $X2=8.725 $Y2=1.16
r271 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.65 $Y=1.085
+ $X2=8.65 $Y2=0.69
r272 14 16 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=6.535 $Y=1.585
+ $X2=6.535 $Y2=0.9
r273 13 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.23 $Y=1.66
+ $X2=6.065 $Y2=1.66
r274 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.46 $Y=1.66
+ $X2=6.535 $Y2=1.585
r275 12 13 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=6.46 $Y=1.66
+ $X2=6.23 $Y2=1.66
r276 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.135 $Y=2.24
+ $X2=6.135 $Y2=2.525
r277 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.135 $Y=2.15 $X2=6.135
+ $Y2=2.24
r278 8 73 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=6.135 $Y=2.15
+ $X2=6.135 $Y2=1.915
r279 2 56 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.96 $X2=5.32 $Y2=2.085
r280 1 29 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=5.23
+ $Y=0.595 $X2=5.37 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%A_1367_112# 1 2 9 12 13 15 18 19 22 24 25
+ 27 33 34
c110 34 0 2.99465e-19 $X=8.57 $Y=0.842
c111 22 0 1.09068e-19 $X=7.325 $Y=1.005
c112 18 0 3.61087e-19 $X=7.19 $Y=1.78
c113 9 0 1.54393e-19 $X=6.91 $Y=0.9
r114 40 42 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=6.91 $Y=1.78
+ $X2=7.025 $Y2=1.78
r115 32 34 3.26203 $w=4.93e-07 $l=1.35e-07 $layer=LI1_cond $X=8.435 $Y=0.842
+ $X2=8.57 $Y2=0.842
r116 32 33 9.48656 $w=4.93e-07 $l=1.65e-07 $layer=LI1_cond $X=8.435 $Y=0.842
+ $X2=8.27 $Y2=0.842
r117 27 29 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=8.9 $Y=1.88 $X2=8.9
+ $Y2=2.59
r118 25 36 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.9 $Y=1.49
+ $X2=8.57 $Y2=1.49
r119 25 27 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=8.9 $Y=1.575
+ $X2=8.9 $Y2=1.88
r120 24 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.57 $Y=1.405
+ $X2=8.57 $Y2=1.49
r121 23 34 7.09362 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=8.57 $Y=1.09
+ $X2=8.57 $Y2=0.842
r122 23 24 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.57 $Y=1.09
+ $X2=8.57 $Y2=1.405
r123 22 33 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=7.325 $Y=1.005
+ $X2=8.27 $Y2=1.005
r124 19 42 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.19 $Y=1.78
+ $X2=7.025 $Y2=1.78
r125 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.19
+ $Y=1.78 $X2=7.19 $Y2=1.78
r126 16 22 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=7.19 $Y=1.09
+ $X2=7.325 $Y2=1.005
r127 16 18 29.4513 $w=2.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.19 $Y=1.09
+ $X2=7.19 $Y2=1.78
r128 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.025 $Y=2.24
+ $X2=7.025 $Y2=2.525
r129 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.025 $Y=2.15
+ $X2=7.025 $Y2=2.24
r130 11 42 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.025 $Y=1.945
+ $X2=7.025 $Y2=1.78
r131 11 12 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=7.025 $Y=1.945
+ $X2=7.025 $Y2=2.15
r132 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.91 $Y=1.615
+ $X2=6.91 $Y2=1.78
r133 7 9 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=6.91 $Y=1.615
+ $X2=6.91 $Y2=0.9
r134 2 29 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=8.75
+ $Y=1.735 $X2=8.9 $Y2=2.59
r135 2 27 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.75
+ $Y=1.735 $X2=8.9 $Y2=1.88
r136 1 32 182 $w=1.7e-07 $l=5.24404e-07 $layer=licon1_NDIFF $count=1 $X=8.25
+ $Y=0.37 $X2=8.435 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%RESET_B 2 6 7 9 10 11 15 16 17 18 20 22 25
+ 28 29 31 33 34 35 36 37 44 45 48 51 53 61 62
c226 53 0 1.27018e-19 $X=7.67 $Y=2.03
c227 10 0 1.62559e-19 $X=7.225 $Y=0.18
c228 7 0 9.42244e-20 $X=3.605 $Y=2.245
r229 60 62 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=10.75 $Y=1.985
+ $X2=10.94 $Y2=1.985
r230 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.75
+ $Y=1.985 $X2=10.75 $Y2=1.985
r231 57 60 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=10.63 $Y=1.985
+ $X2=10.75 $Y2=1.985
r232 53 55 41.7374 $w=3.58e-07 $l=3.1e-07 $layer=POLY_cond $X=7.67 $Y=2.03
+ $X2=7.98 $Y2=2.03
r233 52 53 0.673184 $w=3.58e-07 $l=5e-09 $layer=POLY_cond $X=7.665 $Y=2.03
+ $X2=7.67 $Y2=2.03
r234 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.995 $X2=3.95 $Y2=1.995
r235 48 50 46.4497 $w=3.58e-07 $l=3.45e-07 $layer=POLY_cond $X=3.605 $Y=2.037
+ $X2=3.95 $Y2=2.037
r236 47 48 6.73184 $w=3.58e-07 $l=5e-08 $layer=POLY_cond $X=3.555 $Y=2.037
+ $X2=3.605 $Y2=2.037
r237 45 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r238 44 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.98
+ $Y=1.985 $X2=7.98 $Y2=1.985
r239 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r240 39 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r241 37 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=2.035
+ $X2=7.92 $Y2=2.035
r242 36 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r243 36 37 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=8.065 $Y2=2.035
r244 35 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r245 34 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r246 34 35 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=4.225 $Y2=2.035
r247 32 33 40.1667 $w=1.7e-07 $l=9.5e-08 $layer=POLY_cond $X=3.565 $Y=0.965
+ $X2=3.565 $Y2=1.06
r248 29 31 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.94 $Y=2.465
+ $X2=10.94 $Y2=2.75
r249 28 29 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.94 $Y=2.375
+ $X2=10.94 $Y2=2.465
r250 27 62 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.94 $Y=2.15
+ $X2=10.94 $Y2=1.985
r251 27 28 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=10.94 $Y=2.15
+ $X2=10.94 $Y2=2.375
r252 23 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.63 $Y=1.82
+ $X2=10.63 $Y2=1.985
r253 23 25 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=10.63 $Y=1.82
+ $X2=10.63 $Y2=0.58
r254 22 53 23.1716 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.67 $Y=1.82
+ $X2=7.67 $Y2=2.03
r255 21 22 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=7.67 $Y=1.335
+ $X2=7.67 $Y2=1.82
r256 18 52 23.1716 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.665 $Y=2.24
+ $X2=7.665 $Y2=2.03
r257 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.665 $Y=2.24
+ $X2=7.665 $Y2=2.525
r258 16 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.595 $Y=1.26
+ $X2=7.67 $Y2=1.335
r259 16 17 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=7.595 $Y=1.26
+ $X2=7.375 $Y2=1.26
r260 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.3 $Y=1.185
+ $X2=7.375 $Y2=1.26
r261 13 15 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.3 $Y=1.185
+ $X2=7.3 $Y2=0.9
r262 12 15 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=7.3 $Y=0.255
+ $X2=7.3 $Y2=0.9
r263 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.225 $Y=0.18
+ $X2=7.3 $Y2=0.255
r264 10 11 1833.14 $w=1.5e-07 $l=3.575e-06 $layer=POLY_cond $X=7.225 $Y=0.18
+ $X2=3.65 $Y2=0.18
r265 7 48 23.1716 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.605 $Y=2.245
+ $X2=3.605 $Y2=2.037
r266 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.605 $Y=2.245
+ $X2=3.605 $Y2=2.64
r267 6 32 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.575 $Y=0.615
+ $X2=3.575 $Y2=0.965
r268 3 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.575 $Y=0.255
+ $X2=3.65 $Y2=0.18
r269 3 6 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.575 $Y=0.255
+ $X2=3.575 $Y2=0.615
r270 2 47 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.555 $Y=1.83
+ $X2=3.555 $Y2=2.037
r271 2 33 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=3.555 $Y=1.83
+ $X2=3.555 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%A_1236_138# 1 2 3 12 14 16 18 19 23 26 27
+ 30 31 33 34 37 41
c135 34 0 7.6904e-20 $X=8.15 $Y=1.41
c136 27 0 9.53373e-20 $X=7.495 $Y=2.405
c137 23 0 6.13201e-21 $X=6.715 $Y=0.99
c138 12 0 3.00719e-20 $X=8.175 $Y=0.74
r139 37 39 4.46107 $w=3.08e-07 $l=1.2e-07 $layer=LI1_cond $X=6.315 $Y=0.87
+ $X2=6.315 $Y2=0.99
r140 34 47 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=8.15 $Y=1.41
+ $X2=8.15 $Y2=1.52
r141 34 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.15 $Y=1.41
+ $X2=8.15 $Y2=1.245
r142 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.15
+ $Y=1.41 $X2=8.15 $Y2=1.41
r143 31 33 17.744 $w=3.13e-07 $l=4.85e-07 $layer=LI1_cond $X=7.665 $Y=1.417
+ $X2=8.15 $Y2=1.417
r144 30 44 11.6012 $w=3.26e-07 $l=4.04191e-07 $layer=LI1_cond $X=7.58 $Y=2.32
+ $X2=7.89 $Y2=2.537
r145 29 31 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=7.58 $Y=1.575
+ $X2=7.665 $Y2=1.417
r146 29 30 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.58 $Y=1.575
+ $X2=7.58 $Y2=2.32
r147 28 41 3.70735 $w=2.5e-07 $l=1.69245e-07 $layer=LI1_cond $X=6.885 $Y=2.405
+ $X2=6.8 $Y2=2.537
r148 27 30 5.9625 $w=3.26e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.495 $Y=2.405
+ $X2=7.58 $Y2=2.32
r149 27 28 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.495 $Y=2.405
+ $X2=6.885 $Y2=2.405
r150 26 41 2.76166 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=6.8 $Y=2.32 $X2=6.8
+ $Y2=2.537
r151 25 26 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=6.8 $Y=1.075
+ $X2=6.8 $Y2=2.32
r152 24 39 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=6.47 $Y=0.99
+ $X2=6.315 $Y2=0.99
r153 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.715 $Y=0.99
+ $X2=6.8 $Y2=1.075
r154 23 24 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.715 $Y=0.99
+ $X2=6.47 $Y2=0.99
r155 19 41 3.70735 $w=2.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=6.715 $Y=2.59
+ $X2=6.8 $Y2=2.537
r156 19 21 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.715 $Y=2.59
+ $X2=6.41 $Y2=2.59
r157 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.675 $Y=1.66
+ $X2=8.675 $Y2=2.235
r158 15 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.315 $Y=1.52
+ $X2=8.15 $Y2=1.52
r159 14 16 26.9307 $w=1.5e-07 $l=1.79444e-07 $layer=POLY_cond $X=8.585 $Y=1.52
+ $X2=8.675 $Y2=1.66
r160 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.585 $Y=1.52
+ $X2=8.315 $Y2=1.52
r161 12 46 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.175 $Y=0.74
+ $X2=8.175 $Y2=1.245
r162 3 44 600 $w=1.7e-07 $l=2.85307e-07 $layer=licon1_PDIFF $count=1 $X=7.74
+ $Y=2.315 $X2=7.89 $Y2=2.535
r163 2 21 600 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=6.21
+ $Y=2.315 $X2=6.41 $Y2=2.59
r164 1 37 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.18 $Y=0.69
+ $X2=6.32 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%A_837_98# 1 2 9 13 14 16 17 18 19 20 22 24
+ 25 26 27 29 30 32 33 37 38 39 42 46 48 49 51 52 54 58 60 66 69 70
c205 69 0 3.00264e-19 $X=5.115 $Y=1.485
c206 60 0 9.42244e-20 $X=4.425 $Y=1.905
c207 38 0 1.10364e-19 $X=9.625 $Y=1.585
c208 22 0 6.13201e-21 $X=6.105 $Y=1.185
c209 17 0 4.8605e-20 $X=5.615 $Y=3.075
c210 9 0 4.7366e-20 $X=5.095 $Y=2.46
r211 69 70 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.115 $Y=1.485
+ $X2=5.115 $Y2=1.41
r212 67 72 50.583 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=5.115 $Y=1.61
+ $X2=5.115 $Y2=1.8
r213 67 69 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.115 $Y=1.61
+ $X2=5.115 $Y2=1.485
r214 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.115
+ $Y=1.61 $X2=5.115 $Y2=1.61
r215 60 63 11.0909 $w=1.78e-07 $l=1.8e-07 $layer=LI1_cond $X=4.425 $Y=1.905
+ $X2=4.425 $Y2=2.085
r216 56 58 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=4.33 $Y=0.65
+ $X2=4.45 $Y2=0.65
r217 54 66 10.218 $w=3.43e-07 $l=2.6533e-07 $layer=LI1_cond $X=4.89 $Y=1.41
+ $X2=5.042 $Y2=1.61
r218 53 54 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.89 $Y=1.09
+ $X2=4.89 $Y2=1.41
r219 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.805 $Y=1.005
+ $X2=4.89 $Y2=1.09
r220 51 52 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.805 $Y=1.005
+ $X2=4.535 $Y2=1.005
r221 50 60 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.515 $Y=1.905
+ $X2=4.425 $Y2=1.905
r222 49 66 10.4927 $w=3.43e-07 $l=3.96157e-07 $layer=LI1_cond $X=4.805 $Y=1.905
+ $X2=5.042 $Y2=1.61
r223 49 50 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.805 $Y=1.905
+ $X2=4.515 $Y2=1.905
r224 48 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.45 $Y=0.92
+ $X2=4.535 $Y2=1.005
r225 47 58 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.45 $Y=0.75 $X2=4.45
+ $Y2=0.65
r226 47 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.45 $Y=0.75
+ $X2=4.45 $Y2=0.92
r227 44 45 69.0764 $w=1.57e-07 $l=2.25e-07 $layer=POLY_cond $X=5.63 $Y=1.26
+ $X2=5.63 $Y2=1.485
r228 40 42 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=9.7 $Y=1.51 $X2=9.7
+ $Y2=0.58
r229 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.625 $Y=1.585
+ $X2=9.7 $Y2=1.51
r230 38 39 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=9.625 $Y=1.585
+ $X2=9.2 $Y2=1.585
r231 35 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.125 $Y=2.81
+ $X2=9.125 $Y2=2.235
r232 34 39 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.125 $Y=1.66
+ $X2=9.2 $Y2=1.585
r233 34 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.125 $Y=1.66
+ $X2=9.125 $Y2=2.235
r234 32 35 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.125 $Y=2.9
+ $X2=9.125 $Y2=2.81
r235 32 33 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=9.125 $Y=2.9
+ $X2=9.125 $Y2=3.075
r236 31 46 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.725 $Y=3.15
+ $X2=6.635 $Y2=3.15
r237 30 33 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.035 $Y=3.15
+ $X2=9.125 $Y2=3.075
r238 30 31 1184.49 $w=1.5e-07 $l=2.31e-06 $layer=POLY_cond $X=9.035 $Y=3.15
+ $X2=6.725 $Y2=3.15
r239 27 29 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.635 $Y=2.81
+ $X2=6.635 $Y2=2.525
r240 26 46 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.635 $Y=3.075
+ $X2=6.635 $Y2=3.15
r241 25 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.635 $Y=2.9
+ $X2=6.635 $Y2=2.81
r242 25 26 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=6.635 $Y=2.9
+ $X2=6.635 $Y2=3.075
r243 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.105 $Y=1.185
+ $X2=6.105 $Y2=0.9
r244 21 44 3.92347 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.72 $Y=1.26 $X2=5.63
+ $Y2=1.26
r245 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.03 $Y=1.26
+ $X2=6.105 $Y2=1.185
r246 20 21 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=6.03 $Y=1.26
+ $X2=5.72 $Y2=1.26
r247 18 46 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.545 $Y=3.15
+ $X2=6.635 $Y2=3.15
r248 18 19 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=6.545 $Y=3.15
+ $X2=5.69 $Y2=3.15
r249 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.615 $Y=3.075
+ $X2=5.69 $Y2=3.15
r250 16 45 23.0255 $w=1.57e-07 $l=8.21584e-08 $layer=POLY_cond $X=5.615 $Y=1.56
+ $X2=5.63 $Y2=1.485
r251 16 17 776.84 $w=1.5e-07 $l=1.515e-06 $layer=POLY_cond $X=5.615 $Y=1.56
+ $X2=5.615 $Y2=3.075
r252 15 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.28 $Y=1.485
+ $X2=5.115 $Y2=1.485
r253 14 45 3.92347 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.54 $Y=1.485
+ $X2=5.63 $Y2=1.485
r254 14 15 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=5.54 $Y=1.485
+ $X2=5.28 $Y2=1.485
r255 13 70 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.155 $Y=0.965
+ $X2=5.155 $Y2=1.41
r256 9 72 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.095 $Y=2.46
+ $X2=5.095 $Y2=1.8
r257 2 63 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.96 $X2=4.42 $Y2=2.085
r258 1 56 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=4.185
+ $Y=0.49 $X2=4.33 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%A_2003_48# 1 2 9 12 13 15 16 18 25 27 28 33
+ 34 37
c89 25 0 1.05829e-19 $X=11.5 $Y=1.385
r90 36 37 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.245 $Y=1.47
+ $X2=11.5 $Y2=1.47
r91 33 34 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=11.165 $Y=2.75
+ $X2=11.165 $Y2=2.52
r92 28 41 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.18 $Y=1.39
+ $X2=10.18 $Y2=1.555
r93 28 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.18 $Y=1.39
+ $X2=10.18 $Y2=1.225
r94 27 30 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=10.18 $Y=1.39 $X2=10.18
+ $Y2=1.47
r95 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.18
+ $Y=1.39 $X2=10.18 $Y2=1.39
r96 25 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.5 $Y=1.385
+ $X2=11.5 $Y2=1.47
r97 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.5 $Y=0.715
+ $X2=11.5 $Y2=1.385
r98 22 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.245 $Y=1.555
+ $X2=11.245 $Y2=1.47
r99 22 34 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=11.245 $Y=1.555
+ $X2=11.245 $Y2=2.52
r100 18 24 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.415 $Y=0.55
+ $X2=11.5 $Y2=0.715
r101 18 20 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=11.415 $Y=0.55
+ $X2=11.24 $Y2=0.55
r102 17 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.345 $Y=1.47
+ $X2=10.18 $Y2=1.47
r103 16 36 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=11.16 $Y=1.47
+ $X2=11.245 $Y2=1.47
r104 16 17 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=11.16 $Y=1.47
+ $X2=10.345 $Y2=1.47
r105 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.255 $Y=2.465
+ $X2=10.255 $Y2=2.75
r106 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.255 $Y=2.375
+ $X2=10.255 $Y2=2.465
r107 12 41 318.742 $w=1.8e-07 $l=8.2e-07 $layer=POLY_cond $X=10.255 $Y=2.375
+ $X2=10.255 $Y2=1.555
r108 9 40 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=10.09 $Y=0.58
+ $X2=10.09 $Y2=1.225
r109 2 33 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=11.015
+ $Y=2.54 $X2=11.165 $Y2=2.75
r110 1 20 182 $w=1.7e-07 $l=2.52785e-07 $layer=licon1_NDIFF $count=1 $X=11.065
+ $Y=0.37 $X2=11.24 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%A_1745_74# 1 2 7 9 12 13 14 16 17 19 21 22
+ 24 26 27 29 31 32 33 34 35 39 44 46 47 49 50 52 53 54 64
c164 29 0 1.81891e-19 $X=12.49 $Y=1.765
c165 26 0 1.05829e-19 $X=12.055 $Y=1.615
c166 22 0 1.86508e-19 $X=12.055 $Y=1.185
r167 63 64 35.0294 $w=4.35e-07 $l=7.5e-08 $layer=POLY_cond $X=11.46 $Y=1.117
+ $X2=11.535 $Y2=1.117
r168 58 63 48.5836 $w=4.35e-07 $l=3.8e-07 $layer=POLY_cond $X=11.08 $Y=1.117
+ $X2=11.46 $Y2=1.117
r169 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.08
+ $Y=1.065 $X2=11.08 $Y2=1.065
r170 54 57 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=11.08 $Y=0.97
+ $X2=11.08 $Y2=1.065
r171 51 52 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=10.21 $Y=1.895
+ $X2=10.21 $Y2=2.55
r172 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.125 $Y=1.81
+ $X2=10.21 $Y2=1.895
r173 49 50 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.125 $Y=1.81
+ $X2=9.755 $Y2=1.81
r174 48 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.755 $Y=0.97
+ $X2=9.67 $Y2=0.97
r175 47 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.915 $Y=0.97
+ $X2=11.08 $Y2=0.97
r176 47 48 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=10.915 $Y=0.97
+ $X2=9.755 $Y2=0.97
r177 46 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.67 $Y=1.725
+ $X2=9.755 $Y2=1.81
r178 45 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.67 $Y=1.055
+ $X2=9.67 $Y2=0.97
r179 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.67 $Y=1.055
+ $X2=9.67 $Y2=1.725
r180 44 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.67 $Y=0.885
+ $X2=9.67 $Y2=0.97
r181 43 44 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=9.67 $Y=0.735
+ $X2=9.67 $Y2=0.885
r182 39 52 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.125 $Y=2.715
+ $X2=10.21 $Y2=2.55
r183 39 41 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=10.125 $Y=2.715
+ $X2=9.52 $Y2=2.715
r184 35 43 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.585 $Y=0.57
+ $X2=9.67 $Y2=0.735
r185 35 37 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=9.585 $Y=0.57
+ $X2=9.405 $Y2=0.57
r186 29 31 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=12.49 $Y=1.765
+ $X2=12.49 $Y2=2.26
r187 28 33 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=12.13 $Y=1.69
+ $X2=12.04 $Y2=1.69
r188 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.415 $Y=1.69
+ $X2=12.49 $Y2=1.765
r189 27 28 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.415 $Y=1.69
+ $X2=12.13 $Y2=1.69
r190 26 33 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=12.055 $Y=1.615
+ $X2=12.04 $Y2=1.69
r191 25 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.055 $Y=1.335
+ $X2=12.055 $Y2=1.26
r192 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=12.055 $Y=1.335
+ $X2=12.055 $Y2=1.615
r193 22 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.055 $Y=1.185
+ $X2=12.055 $Y2=1.26
r194 22 24 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=12.055 $Y=1.185
+ $X2=12.055 $Y2=0.74
r195 19 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.04 $Y=1.765
+ $X2=12.04 $Y2=1.69
r196 19 21 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=12.04 $Y=1.765
+ $X2=12.04 $Y2=2.26
r197 17 34 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.98 $Y=1.26
+ $X2=12.055 $Y2=1.26
r198 17 64 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=11.98 $Y=1.26
+ $X2=11.535 $Y2=1.26
r199 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.475 $Y=2.465
+ $X2=11.475 $Y2=2.75
r200 13 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.475 $Y=2.375
+ $X2=11.475 $Y2=2.465
r201 12 32 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.475 $Y=1.665
+ $X2=11.475 $Y2=1.575
r202 12 13 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=11.475 $Y=1.665
+ $X2=11.475 $Y2=2.375
r203 10 63 27.9254 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=11.46 $Y=1.335
+ $X2=11.46 $Y2=1.117
r204 10 32 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=11.46 $Y=1.335
+ $X2=11.46 $Y2=1.575
r205 7 58 11.5066 $w=4.35e-07 $l=9e-08 $layer=POLY_cond $X=10.99 $Y=1.117
+ $X2=11.08 $Y2=1.117
r206 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.99 $Y=0.9
+ $X2=10.99 $Y2=0.58
r207 2 41 600 $w=1.7e-07 $l=1.12872e-06 $layer=licon1_PDIFF $count=1 $X=9.2
+ $Y=1.735 $X2=9.52 $Y2=2.715
r208 1 37 182 $w=1.7e-07 $l=7.73563e-07 $layer=licon1_NDIFF $count=1 $X=8.725
+ $Y=0.37 $X2=9.405 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%A_2339_74# 1 2 7 9 10 11 12 14 15 17 18 20
+ 21 23 24 26 27 29 30 32 35 39 41 46 59
c117 59 0 2.76177e-20 $X=14.375 $Y=1.495
c118 21 0 1.4738e-19 $X=13.925 $Y=1.765
r119 59 60 1.0783 $w=4.47e-07 $l=1e-08 $layer=POLY_cond $X=14.375 $Y=1.495
+ $X2=14.385 $Y2=1.495
r120 58 59 45.2886 $w=4.47e-07 $l=4.2e-07 $layer=POLY_cond $X=13.955 $Y=1.495
+ $X2=14.375 $Y2=1.495
r121 57 58 3.2349 $w=4.47e-07 $l=3e-08 $layer=POLY_cond $X=13.925 $Y=1.495
+ $X2=13.955 $Y2=1.495
r122 54 55 48.5235 $w=4.47e-07 $l=4.5e-07 $layer=POLY_cond $X=13.025 $Y=1.495
+ $X2=13.475 $Y2=1.495
r123 49 51 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=11.84 $Y=1.435
+ $X2=12.265 $Y2=1.435
r124 47 57 25.8792 $w=4.47e-07 $l=2.4e-07 $layer=POLY_cond $X=13.685 $Y=1.495
+ $X2=13.925 $Y2=1.495
r125 47 55 22.6443 $w=4.47e-07 $l=2.1e-07 $layer=POLY_cond $X=13.685 $Y=1.495
+ $X2=13.475 $Y2=1.495
r126 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.685
+ $Y=1.435 $X2=13.685 $Y2=1.435
r127 44 54 2.1566 $w=4.47e-07 $l=2e-08 $layer=POLY_cond $X=13.005 $Y=1.495
+ $X2=13.025 $Y2=1.495
r128 44 52 9.7047 $w=4.47e-07 $l=9e-08 $layer=POLY_cond $X=13.005 $Y=1.495
+ $X2=12.915 $Y2=1.495
r129 43 46 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=13.005 $Y=1.435
+ $X2=13.685 $Y2=1.435
r130 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.005
+ $Y=1.435 $X2=13.005 $Y2=1.435
r131 41 51 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.43 $Y=1.435
+ $X2=12.265 $Y2=1.435
r132 41 43 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=12.43 $Y=1.435
+ $X2=13.005 $Y2=1.435
r133 37 51 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=12.265 $Y=1.6
+ $X2=12.265 $Y2=1.435
r134 37 39 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=12.265 $Y=1.6
+ $X2=12.265 $Y2=1.985
r135 33 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.84 $Y=1.27
+ $X2=11.84 $Y2=1.435
r136 33 35 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=11.84 $Y=1.27
+ $X2=11.84 $Y2=0.515
r137 30 60 28.6003 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=14.385 $Y=1.225
+ $X2=14.385 $Y2=1.495
r138 30 32 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=14.385 $Y=1.225
+ $X2=14.385 $Y2=0.74
r139 27 59 28.6003 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=14.375 $Y=1.765
+ $X2=14.375 $Y2=1.495
r140 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=14.375 $Y=1.765
+ $X2=14.375 $Y2=2.4
r141 24 58 28.6003 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=13.955 $Y=1.225
+ $X2=13.955 $Y2=1.495
r142 24 26 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=13.955 $Y=1.225
+ $X2=13.955 $Y2=0.74
r143 21 57 28.6003 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=13.925 $Y=1.765
+ $X2=13.925 $Y2=1.495
r144 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.925 $Y=1.765
+ $X2=13.925 $Y2=2.4
r145 18 55 28.6003 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=13.475 $Y=1.765
+ $X2=13.475 $Y2=1.495
r146 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.475 $Y=1.765
+ $X2=13.475 $Y2=2.4
r147 15 54 28.6003 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=13.025 $Y=1.765
+ $X2=13.025 $Y2=1.495
r148 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.025 $Y=1.765
+ $X2=13.025 $Y2=2.4
r149 12 52 28.6003 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=12.915 $Y=1.225
+ $X2=12.915 $Y2=1.495
r150 12 14 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=12.915 $Y=1.225
+ $X2=12.915 $Y2=0.74
r151 10 52 30.9047 $w=4.47e-07 $l=2.29456e-07 $layer=POLY_cond $X=12.84 $Y=1.3
+ $X2=12.915 $Y2=1.495
r152 10 11 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=12.84 $Y=1.3
+ $X2=12.56 $Y2=1.3
r153 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.485 $Y=1.225
+ $X2=12.56 $Y2=1.3
r154 7 9 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=12.485 $Y=1.225
+ $X2=12.485 $Y2=0.74
r155 2 39 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=12.115
+ $Y=1.84 $X2=12.265 $Y2=1.985
r156 1 35 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=11.695
+ $Y=0.37 $X2=11.84 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 43 47 53
+ 57 61 65 69 71 73 76 77 79 80 81 83 88 100 114 118 123 129 136 139 142 145 148
+ 151 155
c194 2 0 1.19423e-19 $X=3.11 $Y=2.32
r195 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r196 151 152 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r197 149 152 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r198 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r199 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r200 142 143 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r201 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r202 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r203 129 132 11.1084 $w=9.48e-07 $l=8.65e-07 $layer=LI1_cond $X=1.09 $Y=2.465
+ $X2=1.09 $Y2=3.33
r204 127 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=14.64 $Y2=3.33
r205 127 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r206 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r207 124 151 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.865 $Y=3.33
+ $X2=13.74 $Y2=3.33
r208 124 126 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.865 $Y=3.33
+ $X2=14.16 $Y2=3.33
r209 123 154 4.40486 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=14.47 $Y=3.33
+ $X2=14.675 $Y2=3.33
r210 123 126 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=14.47 $Y=3.33
+ $X2=14.16 $Y2=3.33
r211 122 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r212 122 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r213 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r214 119 145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.9 $Y=3.33
+ $X2=11.775 $Y2=3.33
r215 119 121 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.9 $Y=3.33
+ $X2=12.24 $Y2=3.33
r216 118 148 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.635 $Y=3.33
+ $X2=12.76 $Y2=3.33
r217 118 121 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.635 $Y=3.33
+ $X2=12.24 $Y2=3.33
r218 117 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r219 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r220 114 145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.65 $Y=3.33
+ $X2=11.775 $Y2=3.33
r221 114 116 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=11.65 $Y=3.33
+ $X2=11.28 $Y2=3.33
r222 113 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r223 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r224 110 113 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r225 110 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r226 109 112 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r227 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r228 107 142 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.535 $Y=3.33
+ $X2=8.45 $Y2=3.33
r229 107 109 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.535 $Y=3.33
+ $X2=8.88 $Y2=3.33
r230 105 106 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r231 103 106 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r232 102 105 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r233 102 103 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r234 100 139 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=7.17 $Y=3.33
+ $X2=7.345 $Y2=3.33
r235 100 105 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.17 $Y=3.33
+ $X2=6.96 $Y2=3.33
r236 99 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r237 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r238 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r239 96 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r240 95 98 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r241 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r242 93 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.26 $Y2=3.33
r243 93 95 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.6 $Y2=3.33
r244 92 137 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r245 92 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r246 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r247 89 132 11.3727 $w=1.7e-07 $l=4.75e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.09 $Y2=3.33
r248 89 91 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.68 $Y2=3.33
r249 88 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=3.26 $Y2=3.33
r250 88 91 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=1.68 $Y2=3.33
r251 86 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r252 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r253 83 132 11.3727 $w=1.7e-07 $l=4.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.09 $Y2=3.33
r254 83 85 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r255 81 143 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r256 81 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r257 81 139 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r258 79 112 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=10.465 $Y=3.33
+ $X2=10.32 $Y2=3.33
r259 79 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.465 $Y=3.33
+ $X2=10.63 $Y2=3.33
r260 78 116 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=10.795 $Y=3.33
+ $X2=11.28 $Y2=3.33
r261 78 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.795 $Y=3.33
+ $X2=10.63 $Y2=3.33
r262 76 98 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.56 $Y2=3.33
r263 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.87 $Y2=3.33
r264 75 102 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r265 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.87 $Y2=3.33
r266 71 154 3.07266 $w=2.95e-07 $l=1.1025e-07 $layer=LI1_cond $X=14.617 $Y=3.245
+ $X2=14.675 $Y2=3.33
r267 71 73 37.8939 $w=2.93e-07 $l=9.7e-07 $layer=LI1_cond $X=14.617 $Y=3.245
+ $X2=14.617 $Y2=2.275
r268 67 151 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.74 $Y=3.245
+ $X2=13.74 $Y2=3.33
r269 67 69 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=13.74 $Y=3.245
+ $X2=13.74 $Y2=2.275
r270 66 148 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.885 $Y=3.33
+ $X2=12.76 $Y2=3.33
r271 65 151 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.615 $Y=3.33
+ $X2=13.74 $Y2=3.33
r272 65 66 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=13.615 $Y=3.33
+ $X2=12.885 $Y2=3.33
r273 61 64 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=12.76 $Y=1.985
+ $X2=12.76 $Y2=2.815
r274 59 148 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.76 $Y=3.245
+ $X2=12.76 $Y2=3.33
r275 59 64 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.76 $Y=3.245
+ $X2=12.76 $Y2=2.815
r276 55 145 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.775 $Y=3.245
+ $X2=11.775 $Y2=3.33
r277 55 57 58.0831 $w=2.48e-07 $l=1.26e-06 $layer=LI1_cond $X=11.775 $Y=3.245
+ $X2=11.775 $Y2=1.985
r278 51 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.63 $Y=3.245
+ $X2=10.63 $Y2=3.33
r279 51 53 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.63 $Y=3.245
+ $X2=10.63 $Y2=2.75
r280 47 50 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.45 $Y=1.91
+ $X2=8.45 $Y2=2.59
r281 45 142 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.45 $Y=3.245
+ $X2=8.45 $Y2=3.33
r282 45 50 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=8.45 $Y=3.245
+ $X2=8.45 $Y2=2.59
r283 44 139 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=7.52 $Y=3.33
+ $X2=7.345 $Y2=3.33
r284 43 142 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.365 $Y=3.33
+ $X2=8.45 $Y2=3.33
r285 43 44 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=8.365 $Y=3.33
+ $X2=7.52 $Y2=3.33
r286 39 139 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.345 $Y=3.245
+ $X2=7.345 $Y2=3.33
r287 39 41 13.8293 $w=3.48e-07 $l=4.2e-07 $layer=LI1_cond $X=7.345 $Y=3.245
+ $X2=7.345 $Y2=2.825
r288 35 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=3.33
r289 35 37 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=2.835
r290 31 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=3.33
r291 31 33 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=2.79
r292 10 73 300 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_PDIFF $count=2 $X=14.45
+ $Y=1.84 $X2=14.6 $Y2=2.275
r293 9 69 300 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_PDIFF $count=2 $X=13.55
+ $Y=1.84 $X2=13.7 $Y2=2.275
r294 8 64 600 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=12.565
+ $Y=1.84 $X2=12.8 $Y2=2.815
r295 8 61 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=12.565
+ $Y=1.84 $X2=12.8 $Y2=1.985
r296 7 57 300 $w=1.7e-07 $l=6.74611e-07 $layer=licon1_PDIFF $count=2 $X=11.55
+ $Y=2.54 $X2=11.815 $Y2=1.985
r297 6 53 600 $w=1.7e-07 $l=3.91152e-07 $layer=licon1_PDIFF $count=1 $X=10.33
+ $Y=2.54 $X2=10.63 $Y2=2.75
r298 5 50 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.735 $X2=8.45 $Y2=2.59
r299 5 47 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.735 $X2=8.45 $Y2=1.91
r300 4 41 600 $w=1.7e-07 $l=6.20524e-07 $layer=licon1_PDIFF $count=1 $X=7.1
+ $Y=2.315 $X2=7.345 $Y2=2.825
r301 3 37 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=1.96 $X2=4.87 $Y2=2.835
r302 2 33 600 $w=1.7e-07 $l=5.39815e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=2.32 $X2=3.26 $Y2=2.79
r303 1 129 150 $w=1.7e-07 $l=8.8955e-07 $layer=licon1_PDIFF $count=4 $X=0.58
+ $Y=2.32 $X2=1.4 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%A_415_81# 1 2 3 4 5 18 22 24 27 32 36 39 40
+ 41 42 43 45 47 55 56 57
c158 57 0 4.7366e-20 $X=4.645 $Y=2.5
c159 45 0 4.8605e-20 $X=6.46 $Y=2.085
c160 42 0 1.2914e-19 $X=6.375 $Y=2.17
c161 40 0 1.54393e-19 $X=6.375 $Y=1.33
c162 32 0 7.67579e-20 $X=5.745 $Y=2.495
c163 27 0 1.19423e-19 $X=3.53 $Y=2.33
r164 56 57 4.00505 $w=1.78e-07 $l=6.5e-08 $layer=LI1_cond $X=4.58 $Y=2.5
+ $X2=4.645 $Y2=2.5
r165 54 55 0.976 $w=5e-07 $l=4e-08 $layer=LI1_cond $X=3.72 $Y=2.465 $X2=3.72
+ $Y2=2.505
r166 52 54 0.854 $w=5e-07 $l=3.5e-08 $layer=LI1_cond $X=3.72 $Y=2.43 $X2=3.72
+ $Y2=2.465
r167 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.46 $Y=1.415
+ $X2=6.46 $Y2=2.085
r168 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.375 $Y=2.17
+ $X2=6.46 $Y2=2.085
r169 42 43 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.375 $Y=2.17
+ $X2=6.075 $Y2=2.17
r170 40 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.375 $Y=1.33
+ $X2=6.46 $Y2=1.415
r171 40 41 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.375 $Y=1.33
+ $X2=5.99 $Y2=1.33
r172 39 59 3.26369 $w=2.5e-07 $l=1.90955e-07 $layer=LI1_cond $X=5.95 $Y=2.41
+ $X2=5.91 $Y2=2.582
r173 38 43 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.95 $Y=2.255
+ $X2=6.075 $Y2=2.17
r174 38 39 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=5.95 $Y=2.255
+ $X2=5.95 $Y2=2.41
r175 34 41 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.89 $Y=1.245
+ $X2=5.99 $Y2=1.33
r176 34 36 19.1318 $w=1.98e-07 $l=3.45e-07 $layer=LI1_cond $X=5.89 $Y=1.245
+ $X2=5.89 $Y2=0.9
r177 32 59 3.87948 $w=1.7e-07 $l=2.03912e-07 $layer=LI1_cond $X=5.745 $Y=2.495
+ $X2=5.91 $Y2=2.582
r178 32 57 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=5.745 $Y=2.495
+ $X2=4.645 $Y2=2.495
r179 31 55 7.15667 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.995 $Y=2.505
+ $X2=3.72 $Y2=2.505
r180 31 56 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.995 $Y=2.505
+ $X2=4.58 $Y2=2.505
r181 27 52 8.12146 $w=5e-07 $l=2.34734e-07 $layer=LI1_cond $X=3.53 $Y=2.33
+ $X2=3.72 $Y2=2.43
r182 26 27 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.53 $Y=1.09
+ $X2=3.53 $Y2=2.33
r183 25 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=1.005
+ $X2=2.65 $Y2=1.005
r184 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=3.53 $Y2=1.09
r185 24 25 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=2.735 $Y2=1.005
r186 23 47 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.435 $Y=2.43
+ $X2=2.27 $Y2=2.43
r187 22 52 7.15667 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=3.72 $Y2=2.43
r188 22 23 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=2.435 $Y2=2.43
r189 18 50 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.65 $Y=0.72
+ $X2=2.65 $Y2=1.005
r190 18 20 2.99635 $w=2.48e-07 $l=6.5e-08 $layer=LI1_cond $X=2.565 $Y=0.72
+ $X2=2.5 $Y2=0.72
r191 5 59 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.765
+ $Y=2.315 $X2=5.91 $Y2=2.525
r192 4 54 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.68
+ $Y=2.32 $X2=3.83 $Y2=2.465
r193 3 47 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.12
+ $Y=2.32 $X2=2.27 $Y2=2.465
r194 2 36 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.765
+ $Y=0.69 $X2=5.89 $Y2=0.9
r195 1 20 182 $w=1.7e-07 $l=5.45436e-07 $layer=licon1_NDIFF $count=1 $X=2.075
+ $Y=0.405 $X2=2.5 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%Q 1 2 3 4 15 17 18 21 25 26 29 35 38 40
c67 40 0 1.4738e-19 $X=14.64 $Y=1.665
c68 26 0 1.81891e-19 $X=13.415 $Y=1.855
c69 15 0 1.86508e-19 $X=12.7 $Y=0.515
r70 42 43 0.0389776 $w=6.26e-07 $l=2e-09 $layer=LI1_cond $X=14.17 $Y=1.62
+ $X2=14.172 $Y2=1.62
r71 40 43 9.12077 $w=6.26e-07 $l=4.68e-07 $layer=LI1_cond $X=14.64 $Y=1.62
+ $X2=14.172 $Y2=1.62
r72 38 42 8.59112 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=14.17 $Y=1.3
+ $X2=14.17 $Y2=1.62
r73 37 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.17 $Y=1.1
+ $X2=14.17 $Y2=1.015
r74 37 38 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=14.17 $Y=1.1 $X2=14.17
+ $Y2=1.3
r75 33 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.17 $Y=0.93
+ $X2=14.17 $Y2=1.015
r76 33 35 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=14.17 $Y=0.93
+ $X2=14.17 $Y2=0.515
r77 29 31 44.4897 $w=2.13e-07 $l=8.3e-07 $layer=LI1_cond $X=14.172 $Y=1.985
+ $X2=14.172 $Y2=2.815
r78 27 43 7.10307 $w=2.15e-07 $l=3.2e-07 $layer=LI1_cond $X=14.172 $Y=1.94
+ $X2=14.172 $Y2=1.62
r79 27 29 2.41209 $w=2.13e-07 $l=4.5e-08 $layer=LI1_cond $X=14.172 $Y=1.94
+ $X2=14.172 $Y2=1.985
r80 25 42 9.36281 $w=6.26e-07 $l=2.82666e-07 $layer=LI1_cond $X=14.065 $Y=1.855
+ $X2=14.17 $Y2=1.62
r81 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=14.065 $Y=1.855
+ $X2=13.415 $Y2=1.855
r82 21 23 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=13.25 $Y=1.985
+ $X2=13.25 $Y2=2.815
r83 19 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.25 $Y=1.94
+ $X2=13.415 $Y2=1.855
r84 19 21 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=13.25 $Y=1.94
+ $X2=13.25 $Y2=1.985
r85 17 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.085 $Y=1.015
+ $X2=14.17 $Y2=1.015
r86 17 18 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=14.085 $Y=1.015
+ $X2=12.865 $Y2=1.015
r87 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.7 $Y=0.93
+ $X2=12.865 $Y2=1.015
r88 13 15 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=12.7 $Y=0.93
+ $X2=12.7 $Y2=0.515
r89 4 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=14
+ $Y=1.84 $X2=14.15 $Y2=2.815
r90 4 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=14
+ $Y=1.84 $X2=14.15 $Y2=1.985
r91 3 23 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.1
+ $Y=1.84 $X2=13.25 $Y2=2.815
r92 3 21 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.1
+ $Y=1.84 $X2=13.25 $Y2=1.985
r93 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.03
+ $Y=0.37 $X2=14.17 $Y2=0.515
r94 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.56
+ $Y=0.37 $X2=12.7 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%VGND 1 2 3 4 5 6 7 8 27 31 35 37 41 45 47
+ 49 52 53 54 56 68 72 80 93 99 102 106 112 115 120 126 129
c145 129 0 3.56444e-20 $X=14.64 $Y=0
c146 49 0 2.76177e-20 $X=14.6 $Y=0.515
r147 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r148 125 126 11.7074 $w=8.43e-07 $l=1.65e-07 $layer=LI1_cond $X=13.74 $Y=0.337
+ $X2=13.905 $Y2=0.337
r149 122 125 0.849286 $w=8.43e-07 $l=6e-08 $layer=LI1_cond $X=13.68 $Y=0.337
+ $X2=13.74 $Y2=0.337
r150 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r151 119 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r152 118 122 6.79429 $w=8.43e-07 $l=4.8e-07 $layer=LI1_cond $X=13.2 $Y=0.337
+ $X2=13.68 $Y2=0.337
r153 118 120 11.7074 $w=8.43e-07 $l=1.65e-07 $layer=LI1_cond $X=13.2 $Y=0.337
+ $X2=13.035 $Y2=0.337
r154 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r155 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r156 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r157 106 109 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.595 $Y2=0.325
r158 102 103 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r159 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r160 97 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r161 97 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=13.68 $Y2=0
r162 96 126 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=14.16 $Y=0
+ $X2=13.905 $Y2=0
r163 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r164 93 128 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=14.435 $Y=0
+ $X2=14.657 $Y2=0
r165 93 96 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=14.435 $Y=0
+ $X2=14.16 $Y2=0
r166 92 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r167 92 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r168 91 120 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.72 $Y=0
+ $X2=13.035 $Y2=0
r169 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r170 89 115 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.365 $Y=0
+ $X2=12.235 $Y2=0
r171 89 91 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=12.365 $Y=0
+ $X2=12.72 $Y2=0
r172 87 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r173 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r174 84 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.76 $Y2=0
r175 84 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r176 83 86 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=10.8 $Y=0 $X2=11.76
+ $Y2=0
r177 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r178 81 112 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=10.58 $Y=0
+ $X2=10.36 $Y2=0
r179 81 83 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=10.58 $Y=0 $X2=10.8
+ $Y2=0
r180 80 115 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.105 $Y=0
+ $X2=12.235 $Y2=0
r181 80 86 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.105 $Y=0
+ $X2=11.76 $Y2=0
r182 79 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r183 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r184 76 79 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=9.84 $Y2=0
r185 75 78 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=0 $X2=9.84
+ $Y2=0
r186 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r187 73 106 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.76 $Y=0
+ $X2=7.595 $Y2=0
r188 73 75 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.76 $Y=0 $X2=7.92
+ $Y2=0
r189 72 112 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=10.14 $Y=0
+ $X2=10.36 $Y2=0
r190 72 78 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=10.14 $Y=0 $X2=9.84
+ $Y2=0
r191 71 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r192 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r193 68 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=0
+ $X2=4.88 $Y2=0
r194 68 70 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.715 $Y=0
+ $X2=4.56 $Y2=0
r195 67 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r196 66 67 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r197 64 67 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r198 64 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r199 63 66 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r200 63 64 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r201 61 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r202 61 63 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r203 59 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r204 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r205 56 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r206 56 58 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r207 54 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r208 54 103 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=5.04 $Y2=0
r209 54 106 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r210 52 66 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.6
+ $Y2=0
r211 52 53 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.832
+ $Y2=0
r212 51 70 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=4.56
+ $Y2=0
r213 51 53 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=3.832
+ $Y2=0
r214 47 128 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=14.6 $Y=0.085
+ $X2=14.657 $Y2=0
r215 47 49 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=14.6 $Y=0.085
+ $X2=14.6 $Y2=0.515
r216 43 115 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=12.235 $Y=0.085
+ $X2=12.235 $Y2=0
r217 43 45 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=12.235 $Y=0.085
+ $X2=12.235 $Y2=0.515
r218 39 112 1.73497 $w=4.4e-07 $l=8.5e-08 $layer=LI1_cond $X=10.36 $Y=0.085
+ $X2=10.36 $Y2=0
r219 39 41 11.2625 $w=4.38e-07 $l=4.3e-07 $layer=LI1_cond $X=10.36 $Y=0.085
+ $X2=10.36 $Y2=0.515
r220 38 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=0
+ $X2=4.88 $Y2=0
r221 37 106 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.43 $Y=0
+ $X2=7.595 $Y2=0
r222 37 38 155.599 $w=1.68e-07 $l=2.385e-06 $layer=LI1_cond $X=7.43 $Y=0
+ $X2=5.045 $Y2=0
r223 33 102 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0
r224 33 35 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0.665
r225 29 53 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.832 $Y=0.085
+ $X2=3.832 $Y2=0
r226 29 31 17.7299 $w=3.23e-07 $l=5e-07 $layer=LI1_cond $X=3.832 $Y=0.085
+ $X2=3.832 $Y2=0.585
r227 25 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r228 25 27 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.555
r229 8 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.46
+ $Y=0.37 $X2=14.6 $Y2=0.515
r230 7 125 91 $w=1.7e-07 $l=8.55132e-07 $layer=licon1_NDIFF $count=2 $X=12.99
+ $Y=0.37 $X2=13.74 $Y2=0.595
r231 6 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.13
+ $Y=0.37 $X2=12.27 $Y2=0.515
r232 5 41 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=10.165
+ $Y=0.37 $X2=10.36 $Y2=0.515
r233 4 109 182 $w=1.7e-07 $l=4.62088e-07 $layer=licon1_NDIFF $count=1 $X=7.375
+ $Y=0.69 $X2=7.595 $Y2=0.325
r234 3 35 182 $w=1.7e-07 $l=2.32379e-07 $layer=licon1_NDIFF $count=1 $X=4.68
+ $Y=0.595 $X2=4.88 $Y2=0.665
r235 2 31 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.65
+ $Y=0.405 $X2=3.79 $Y2=0.585
r236 1 27 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LS__SDFRTP_4%noxref_24 1 2 7 11 13
r27 13 16 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.27 $Y=0.34
+ $X2=1.27 $Y2=0.55
r28 9 11 6.70512 $w=2.73e-07 $l=1.6e-07 $layer=LI1_cond $X=3.362 $Y=0.425
+ $X2=3.362 $Y2=0.585
r29 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=0.34
+ $X2=1.27 $Y2=0.34
r30 7 9 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=3.225 $Y=0.34
+ $X2=3.362 $Y2=0.425
r31 7 8 116.781 $w=1.68e-07 $l=1.79e-06 $layer=LI1_cond $X=3.225 $Y=0.34
+ $X2=1.435 $Y2=0.34
r32 2 11 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.22 $Y=0.405
+ $X2=3.36 $Y2=0.585
r33 1 16 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.405 $X2=1.27 $Y2=0.55
.ends

