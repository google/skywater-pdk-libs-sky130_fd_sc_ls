* File: sky130_fd_sc_ls__fa_4.pxi.spice
* Created: Fri Aug 28 13:25:31 2020
* 
x_PM_SKY130_FD_SC_LS__FA_4%B N_B_c_204_n N_B_M1010_g N_B_M1026_g N_B_M1023_g
+ N_B_c_195_n N_B_M1000_g N_B_M1030_g N_B_c_197_n N_B_M1003_g N_B_c_198_n
+ N_B_M1011_g N_B_M1037_g N_B_c_200_n N_B_c_201_n N_B_c_209_n N_B_c_222_p
+ N_B_c_281_p N_B_c_202_n N_B_c_226_p N_B_c_211_n N_B_c_305_p N_B_c_212_n B B
+ PM_SKY130_FD_SC_LS__FA_4%B
x_PM_SKY130_FD_SC_LS__FA_4%CIN N_CIN_c_419_n N_CIN_M1038_g N_CIN_c_420_n
+ N_CIN_M1029_g N_CIN_M1027_g N_CIN_c_422_n N_CIN_M1005_g N_CIN_c_423_n
+ N_CIN_M1017_g N_CIN_c_424_n N_CIN_M1025_g N_CIN_c_425_n N_CIN_c_426_n
+ N_CIN_c_427_n N_CIN_c_428_n N_CIN_c_429_n N_CIN_c_430_n N_CIN_c_431_n CIN
+ N_CIN_c_432_n N_CIN_c_433_n PM_SKY130_FD_SC_LS__FA_4%CIN
x_PM_SKY130_FD_SC_LS__FA_4%A_418_74# N_A_418_74#_M1038_d N_A_418_74#_M1029_d
+ N_A_418_74#_c_570_n N_A_418_74#_M1016_g N_A_418_74#_c_571_n
+ N_A_418_74#_M1006_g N_A_418_74#_c_585_n N_A_418_74#_M1008_g
+ N_A_418_74#_M1013_g N_A_418_74#_c_586_n N_A_418_74#_M1009_g
+ N_A_418_74#_M1014_g N_A_418_74#_c_587_n N_A_418_74#_M1018_g
+ N_A_418_74#_M1022_g N_A_418_74#_c_588_n N_A_418_74#_M1019_g
+ N_A_418_74#_M1035_g N_A_418_74#_c_576_n N_A_418_74#_c_669_p
+ N_A_418_74#_c_599_n N_A_418_74#_c_602_n N_A_418_74#_c_604_n
+ N_A_418_74#_c_638_n N_A_418_74#_c_577_n N_A_418_74#_c_606_n
+ N_A_418_74#_c_644_n N_A_418_74#_c_578_n N_A_418_74#_c_579_n
+ N_A_418_74#_c_613_n N_A_418_74#_c_683_p N_A_418_74#_c_614_n
+ N_A_418_74#_c_580_n N_A_418_74#_c_581_n N_A_418_74#_c_764_p
+ N_A_418_74#_c_615_n N_A_418_74#_c_619_n N_A_418_74#_c_622_n
+ N_A_418_74#_c_647_n N_A_418_74#_c_590_n N_A_418_74#_c_626_n
+ N_A_418_74#_c_629_n N_A_418_74#_c_582_n N_A_418_74#_c_583_n
+ PM_SKY130_FD_SC_LS__FA_4%A_418_74#
x_PM_SKY130_FD_SC_LS__FA_4%A N_A_c_863_n N_A_M1032_g N_A_c_876_n N_A_M1028_g
+ N_A_c_878_n N_A_c_879_n N_A_c_865_n N_A_c_866_n N_A_c_881_n N_A_c_882_n
+ N_A_c_883_n N_A_M1001_g N_A_M1033_g N_A_c_885_n N_A_M1015_g N_A_c_867_n
+ N_A_c_868_n N_A_c_887_n N_A_c_888_n N_A_c_889_n N_A_M1004_g N_A_c_891_n
+ N_A_M1039_g N_A_c_870_n N_A_M1012_g N_A_c_871_n N_A_c_895_n N_A_c_872_n
+ N_A_c_896_n N_A_c_897_n A A N_A_c_874_n PM_SKY130_FD_SC_LS__FA_4%A
x_PM_SKY130_FD_SC_LS__FA_4%A_1024_74# N_A_1024_74#_M1016_d N_A_1024_74#_M1006_d
+ N_A_1024_74#_c_1072_n N_A_1024_74#_M1002_g N_A_1024_74#_M1020_g
+ N_A_1024_74#_c_1073_n N_A_1024_74#_M1007_g N_A_1024_74#_M1021_g
+ N_A_1024_74#_c_1074_n N_A_1024_74#_M1024_g N_A_1024_74#_M1034_g
+ N_A_1024_74#_c_1075_n N_A_1024_74#_M1031_g N_A_1024_74#_M1036_g
+ N_A_1024_74#_c_1081_n N_A_1024_74#_c_1084_n N_A_1024_74#_c_1087_n
+ N_A_1024_74#_c_1068_n N_A_1024_74#_c_1076_n N_A_1024_74#_c_1069_n
+ N_A_1024_74#_c_1078_n N_A_1024_74#_c_1092_n N_A_1024_74#_c_1104_n
+ N_A_1024_74#_c_1093_n N_A_1024_74#_c_1095_n N_A_1024_74#_c_1070_n
+ N_A_1024_74#_c_1071_n PM_SKY130_FD_SC_LS__FA_4%A_1024_74#
x_PM_SKY130_FD_SC_LS__FA_4%A_27_392# N_A_27_392#_M1028_s N_A_27_392#_M1010_d
+ N_A_27_392#_c_1223_n N_A_27_392#_c_1224_n N_A_27_392#_c_1232_n
+ N_A_27_392#_c_1233_n N_A_27_392#_c_1225_n N_A_27_392#_c_1226_n
+ PM_SKY130_FD_SC_LS__FA_4%A_27_392#
x_PM_SKY130_FD_SC_LS__FA_4%VPWR N_VPWR_M1028_d N_VPWR_M1001_d N_VPWR_M1003_d
+ N_VPWR_M1012_d N_VPWR_M1007_s N_VPWR_M1031_s N_VPWR_M1009_d N_VPWR_M1019_d
+ N_VPWR_c_1275_n N_VPWR_c_1276_n N_VPWR_c_1277_n N_VPWR_c_1278_n
+ N_VPWR_c_1279_n N_VPWR_c_1280_n N_VPWR_c_1281_n N_VPWR_c_1282_n
+ N_VPWR_c_1283_n N_VPWR_c_1284_n N_VPWR_c_1285_n VPWR N_VPWR_c_1286_n
+ N_VPWR_c_1287_n N_VPWR_c_1288_n N_VPWR_c_1289_n N_VPWR_c_1290_n
+ N_VPWR_c_1291_n N_VPWR_c_1292_n N_VPWR_c_1293_n N_VPWR_c_1294_n
+ N_VPWR_c_1295_n N_VPWR_c_1296_n N_VPWR_c_1297_n N_VPWR_c_1274_n
+ PM_SKY130_FD_SC_LS__FA_4%VPWR
x_PM_SKY130_FD_SC_LS__FA_4%A_737_347# N_A_737_347#_M1005_d N_A_737_347#_M1004_d
+ N_A_737_347#_c_1431_n N_A_737_347#_c_1434_n N_A_737_347#_c_1427_n
+ N_A_737_347#_c_1428_n PM_SKY130_FD_SC_LS__FA_4%A_737_347#
x_PM_SKY130_FD_SC_LS__FA_4%SUM N_SUM_M1020_s N_SUM_M1034_s N_SUM_M1002_d
+ N_SUM_M1024_d N_SUM_c_1466_n N_SUM_c_1467_n N_SUM_c_1463_n N_SUM_c_1494_n
+ N_SUM_c_1464_n N_SUM_c_1465_n SUM SUM SUM SUM PM_SKY130_FD_SC_LS__FA_4%SUM
x_PM_SKY130_FD_SC_LS__FA_4%COUT N_COUT_M1013_d N_COUT_M1022_d N_COUT_M1008_s
+ N_COUT_M1018_s N_COUT_c_1530_n N_COUT_c_1531_n N_COUT_c_1526_n N_COUT_c_1532_n
+ N_COUT_c_1548_n N_COUT_c_1527_n N_COUT_c_1528_n N_COUT_c_1529_n
+ N_COUT_c_1563_n COUT COUT COUT COUT N_COUT_c_1533_n COUT
+ PM_SKY130_FD_SC_LS__FA_4%COUT
x_PM_SKY130_FD_SC_LS__FA_4%A_27_74# N_A_27_74#_M1032_s N_A_27_74#_M1026_d
+ N_A_27_74#_c_1595_n N_A_27_74#_c_1596_n N_A_27_74#_c_1599_n
+ N_A_27_74#_c_1597_n PM_SKY130_FD_SC_LS__FA_4%A_27_74#
x_PM_SKY130_FD_SC_LS__FA_4%VGND N_VGND_M1032_d N_VGND_M1033_d N_VGND_M1030_d
+ N_VGND_M1039_d N_VGND_M1021_d N_VGND_M1036_d N_VGND_M1014_s N_VGND_M1035_s
+ N_VGND_c_1627_n N_VGND_c_1628_n N_VGND_c_1629_n N_VGND_c_1630_n
+ N_VGND_c_1631_n N_VGND_c_1632_n N_VGND_c_1633_n N_VGND_c_1634_n VGND
+ N_VGND_c_1635_n N_VGND_c_1636_n N_VGND_c_1637_n N_VGND_c_1638_n
+ N_VGND_c_1639_n N_VGND_c_1640_n N_VGND_c_1641_n N_VGND_c_1642_n
+ N_VGND_c_1643_n N_VGND_c_1644_n N_VGND_c_1645_n N_VGND_c_1646_n
+ PM_SKY130_FD_SC_LS__FA_4%VGND
x_PM_SKY130_FD_SC_LS__FA_4%A_734_74# N_A_734_74#_M1027_d N_A_734_74#_M1015_d
+ N_A_734_74#_c_1776_n N_A_734_74#_c_1774_n N_A_734_74#_c_1775_n
+ PM_SKY130_FD_SC_LS__FA_4%A_734_74#
cc_1 VNB N_B_M1026_g 0.0209127f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=0.74
cc_2 VNB N_B_M1023_g 0.0210869f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.74
cc_3 VNB N_B_c_195_n 0.0248541f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.66
cc_4 VNB N_B_M1030_g 0.0203825f $X=-0.19 $Y=-0.245 $X2=4.025 $Y2=0.74
cc_5 VNB N_B_c_197_n 0.0265492f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=1.66
cc_6 VNB N_B_c_198_n 0.0217205f $X=-0.19 $Y=-0.245 $X2=6.1 $Y2=1.66
cc_7 VNB N_B_M1037_g 0.0183203f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=0.74
cc_8 VNB N_B_c_200_n 0.00309095f $X=-0.19 $Y=-0.245 $X2=1.665 $Y2=1.417
cc_9 VNB N_B_c_201_n 0.0397216f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.41
cc_10 VNB N_B_c_202_n 8.09421e-19 $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.41
cc_11 VNB B 0.00826485f $X=-0.19 $Y=-0.245 $X2=6.395 $Y2=1.58
cc_12 VNB N_CIN_c_419_n 0.018815f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.66
cc_13 VNB N_CIN_c_420_n 0.0309653f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=1.245
cc_14 VNB N_CIN_M1027_g 0.019466f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.74
cc_15 VNB N_CIN_c_422_n 0.0232802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_CIN_c_423_n 0.0296271f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=2.235
cc_17 VNB N_CIN_c_424_n 0.0178512f $X=-0.19 $Y=-0.245 $X2=4.025 $Y2=0.74
cc_18 VNB N_CIN_c_425_n 0.0025906f $X=-0.19 $Y=-0.245 $X2=6.1 $Y2=1.66
cc_19 VNB N_CIN_c_426_n 0.0071807f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=1.245
cc_20 VNB N_CIN_c_427_n 0.00290723f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=0.74
cc_21 VNB N_CIN_c_428_n 0.018935f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=0.74
cc_22 VNB N_CIN_c_429_n 0.00298431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_CIN_c_430_n 0.00460694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_CIN_c_431_n 0.00274216f $X=-0.19 $Y=-0.245 $X2=1.75 $Y2=1.575
cc_25 VNB N_CIN_c_432_n 0.00310764f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.41
cc_26 VNB N_CIN_c_433_n 0.00361772f $X=-0.19 $Y=-0.245 $X2=6.395 $Y2=1.58
cc_27 VNB N_A_418_74#_c_570_n 0.0177385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_418_74#_c_571_n 0.0279921f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.74
cc_29 VNB N_A_418_74#_M1013_g 0.0209667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_418_74#_M1014_g 0.0185701f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=1.245
cc_31 VNB N_A_418_74#_M1022_g 0.0182888f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.41
cc_32 VNB N_A_418_74#_M1035_g 0.0251724f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.41
cc_33 VNB N_A_418_74#_c_576_n 0.00500716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_418_74#_c_577_n 0.00333942f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.817
cc_35 VNB N_A_418_74#_c_578_n 0.00802253f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=1.452
cc_36 VNB N_A_418_74#_c_579_n 9.82756e-19 $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.41
cc_37 VNB N_A_418_74#_c_580_n 0.00296963f $X=-0.19 $Y=-0.245 $X2=5.915 $Y2=1.805
cc_38 VNB N_A_418_74#_c_581_n 0.00392926f $X=-0.19 $Y=-0.245 $X2=6 $Y2=1.575
cc_39 VNB N_A_418_74#_c_582_n 0.00879717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_418_74#_c_583_n 0.120757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_c_863_n 0.00564717f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=2.235
cc_42 VNB N_A_M1032_g 0.0277073f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=0.74
cc_43 VNB N_A_c_865_n 0.00506139f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=2.235
cc_44 VNB N_A_c_866_n 0.0110176f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=2.235
cc_45 VNB N_A_c_867_n 0.00548129f $X=-0.19 $Y=-0.245 $X2=1.665 $Y2=1.417
cc_46 VNB N_A_c_868_n 0.0140582f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.417
cc_47 VNB N_A_M1039_g 0.0403652f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.41
cc_48 VNB N_A_c_870_n 0.0024482f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=1.83
cc_49 VNB N_A_c_871_n 0.0161869f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.41
cc_50 VNB N_A_c_872_n 0.0169826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB A 0.0194965f $X=-0.19 $Y=-0.245 $X2=6.395 $Y2=1.58
cc_52 VNB N_A_c_874_n 0.0599859f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.41
cc_53 VNB N_A_1024_74#_M1020_g 0.0221413f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.66
cc_54 VNB N_A_1024_74#_M1021_g 0.0217363f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=1.66
cc_55 VNB N_A_1024_74#_M1034_g 0.0210584f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=0.74
cc_56 VNB N_A_1024_74#_M1036_g 0.0220203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1024_74#_c_1068_n 0.00361783f $X=-0.19 $Y=-0.245 $X2=4.115
+ $Y2=1.41
cc_58 VNB N_A_1024_74#_c_1069_n 3.03738e-19 $X=-0.19 $Y=-0.245 $X2=5.915
+ $Y2=1.58
cc_59 VNB N_A_1024_74#_c_1070_n 0.0029978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1024_74#_c_1071_n 0.0830321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VPWR_c_1274_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_SUM_c_1463_n 0.00586669f $X=-0.19 $Y=-0.245 $X2=4.025 $Y2=0.74
cc_63 VNB N_SUM_c_1464_n 0.00234369f $X=-0.19 $Y=-0.245 $X2=6.1 $Y2=2.235
cc_64 VNB N_SUM_c_1465_n 0.00137885f $X=-0.19 $Y=-0.245 $X2=6.1 $Y2=2.235
cc_65 VNB N_COUT_c_1526_n 0.00220089f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=1.66
cc_66 VNB N_COUT_c_1527_n 0.00123375f $X=-0.19 $Y=-0.245 $X2=6.1 $Y2=2.235
cc_67 VNB N_COUT_c_1528_n 0.00229206f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=0.74
cc_68 VNB N_COUT_c_1529_n 0.00154258f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.417
cc_69 VNB N_A_27_74#_c_1595_n 0.00249128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_27_74#_c_1596_n 0.0306363f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=2.235
cc_71 VNB N_A_27_74#_c_1597_n 0.00162437f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=1.66
cc_72 VNB N_VGND_c_1627_n 0.00574325f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=0.74
cc_73 VNB N_VGND_c_1628_n 0.00546039f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.41
cc_74 VNB N_VGND_c_1629_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1630_n 0.0471419f $X=-0.19 $Y=-0.245 $X2=1.75 $Y2=1.95
cc_76 VNB N_VGND_c_1631_n 0.0556692f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.745
cc_77 VNB N_VGND_c_1632_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.41
cc_78 VNB N_VGND_c_1633_n 0.0133472f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.41
cc_79 VNB N_VGND_c_1634_n 0.0178103f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.41
cc_80 VNB N_VGND_c_1635_n 0.0547728f $X=-0.19 $Y=-0.245 $X2=6.175 $Y2=1.41
cc_81 VNB N_VGND_c_1636_n 0.0185379f $X=-0.19 $Y=-0.245 $X2=6.175 $Y2=1.575
cc_82 VNB N_VGND_c_1637_n 0.0185379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1638_n 0.0175388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1639_n 0.0174844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1640_n 0.0185699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1641_n 0.01914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1642_n 0.0153962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1643_n 0.0170767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1644_n 0.015362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1645_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1646_n 0.579257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_734_74#_c_1774_n 0.00205545f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.74
cc_93 VNB N_A_734_74#_c_1775_n 0.00203932f $X=-0.19 $Y=-0.245 $X2=4.025
+ $Y2=1.245
cc_94 VPB N_B_c_204_n 0.0144816f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.66
cc_95 VPB N_B_c_195_n 0.0237816f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.66
cc_96 VPB N_B_c_197_n 0.0242762f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=1.66
cc_97 VPB N_B_c_198_n 0.0242613f $X=-0.19 $Y=1.66 $X2=6.1 $Y2=1.66
cc_98 VPB N_B_c_201_n 0.0238543f $X=-0.19 $Y=1.66 $X2=1.51 $Y2=1.41
cc_99 VPB N_B_c_209_n 0.00260578f $X=-0.19 $Y=1.66 $X2=1.75 $Y2=1.95
cc_100 VPB N_B_c_202_n 0.00278934f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.41
cc_101 VPB N_B_c_211_n 0.00346695f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.41
cc_102 VPB N_B_c_212_n 0.00138677f $X=-0.19 $Y=1.66 $X2=4.62 $Y2=1.805
cc_103 VPB B 0.0115641f $X=-0.19 $Y=1.66 $X2=5.915 $Y2=1.58
cc_104 VPB B 0.00306973f $X=-0.19 $Y=1.66 $X2=6.395 $Y2=1.58
cc_105 VPB N_CIN_c_420_n 0.0211184f $X=-0.19 $Y=1.66 $X2=1.585 $Y2=1.245
cc_106 VPB N_CIN_c_422_n 0.024478f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_CIN_c_423_n 0.0210283f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=2.235
cc_108 VPB N_CIN_c_425_n 0.00192839f $X=-0.19 $Y=1.66 $X2=6.1 $Y2=1.66
cc_109 VPB N_CIN_c_432_n 0.00280188f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.41
cc_110 VPB N_CIN_c_433_n 4.02791e-19 $X=-0.19 $Y=1.66 $X2=6.395 $Y2=1.58
cc_111 VPB N_A_418_74#_c_571_n 0.021378f $X=-0.19 $Y=1.66 $X2=2.585 $Y2=0.74
cc_112 VPB N_A_418_74#_c_585_n 0.0161792f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=2.235
cc_113 VPB N_A_418_74#_c_586_n 0.0157671f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=2.235
cc_114 VPB N_A_418_74#_c_587_n 0.0157695f $X=-0.19 $Y=1.66 $X2=6.115 $Y2=0.74
cc_115 VPB N_A_418_74#_c_588_n 0.0174317f $X=-0.19 $Y=1.66 $X2=1.75 $Y2=1.575
cc_116 VPB N_A_418_74#_c_576_n 0.00121453f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_418_74#_c_590_n 0.00242081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_418_74#_c_583_n 0.0298035f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_c_863_n 0.00941817f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=2.235
cc_120 VPB N_A_c_876_n 0.00913453f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_M1028_g 0.0122398f $X=-0.19 $Y=1.66 $X2=2.585 $Y2=0.74
cc_122 VPB N_A_c_878_n 0.186653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_c_879_n 0.0188978f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.66
cc_124 VPB N_A_c_866_n 5.52855e-19 $X=-0.19 $Y=1.66 $X2=2.6 $Y2=2.235
cc_125 VPB N_A_c_881_n 0.00765451f $X=-0.19 $Y=1.66 $X2=4.025 $Y2=1.245
cc_126 VPB N_A_c_882_n 0.0165566f $X=-0.19 $Y=1.66 $X2=4.025 $Y2=0.74
cc_127 VPB N_A_c_883_n 0.00599309f $X=-0.19 $Y=1.66 $X2=4.025 $Y2=0.74
cc_128 VPB N_A_M1001_g 0.00836775f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=2.235
cc_129 VPB N_A_c_885_n 0.0926755f $X=-0.19 $Y=1.66 $X2=6.1 $Y2=2.235
cc_130 VPB N_A_c_868_n 8.14877e-19 $X=-0.19 $Y=1.66 $X2=1.51 $Y2=1.417
cc_131 VPB N_A_c_887_n 0.00746422f $X=-0.19 $Y=1.66 $X2=1.51 $Y2=1.41
cc_132 VPB N_A_c_888_n 0.0165566f $X=-0.19 $Y=1.66 $X2=1.51 $Y2=1.41
cc_133 VPB N_A_c_889_n 0.00635539f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_M1004_g 0.00842308f $X=-0.19 $Y=1.66 $X2=2.48 $Y2=2.035
cc_135 VPB N_A_c_891_n 0.149049f $X=-0.19 $Y=1.66 $X2=1.835 $Y2=2.035
cc_136 VPB N_A_M1039_g 0.00127901f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.41
cc_137 VPB N_A_c_870_n 0.00790577f $X=-0.19 $Y=1.66 $X2=3.95 $Y2=1.83
cc_138 VPB N_A_M1012_g 0.0102158f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.41
cc_139 VPB N_A_c_895_n 0.00879521f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.41
cc_140 VPB N_A_c_896_n 0.00879521f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.83
cc_141 VPB N_A_c_897_n 0.0297098f $X=-0.19 $Y=1.66 $X2=4.62 $Y2=1.805
cc_142 VPB A 0.0114344f $X=-0.19 $Y=1.66 $X2=6.395 $Y2=1.58
cc_143 VPB N_A_c_874_n 0.00515871f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.41
cc_144 VPB N_A_1024_74#_c_1072_n 0.0164592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_1024_74#_c_1073_n 0.0159404f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=2.235
cc_146 VPB N_A_1024_74#_c_1074_n 0.0159197f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=2.235
cc_147 VPB N_A_1024_74#_c_1075_n 0.0159594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_1024_74#_c_1076_n 0.00296107f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.41
cc_149 VPB N_A_1024_74#_c_1069_n 7.08103e-19 $X=-0.19 $Y=1.66 $X2=5.915 $Y2=1.58
cc_150 VPB N_A_1024_74#_c_1078_n 0.00275922f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_1024_74#_c_1071_n 0.0492224f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_27_392#_c_1223_n 0.0147058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_27_392#_c_1224_n 0.0302206f $X=-0.19 $Y=1.66 $X2=2.585 $Y2=0.74
cc_154 VPB N_A_27_392#_c_1225_n 0.00250926f $X=-0.19 $Y=1.66 $X2=4.025 $Y2=1.245
cc_155 VPB N_A_27_392#_c_1226_n 0.0103587f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=1.66
cc_156 VPB N_VPWR_c_1275_n 0.00542282f $X=-0.19 $Y=1.66 $X2=1.665 $Y2=1.417
cc_157 VPB N_VPWR_c_1276_n 0.00532455f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_1277_n 0.00573955f $X=-0.19 $Y=1.66 $X2=1.835 $Y2=2.035
cc_159 VPB N_VPWR_c_1278_n 0.0102422f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.41
cc_160 VPB N_VPWR_c_1279_n 0.00886117f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.41
cc_161 VPB N_VPWR_c_1280_n 0.0186447f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=2.035
cc_162 VPB N_VPWR_c_1281_n 0.00886117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1282_n 0.012247f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.452
cc_164 VPB N_VPWR_c_1283_n 0.0587025f $X=-0.19 $Y=1.66 $X2=1.585 $Y2=1.452
cc_165 VPB N_VPWR_c_1284_n 0.0634767f $X=-0.19 $Y=1.66 $X2=6.175 $Y2=1.41
cc_166 VPB N_VPWR_c_1285_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_1286_n 0.0175187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1287_n 0.0664038f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_1288_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1289_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1290_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1291_n 0.0195713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1292_n 0.0212973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1293_n 0.00530087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1294_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1295_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1296_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1297_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1274_n 0.0797771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_737_347#_c_1427_n 0.00275723f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=2.235
cc_181 VPB N_A_737_347#_c_1428_n 0.00243973f $X=-0.19 $Y=1.66 $X2=4.025 $Y2=0.74
cc_182 VPB N_SUM_c_1466_n 0.001142f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=2.235
cc_183 VPB N_SUM_c_1467_n 0.00257348f $X=-0.19 $Y=1.66 $X2=4.025 $Y2=1.245
cc_184 VPB N_SUM_c_1465_n 0.00160668f $X=-0.19 $Y=1.66 $X2=6.1 $Y2=2.235
cc_185 VPB SUM 0.00257348f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.745
cc_186 VPB N_COUT_c_1530_n 0.00183525f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=2.235
cc_187 VPB N_COUT_c_1531_n 0.00257348f $X=-0.19 $Y=1.66 $X2=4.025 $Y2=1.245
cc_188 VPB N_COUT_c_1532_n 0.00211023f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=2.235
cc_189 VPB N_COUT_c_1533_n 0.00202275f $X=-0.19 $Y=1.66 $X2=3.95 $Y2=1.83
cc_190 VPB COUT 0.00257348f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.745
cc_191 N_B_M1026_g N_CIN_c_419_n 0.0288887f $X=1.585 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_192 N_B_M1023_g N_CIN_c_419_n 0.0240859f $X=2.585 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_193 N_B_M1023_g N_CIN_c_420_n 0.00136863f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_194 N_B_c_195_n N_CIN_c_420_n 0.0592054f $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_195 N_B_c_200_n N_CIN_c_420_n 0.00227128f $X=1.665 $Y=1.417 $X2=0 $Y2=0
cc_196 N_B_c_201_n N_CIN_c_420_n 0.0149145f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B_c_209_n N_CIN_c_420_n 0.00492077f $X=1.75 $Y=1.95 $X2=0 $Y2=0
cc_198 N_B_c_222_p N_CIN_c_420_n 0.0144657f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_199 N_B_c_202_n N_CIN_c_420_n 0.00103514f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_200 N_B_M1030_g N_CIN_M1027_g 0.0293113f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_201 N_B_c_197_n N_CIN_c_422_n 0.044476f $X=4.06 $Y=1.66 $X2=0 $Y2=0
cc_202 N_B_c_226_p N_CIN_c_422_n 0.0173647f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_203 N_B_c_211_n N_CIN_c_422_n 0.00388862f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B_c_198_n N_CIN_c_423_n 0.071327f $X=6.1 $Y=1.66 $X2=0 $Y2=0
cc_205 B N_CIN_c_423_n 0.0163416f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_206 B N_CIN_c_423_n 0.006389f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_207 N_B_M1037_g N_CIN_c_424_n 0.0538055f $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_208 N_B_c_197_n N_CIN_c_425_n 0.00108757f $X=4.06 $Y=1.66 $X2=0 $Y2=0
cc_209 N_B_c_211_n N_CIN_c_425_n 0.0194879f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_210 N_B_M1023_g N_CIN_c_426_n 0.00166151f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_211 N_B_c_195_n N_CIN_c_426_n 0.00263938f $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_212 N_B_c_222_p N_CIN_c_426_n 0.00534188f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_213 N_B_c_202_n N_CIN_c_426_n 0.025012f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_214 N_B_c_226_p N_CIN_c_426_n 0.00606814f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_215 N_B_M1023_g N_CIN_c_427_n 7.01969e-19 $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_216 N_B_c_195_n N_CIN_c_427_n 6.81723e-19 $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_217 N_B_c_200_n N_CIN_c_427_n 0.00117817f $X=1.665 $Y=1.417 $X2=0 $Y2=0
cc_218 N_B_c_222_p N_CIN_c_427_n 0.0019211f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_219 N_B_c_202_n N_CIN_c_427_n 0.0013005f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_220 N_B_M1030_g N_CIN_c_428_n 0.00157687f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_221 N_B_c_197_n N_CIN_c_428_n 0.00277849f $X=4.06 $Y=1.66 $X2=0 $Y2=0
cc_222 N_B_c_226_p N_CIN_c_428_n 0.00741335f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_223 N_B_c_211_n N_CIN_c_428_n 0.0245256f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_224 N_B_c_212_n N_CIN_c_428_n 0.00817269f $X=4.62 $Y=1.805 $X2=0 $Y2=0
cc_225 B N_CIN_c_428_n 0.0132988f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_226 N_B_M1023_g N_CIN_c_429_n 6.4019e-19 $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_227 N_B_c_195_n N_CIN_c_429_n 6.86607e-19 $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_228 N_B_c_202_n N_CIN_c_429_n 0.00130776f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_229 N_B_c_226_p N_CIN_c_429_n 0.00249006f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_230 B N_CIN_c_430_n 0.0035103f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_231 B N_CIN_c_430_n 9.68406e-19 $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_232 N_B_c_198_n N_CIN_c_431_n 3.67751e-19 $X=6.1 $Y=1.66 $X2=0 $Y2=0
cc_233 N_B_M1037_g N_CIN_c_431_n 3.61499e-19 $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_234 B N_CIN_c_431_n 0.022365f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_235 B N_CIN_c_431_n 0.0224776f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_236 N_B_M1026_g N_CIN_c_432_n 3.51335e-19 $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_237 N_B_M1023_g N_CIN_c_432_n 0.00105583f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_238 N_B_c_195_n N_CIN_c_432_n 0.00218974f $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_239 N_B_c_200_n N_CIN_c_432_n 0.0243757f $X=1.665 $Y=1.417 $X2=0 $Y2=0
cc_240 N_B_c_201_n N_CIN_c_432_n 4.09781e-19 $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_241 N_B_c_209_n N_CIN_c_432_n 0.0158327f $X=1.75 $Y=1.95 $X2=0 $Y2=0
cc_242 N_B_c_222_p N_CIN_c_432_n 0.0119597f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_243 N_B_c_202_n N_CIN_c_432_n 0.0317861f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_244 N_B_M1023_g N_CIN_c_433_n 8.34658e-19 $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_245 N_B_c_195_n N_CIN_c_433_n 0.00176431f $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_246 N_B_c_202_n N_CIN_c_433_n 0.0223381f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_247 N_B_c_226_p N_CIN_c_433_n 0.0451733f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_248 N_B_c_222_p N_A_418_74#_M1029_d 0.00566684f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_249 B N_A_418_74#_c_571_n 0.0171659f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_250 N_B_c_204_n N_A_418_74#_c_576_n 0.00304206f $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_251 N_B_M1026_g N_A_418_74#_c_576_n 0.00442274f $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_252 N_B_c_200_n N_A_418_74#_c_576_n 0.0232015f $X=1.665 $Y=1.417 $X2=0 $Y2=0
cc_253 N_B_c_201_n N_A_418_74#_c_576_n 0.015156f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_254 N_B_c_209_n N_A_418_74#_c_576_n 0.00545885f $X=1.75 $Y=1.95 $X2=0 $Y2=0
cc_255 N_B_c_204_n N_A_418_74#_c_599_n 0.0105918f $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_256 N_B_c_209_n N_A_418_74#_c_599_n 0.00250585f $X=1.75 $Y=1.95 $X2=0 $Y2=0
cc_257 N_B_c_281_p N_A_418_74#_c_599_n 0.0138309f $X=1.835 $Y=2.035 $X2=0 $Y2=0
cc_258 N_B_c_222_p N_A_418_74#_c_602_n 0.0224059f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_259 N_B_c_281_p N_A_418_74#_c_602_n 0.0137412f $X=1.835 $Y=2.035 $X2=0 $Y2=0
cc_260 N_B_c_204_n N_A_418_74#_c_604_n 0.00372332f $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_261 N_B_M1023_g N_A_418_74#_c_577_n 0.00341585f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_262 N_B_M1030_g N_A_418_74#_c_606_n 0.0110518f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_263 N_B_c_197_n N_A_418_74#_c_606_n 0.00309208f $X=4.06 $Y=1.66 $X2=0 $Y2=0
cc_264 N_B_c_226_p N_A_418_74#_c_606_n 0.00177476f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_265 N_B_c_211_n N_A_418_74#_c_606_n 0.0184553f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_266 N_B_c_212_n N_A_418_74#_c_606_n 0.00330149f $X=4.62 $Y=1.805 $X2=0 $Y2=0
cc_267 B N_A_418_74#_c_606_n 0.00301153f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_268 N_B_M1037_g N_A_418_74#_c_578_n 0.0102703f $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_269 N_B_M1037_g N_A_418_74#_c_613_n 0.00376916f $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_270 N_B_M1037_g N_A_418_74#_c_614_n 0.00295923f $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_271 N_B_c_204_n N_A_418_74#_c_615_n 0.0132744f $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_272 N_B_c_200_n N_A_418_74#_c_615_n 0.0110357f $X=1.665 $Y=1.417 $X2=0 $Y2=0
cc_273 N_B_c_201_n N_A_418_74#_c_615_n 0.00579157f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B_c_209_n N_A_418_74#_c_615_n 0.0133105f $X=1.75 $Y=1.95 $X2=0 $Y2=0
cc_275 N_B_M1026_g N_A_418_74#_c_619_n 0.0124111f $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_276 N_B_c_200_n N_A_418_74#_c_619_n 0.0208902f $X=1.665 $Y=1.417 $X2=0 $Y2=0
cc_277 N_B_c_201_n N_A_418_74#_c_619_n 0.00858317f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_278 N_B_c_200_n N_A_418_74#_c_622_n 0.0124459f $X=1.665 $Y=1.417 $X2=0 $Y2=0
cc_279 N_B_c_195_n N_A_418_74#_c_590_n 0.0104027f $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_280 N_B_c_222_p N_A_418_74#_c_590_n 0.0156687f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_281 N_B_c_305_p N_A_418_74#_c_590_n 0.00111187f $X=2.645 $Y=1.83 $X2=0 $Y2=0
cc_282 N_B_M1023_g N_A_418_74#_c_626_n 0.0133548f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_283 N_B_c_195_n N_A_418_74#_c_626_n 8.31921e-19 $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_284 N_B_c_202_n N_A_418_74#_c_626_n 0.0122929f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_285 N_B_M1030_g N_A_418_74#_c_629_n 3.88992e-19 $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_286 N_B_c_211_n N_A_418_74#_c_582_n 0.00547767f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_287 B N_A_418_74#_c_582_n 0.0243477f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_288 N_B_c_204_n N_A_c_863_n 0.00448518f $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_289 N_B_c_201_n N_A_c_863_n 0.00181091f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_290 N_B_c_204_n N_A_M1028_g 0.0159616f $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_291 N_B_c_204_n N_A_c_878_n 0.00885198f $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_292 N_B_c_195_n N_A_c_878_n 0.0103487f $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_293 N_B_M1023_g N_A_c_865_n 0.00188318f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_294 N_B_c_195_n N_A_c_865_n 0.0212026f $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_295 N_B_c_202_n N_A_c_865_n 4.82448e-19 $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_296 N_B_c_195_n N_A_c_881_n 0.00206952f $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_297 N_B_c_195_n N_A_c_883_n 0.00281869f $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_298 N_B_c_202_n N_A_c_883_n 0.00196148f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_299 N_B_c_195_n N_A_M1001_g 0.0367853f $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_300 N_B_c_202_n N_A_M1001_g 0.00191446f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_301 N_B_c_226_p N_A_M1001_g 0.0153252f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_302 N_B_c_305_p N_A_M1001_g 0.00107976f $X=2.645 $Y=1.83 $X2=0 $Y2=0
cc_303 N_B_c_197_n N_A_c_885_n 0.0103487f $X=4.06 $Y=1.66 $X2=0 $Y2=0
cc_304 N_B_c_197_n N_A_c_867_n 0.0169287f $X=4.06 $Y=1.66 $X2=0 $Y2=0
cc_305 N_B_c_211_n N_A_c_867_n 0.00145815f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_306 N_B_c_197_n N_A_c_887_n 0.00129916f $X=4.06 $Y=1.66 $X2=0 $Y2=0
cc_307 N_B_c_197_n N_A_c_889_n 0.00224408f $X=4.06 $Y=1.66 $X2=0 $Y2=0
cc_308 N_B_c_211_n N_A_c_889_n 0.00189295f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_309 N_B_c_212_n N_A_c_889_n 5.3878e-19 $X=4.62 $Y=1.805 $X2=0 $Y2=0
cc_310 B N_A_c_889_n 4.9691e-19 $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_311 N_B_c_197_n N_A_M1004_g 0.0253033f $X=4.06 $Y=1.66 $X2=0 $Y2=0
cc_312 N_B_c_211_n N_A_M1004_g 0.00138719f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_313 N_B_c_212_n N_A_M1004_g 0.00716159f $X=4.62 $Y=1.805 $X2=0 $Y2=0
cc_314 B N_A_M1004_g 0.00707418f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_315 N_B_c_198_n N_A_c_891_n 0.0104164f $X=6.1 $Y=1.66 $X2=0 $Y2=0
cc_316 N_B_c_198_n N_A_M1039_g 0.0226014f $X=6.1 $Y=1.66 $X2=0 $Y2=0
cc_317 N_B_M1037_g N_A_M1039_g 0.0321719f $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_318 B N_A_M1039_g 0.00394145f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_319 N_B_c_198_n N_A_c_870_n 0.00318167f $X=6.1 $Y=1.66 $X2=0 $Y2=0
cc_320 B N_A_c_870_n 0.00474782f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_321 N_B_c_198_n N_A_M1012_g 0.034867f $X=6.1 $Y=1.66 $X2=0 $Y2=0
cc_322 B N_A_M1012_g 0.00135925f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_323 N_B_M1023_g N_A_c_871_n 0.0295343f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_324 N_B_M1030_g N_A_c_872_n 0.0260938f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_325 N_B_c_204_n A 4.48262e-19 $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_326 N_B_c_201_n A 0.00146034f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_327 N_B_c_201_n N_A_c_874_n 0.0157952f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_328 B N_A_1024_74#_M1006_d 0.00250873f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_329 N_B_c_198_n N_A_1024_74#_c_1081_n 0.0148981f $X=6.1 $Y=1.66 $X2=0 $Y2=0
cc_330 B N_A_1024_74#_c_1081_n 0.020193f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_331 B N_A_1024_74#_c_1081_n 0.0145837f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_332 N_B_c_198_n N_A_1024_74#_c_1084_n 0.00329274f $X=6.1 $Y=1.66 $X2=0 $Y2=0
cc_333 N_B_M1037_g N_A_1024_74#_c_1084_n 0.00801378f $X=6.115 $Y=0.74 $X2=0
+ $Y2=0
cc_334 B N_A_1024_74#_c_1084_n 0.00823733f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_335 B N_A_1024_74#_c_1087_n 0.0106484f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_336 B N_A_1024_74#_c_1068_n 0.00244385f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_337 B N_A_1024_74#_c_1076_n 0.00554062f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_338 N_B_c_198_n N_A_1024_74#_c_1078_n 0.00246868f $X=6.1 $Y=1.66 $X2=0 $Y2=0
cc_339 B N_A_1024_74#_c_1078_n 0.0203373f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_340 N_B_M1037_g N_A_1024_74#_c_1092_n 9.8919e-19 $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_341 N_B_M1037_g N_A_1024_74#_c_1093_n 0.00623463f $X=6.115 $Y=0.74 $X2=0
+ $Y2=0
cc_342 B N_A_1024_74#_c_1093_n 0.0290034f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_343 N_B_c_198_n N_A_1024_74#_c_1095_n 0.00345516f $X=6.1 $Y=1.66 $X2=0 $Y2=0
cc_344 B N_A_1024_74#_c_1095_n 0.0135032f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_345 B N_A_1024_74#_c_1070_n 0.0140535f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_346 N_B_c_209_n N_A_27_392#_M1010_d 0.00660674f $X=1.75 $Y=1.95 $X2=0 $Y2=0
cc_347 N_B_c_222_p N_A_27_392#_M1010_d 0.00745696f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_348 N_B_c_281_p N_A_27_392#_M1010_d 0.00510287f $X=1.835 $Y=2.035 $X2=0 $Y2=0
cc_349 N_B_c_204_n N_A_27_392#_c_1223_n 5.81223e-19 $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_350 N_B_c_204_n N_A_27_392#_c_1224_n 2.38328e-19 $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_351 N_B_c_204_n N_A_27_392#_c_1232_n 0.00647737f $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_352 N_B_c_204_n N_A_27_392#_c_1233_n 0.0141409f $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_353 N_B_c_204_n N_A_27_392#_c_1225_n 0.00435061f $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_354 N_B_c_204_n N_A_27_392#_c_1226_n 0.0111103f $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_355 N_B_c_226_p N_VPWR_M1001_d 0.00476945f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_356 N_B_c_212_n N_VPWR_M1003_d 0.00699981f $X=4.62 $Y=1.805 $X2=0 $Y2=0
cc_357 N_B_c_204_n N_VPWR_c_1275_n 0.00130424f $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_358 N_B_c_195_n N_VPWR_c_1276_n 0.00280645f $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_359 N_B_c_226_p N_VPWR_c_1276_n 0.0202249f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_360 N_B_c_305_p N_VPWR_c_1276_n 0.00111629f $X=2.645 $Y=1.83 $X2=0 $Y2=0
cc_361 N_B_c_197_n N_VPWR_c_1277_n 0.00401111f $X=4.06 $Y=1.66 $X2=0 $Y2=0
cc_362 N_B_c_195_n N_VPWR_c_1274_n 9.39239e-19 $X=2.6 $Y=1.66 $X2=0 $Y2=0
cc_363 N_B_c_197_n N_VPWR_c_1274_n 9.39239e-19 $X=4.06 $Y=1.66 $X2=0 $Y2=0
cc_364 N_B_c_198_n N_VPWR_c_1274_n 9.39239e-19 $X=6.1 $Y=1.66 $X2=0 $Y2=0
cc_365 N_B_c_226_p A_535_347# 0.00904452f $X=3.95 $Y=1.83 $X2=-0.19 $Y2=-0.245
cc_366 N_B_c_305_p A_535_347# 0.00346735f $X=2.645 $Y=1.83 $X2=-0.19 $Y2=-0.245
cc_367 N_B_c_226_p N_A_737_347#_M1005_d 0.00546464f $X=3.95 $Y=1.83 $X2=-0.19
+ $Y2=-0.245
cc_368 B N_A_737_347#_M1004_d 0.00266f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_369 N_B_c_197_n N_A_737_347#_c_1431_n 0.0126926f $X=4.06 $Y=1.66 $X2=0 $Y2=0
cc_370 N_B_c_212_n N_A_737_347#_c_1431_n 0.0377865f $X=4.62 $Y=1.805 $X2=0 $Y2=0
cc_371 B N_A_737_347#_c_1431_n 0.00513153f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_372 B N_A_737_347#_c_1434_n 0.0182961f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_373 N_B_c_197_n N_A_737_347#_c_1428_n 0.00769916f $X=4.06 $Y=1.66 $X2=0 $Y2=0
cc_374 N_B_c_226_p N_A_737_347#_c_1428_n 0.0162136f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_375 N_B_c_212_n N_A_737_347#_c_1428_n 0.00122259f $X=4.62 $Y=1.805 $X2=0
+ $Y2=0
cc_376 B A_1141_347# 0.00161973f $X=5.915 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_377 B A_1141_347# 5.86586e-19 $X=6.395 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_378 B A_1235_347# 0.00230047f $X=6.395 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_379 N_B_M1026_g N_A_27_74#_c_1595_n 0.0150217f $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_380 N_B_c_201_n N_A_27_74#_c_1599_n 7.61744e-19 $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_381 N_B_M1023_g N_VGND_c_1627_n 0.00200275f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_382 N_B_M1026_g N_VGND_c_1631_n 0.00291649f $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_383 N_B_M1023_g N_VGND_c_1631_n 0.00461464f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_384 N_B_M1030_g N_VGND_c_1633_n 0.00220663f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_385 N_B_M1030_g N_VGND_c_1634_n 0.00316493f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_386 N_B_M1037_g N_VGND_c_1635_n 0.00278271f $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_387 N_B_M1026_g N_VGND_c_1641_n 0.00383588f $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_388 N_B_M1026_g N_VGND_c_1646_n 0.00364217f $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_389 N_B_M1023_g N_VGND_c_1646_n 0.0046687f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_390 N_B_M1030_g N_VGND_c_1646_n 0.00393316f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_391 N_B_M1037_g N_VGND_c_1646_n 0.00353931f $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_392 N_B_M1030_g N_A_734_74#_c_1776_n 0.00936301f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_393 N_B_M1030_g N_A_734_74#_c_1774_n 0.00573013f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_394 N_B_M1030_g N_A_734_74#_c_1775_n 8.6409e-19 $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_395 N_CIN_c_424_n N_A_418_74#_c_570_n 0.0134862f $X=5.725 $Y=1.22 $X2=0 $Y2=0
cc_396 N_CIN_c_423_n N_A_418_74#_c_571_n 0.0536236f $X=5.63 $Y=1.66 $X2=0 $Y2=0
cc_397 N_CIN_c_428_n N_A_418_74#_c_571_n 0.0013891f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_398 N_CIN_c_431_n N_A_418_74#_c_571_n 9.45146e-19 $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_399 N_CIN_c_420_n N_A_418_74#_c_599_n 0.0043641f $X=2.15 $Y=1.66 $X2=0 $Y2=0
cc_400 N_CIN_c_420_n N_A_418_74#_c_602_n 0.0111182f $X=2.15 $Y=1.66 $X2=0 $Y2=0
cc_401 N_CIN_c_419_n N_A_418_74#_c_638_n 0.0139672f $X=2.015 $Y=1.22 $X2=0 $Y2=0
cc_402 N_CIN_c_427_n N_A_418_74#_c_638_n 8.8084e-19 $X=2.305 $Y=1.295 $X2=0
+ $Y2=0
cc_403 N_CIN_c_432_n N_A_418_74#_c_638_n 0.00689032f $X=2.16 $Y=1.295 $X2=0
+ $Y2=0
cc_404 N_CIN_c_419_n N_A_418_74#_c_577_n 0.00305832f $X=2.015 $Y=1.22 $X2=0
+ $Y2=0
cc_405 N_CIN_M1027_g N_A_418_74#_c_606_n 0.0102982f $X=3.595 $Y=0.74 $X2=0 $Y2=0
cc_406 N_CIN_c_422_n N_A_418_74#_c_606_n 0.00112445f $X=3.61 $Y=1.66 $X2=0 $Y2=0
cc_407 N_CIN_c_424_n N_A_418_74#_c_644_n 0.00343696f $X=5.725 $Y=1.22 $X2=0
+ $Y2=0
cc_408 N_CIN_c_424_n N_A_418_74#_c_578_n 0.0109994f $X=5.725 $Y=1.22 $X2=0 $Y2=0
cc_409 N_CIN_c_419_n N_A_418_74#_c_622_n 0.00235187f $X=2.015 $Y=1.22 $X2=0
+ $Y2=0
cc_410 N_CIN_c_420_n N_A_418_74#_c_647_n 9.10263e-19 $X=2.15 $Y=1.66 $X2=0 $Y2=0
cc_411 N_CIN_c_426_n N_A_418_74#_c_647_n 0.00798157f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_412 N_CIN_c_427_n N_A_418_74#_c_647_n 0.00288269f $X=2.305 $Y=1.295 $X2=0
+ $Y2=0
cc_413 N_CIN_c_432_n N_A_418_74#_c_647_n 0.0098023f $X=2.16 $Y=1.295 $X2=0 $Y2=0
cc_414 N_CIN_c_420_n N_A_418_74#_c_590_n 0.0110727f $X=2.15 $Y=1.66 $X2=0 $Y2=0
cc_415 N_CIN_c_425_n N_A_418_74#_c_626_n 0.00659689f $X=3.575 $Y=1.41 $X2=0
+ $Y2=0
cc_416 N_CIN_c_426_n N_A_418_74#_c_626_n 0.0153931f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_417 N_CIN_c_428_n N_A_418_74#_c_626_n 0.00299186f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_418 N_CIN_c_429_n N_A_418_74#_c_626_n 0.00799415f $X=3.265 $Y=1.295 $X2=0
+ $Y2=0
cc_419 N_CIN_c_433_n N_A_418_74#_c_626_n 0.0111957f $X=3.215 $Y=1.377 $X2=0
+ $Y2=0
cc_420 N_CIN_M1027_g N_A_418_74#_c_629_n 0.00631936f $X=3.595 $Y=0.74 $X2=0
+ $Y2=0
cc_421 N_CIN_c_422_n N_A_418_74#_c_629_n 0.0018054f $X=3.61 $Y=1.66 $X2=0 $Y2=0
cc_422 N_CIN_c_425_n N_A_418_74#_c_629_n 0.0185241f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_423 N_CIN_c_428_n N_A_418_74#_c_629_n 0.0441427f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_424 N_CIN_c_423_n N_A_418_74#_c_582_n 4.59775e-19 $X=5.63 $Y=1.66 $X2=0 $Y2=0
cc_425 N_CIN_c_424_n N_A_418_74#_c_582_n 0.00293705f $X=5.725 $Y=1.22 $X2=0
+ $Y2=0
cc_426 N_CIN_c_428_n N_A_418_74#_c_582_n 0.0310488f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_427 N_CIN_c_430_n N_A_418_74#_c_582_n 0.0027738f $X=5.52 $Y=1.295 $X2=0 $Y2=0
cc_428 N_CIN_c_431_n N_A_418_74#_c_582_n 0.0267617f $X=5.52 $Y=1.295 $X2=0 $Y2=0
cc_429 N_CIN_c_420_n N_A_c_878_n 0.0100467f $X=2.15 $Y=1.66 $X2=0 $Y2=0
cc_430 N_CIN_c_422_n N_A_c_865_n 0.0213361f $X=3.61 $Y=1.66 $X2=0 $Y2=0
cc_431 N_CIN_c_433_n N_A_c_865_n 0.00270838f $X=3.215 $Y=1.377 $X2=0 $Y2=0
cc_432 N_CIN_c_433_n N_A_c_866_n 0.0080712f $X=3.215 $Y=1.377 $X2=0 $Y2=0
cc_433 N_CIN_c_422_n N_A_c_881_n 0.00171838f $X=3.61 $Y=1.66 $X2=0 $Y2=0
cc_434 N_CIN_c_422_n N_A_c_883_n 0.0039344f $X=3.61 $Y=1.66 $X2=0 $Y2=0
cc_435 N_CIN_c_433_n N_A_c_883_n 0.00242018f $X=3.215 $Y=1.377 $X2=0 $Y2=0
cc_436 N_CIN_c_422_n N_A_M1001_g 0.0248211f $X=3.61 $Y=1.66 $X2=0 $Y2=0
cc_437 N_CIN_c_422_n N_A_c_885_n 0.0103487f $X=3.61 $Y=1.66 $X2=0 $Y2=0
cc_438 N_CIN_c_428_n N_A_c_867_n 0.00251789f $X=5.375 $Y=1.295 $X2=0 $Y2=0
cc_439 N_CIN_c_428_n N_A_c_868_n 0.0036588f $X=5.375 $Y=1.295 $X2=0 $Y2=0
cc_440 N_CIN_c_423_n N_A_c_891_n 0.0103487f $X=5.63 $Y=1.66 $X2=0 $Y2=0
cc_441 N_CIN_M1027_g N_A_c_871_n 0.0241987f $X=3.595 $Y=0.74 $X2=0 $Y2=0
cc_442 N_CIN_c_429_n N_A_c_871_n 0.00140441f $X=3.265 $Y=1.295 $X2=0 $Y2=0
cc_443 N_CIN_c_433_n N_A_c_871_n 0.00117185f $X=3.215 $Y=1.377 $X2=0 $Y2=0
cc_444 N_CIN_c_423_n N_A_1024_74#_c_1081_n 0.0118586f $X=5.63 $Y=1.66 $X2=0
+ $Y2=0
cc_445 N_CIN_c_423_n N_A_1024_74#_c_1078_n 0.0109951f $X=5.63 $Y=1.66 $X2=0
+ $Y2=0
cc_446 N_CIN_c_423_n N_A_1024_74#_c_1092_n 0.00107113f $X=5.63 $Y=1.66 $X2=0
+ $Y2=0
cc_447 N_CIN_c_424_n N_A_1024_74#_c_1092_n 0.00623624f $X=5.725 $Y=1.22 $X2=0
+ $Y2=0
cc_448 N_CIN_c_430_n N_A_1024_74#_c_1092_n 0.00673868f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_449 N_CIN_c_431_n N_A_1024_74#_c_1092_n 0.0151874f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_450 N_CIN_c_424_n N_A_1024_74#_c_1104_n 0.0102416f $X=5.725 $Y=1.22 $X2=0
+ $Y2=0
cc_451 N_CIN_c_431_n N_A_1024_74#_c_1104_n 0.00504528f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_452 N_CIN_c_424_n N_A_1024_74#_c_1093_n 0.00111404f $X=5.725 $Y=1.22 $X2=0
+ $Y2=0
cc_453 N_CIN_c_432_n N_A_27_392#_M1010_d 6.19023e-19 $X=2.16 $Y=1.295 $X2=0
+ $Y2=0
cc_454 N_CIN_c_420_n N_A_27_392#_c_1226_n 0.00793173f $X=2.15 $Y=1.66 $X2=0
+ $Y2=0
cc_455 N_CIN_c_422_n N_VPWR_c_1276_n 0.00537823f $X=3.61 $Y=1.66 $X2=0 $Y2=0
cc_456 N_CIN_c_420_n N_VPWR_c_1274_n 9.39239e-19 $X=2.15 $Y=1.66 $X2=0 $Y2=0
cc_457 N_CIN_c_422_n N_VPWR_c_1274_n 9.39239e-19 $X=3.61 $Y=1.66 $X2=0 $Y2=0
cc_458 N_CIN_c_423_n N_VPWR_c_1274_n 9.39239e-19 $X=5.63 $Y=1.66 $X2=0 $Y2=0
cc_459 N_CIN_c_422_n N_A_737_347#_c_1428_n 0.0073664f $X=3.61 $Y=1.66 $X2=0
+ $Y2=0
cc_460 N_CIN_c_419_n N_A_27_74#_c_1595_n 0.00409096f $X=2.015 $Y=1.22 $X2=0
+ $Y2=0
cc_461 N_CIN_M1027_g N_VGND_c_1627_n 0.00193337f $X=3.595 $Y=0.74 $X2=0 $Y2=0
cc_462 N_CIN_c_419_n N_VGND_c_1631_n 0.00433162f $X=2.015 $Y=1.22 $X2=0 $Y2=0
cc_463 N_CIN_M1027_g N_VGND_c_1634_n 0.00461464f $X=3.595 $Y=0.74 $X2=0 $Y2=0
cc_464 N_CIN_c_424_n N_VGND_c_1635_n 0.00278271f $X=5.725 $Y=1.22 $X2=0 $Y2=0
cc_465 N_CIN_c_419_n N_VGND_c_1646_n 0.0044836f $X=2.015 $Y=1.22 $X2=0 $Y2=0
cc_466 N_CIN_M1027_g N_VGND_c_1646_n 0.00804222f $X=3.595 $Y=0.74 $X2=0 $Y2=0
cc_467 N_CIN_c_424_n N_VGND_c_1646_n 0.00354203f $X=5.725 $Y=1.22 $X2=0 $Y2=0
cc_468 N_A_418_74#_c_576_n N_A_c_863_n 3.57059e-19 $X=1.09 $Y=1.745 $X2=0 $Y2=0
cc_469 N_A_418_74#_c_615_n N_A_c_863_n 0.00228655f $X=1.41 $Y=1.83 $X2=0 $Y2=0
cc_470 N_A_418_74#_c_576_n N_A_M1032_g 0.00398634f $X=1.09 $Y=1.745 $X2=0 $Y2=0
cc_471 N_A_418_74#_c_669_p N_A_M1032_g 0.00328708f $X=1.175 $Y=1.005 $X2=0 $Y2=0
cc_472 N_A_418_74#_c_615_n N_A_M1028_g 5.8864e-19 $X=1.41 $Y=1.83 $X2=0 $Y2=0
cc_473 N_A_418_74#_c_602_n N_A_c_878_n 0.00180339f $X=2.21 $Y=2.375 $X2=0 $Y2=0
cc_474 N_A_418_74#_c_590_n N_A_c_878_n 0.00600601f $X=2.375 $Y=2.375 $X2=0 $Y2=0
cc_475 N_A_418_74#_c_590_n N_A_M1001_g 0.00141636f $X=2.375 $Y=2.375 $X2=0 $Y2=0
cc_476 N_A_418_74#_c_570_n N_A_c_867_n 0.00165443f $X=5.045 $Y=1.22 $X2=0 $Y2=0
cc_477 N_A_418_74#_c_571_n N_A_c_867_n 0.0208244f $X=5.13 $Y=1.66 $X2=0 $Y2=0
cc_478 N_A_418_74#_c_582_n N_A_c_867_n 0.00253264f $X=5.095 $Y=1.005 $X2=0 $Y2=0
cc_479 N_A_418_74#_c_571_n N_A_c_868_n 0.00506843f $X=5.13 $Y=1.66 $X2=0 $Y2=0
cc_480 N_A_418_74#_c_571_n N_A_c_887_n 0.00213258f $X=5.13 $Y=1.66 $X2=0 $Y2=0
cc_481 N_A_418_74#_c_571_n N_A_M1004_g 0.0256634f $X=5.13 $Y=1.66 $X2=0 $Y2=0
cc_482 N_A_418_74#_c_571_n N_A_c_891_n 0.0103487f $X=5.13 $Y=1.66 $X2=0 $Y2=0
cc_483 N_A_418_74#_c_578_n N_A_M1039_g 0.00209511f $X=6.255 $Y=0.34 $X2=0 $Y2=0
cc_484 N_A_418_74#_c_613_n N_A_M1039_g 0.00349056f $X=6.34 $Y=0.58 $X2=0 $Y2=0
cc_485 N_A_418_74#_c_683_p N_A_M1039_g 0.012131f $X=8.965 $Y=0.665 $X2=0 $Y2=0
cc_486 N_A_418_74#_c_626_n N_A_c_871_n 0.0122961f $X=3.385 $Y=0.965 $X2=0 $Y2=0
cc_487 N_A_418_74#_c_629_n N_A_c_871_n 0.00216961f $X=3.555 $Y=0.965 $X2=0 $Y2=0
cc_488 N_A_418_74#_c_570_n N_A_c_872_n 0.0249033f $X=5.045 $Y=1.22 $X2=0 $Y2=0
cc_489 N_A_418_74#_c_606_n N_A_c_872_n 0.0127471f $X=4.93 $Y=1.005 $X2=0 $Y2=0
cc_490 N_A_418_74#_c_644_n N_A_c_872_n 9.47922e-19 $X=5.17 $Y=0.92 $X2=0 $Y2=0
cc_491 N_A_418_74#_c_579_n N_A_c_872_n 3.23044e-19 $X=5.255 $Y=0.34 $X2=0 $Y2=0
cc_492 N_A_418_74#_c_582_n N_A_c_872_n 0.00165995f $X=5.095 $Y=1.005 $X2=0 $Y2=0
cc_493 N_A_418_74#_c_576_n A 0.0422556f $X=1.09 $Y=1.745 $X2=0 $Y2=0
cc_494 N_A_418_74#_c_615_n A 0.00291429f $X=1.41 $Y=1.83 $X2=0 $Y2=0
cc_495 N_A_418_74#_c_576_n N_A_c_874_n 9.1952e-19 $X=1.09 $Y=1.745 $X2=0 $Y2=0
cc_496 N_A_418_74#_c_644_n N_A_1024_74#_M1016_d 0.00532706f $X=5.17 $Y=0.92
+ $X2=-0.19 $Y2=-0.245
cc_497 N_A_418_74#_c_578_n N_A_1024_74#_M1016_d 0.0087698f $X=6.255 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_498 N_A_418_74#_c_582_n N_A_1024_74#_M1016_d 0.00250765f $X=5.095 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_499 N_A_418_74#_c_683_p N_A_1024_74#_M1020_g 0.0136954f $X=8.965 $Y=0.665
+ $X2=0 $Y2=0
cc_500 N_A_418_74#_c_683_p N_A_1024_74#_M1021_g 0.0120977f $X=8.965 $Y=0.665
+ $X2=0 $Y2=0
cc_501 N_A_418_74#_c_683_p N_A_1024_74#_M1034_g 0.0120967f $X=8.965 $Y=0.665
+ $X2=0 $Y2=0
cc_502 N_A_418_74#_c_585_n N_A_1024_74#_c_1075_n 0.0204913f $X=9.085 $Y=1.765
+ $X2=0 $Y2=0
cc_503 N_A_418_74#_M1013_g N_A_1024_74#_M1036_g 0.021129f $X=9.255 $Y=0.78 $X2=0
+ $Y2=0
cc_504 N_A_418_74#_c_683_p N_A_1024_74#_M1036_g 0.0156149f $X=8.965 $Y=0.665
+ $X2=0 $Y2=0
cc_505 N_A_418_74#_c_580_n N_A_1024_74#_M1036_g 0.00692925f $X=9.05 $Y=1.32
+ $X2=0 $Y2=0
cc_506 N_A_418_74#_c_581_n N_A_1024_74#_M1036_g 0.0017339f $X=9.135 $Y=1.485
+ $X2=0 $Y2=0
cc_507 N_A_418_74#_c_583_n N_A_1024_74#_M1036_g 0.00877228f $X=10.485 $Y=1.542
+ $X2=0 $Y2=0
cc_508 N_A_418_74#_c_578_n N_A_1024_74#_c_1084_n 0.00321187f $X=6.255 $Y=0.34
+ $X2=0 $Y2=0
cc_509 N_A_418_74#_c_683_p N_A_1024_74#_c_1084_n 0.0396142f $X=8.965 $Y=0.665
+ $X2=0 $Y2=0
cc_510 N_A_418_74#_c_614_n N_A_1024_74#_c_1084_n 0.0134799f $X=6.425 $Y=0.665
+ $X2=0 $Y2=0
cc_511 N_A_418_74#_c_683_p N_A_1024_74#_c_1069_n 0.00424675f $X=8.965 $Y=0.665
+ $X2=0 $Y2=0
cc_512 N_A_418_74#_c_571_n N_A_1024_74#_c_1078_n 0.00285784f $X=5.13 $Y=1.66
+ $X2=0 $Y2=0
cc_513 N_A_418_74#_c_570_n N_A_1024_74#_c_1092_n 0.0012068f $X=5.045 $Y=1.22
+ $X2=0 $Y2=0
cc_514 N_A_418_74#_c_644_n N_A_1024_74#_c_1092_n 0.0242712f $X=5.17 $Y=0.92
+ $X2=0 $Y2=0
cc_515 N_A_418_74#_c_578_n N_A_1024_74#_c_1092_n 0.0138888f $X=6.255 $Y=0.34
+ $X2=0 $Y2=0
cc_516 N_A_418_74#_c_614_n N_A_1024_74#_c_1092_n 0.0047823f $X=6.425 $Y=0.665
+ $X2=0 $Y2=0
cc_517 N_A_418_74#_c_582_n N_A_1024_74#_c_1092_n 0.00751744f $X=5.095 $Y=1.005
+ $X2=0 $Y2=0
cc_518 N_A_418_74#_c_578_n N_A_1024_74#_c_1104_n 0.00892235f $X=6.255 $Y=0.34
+ $X2=0 $Y2=0
cc_519 N_A_418_74#_c_582_n N_A_1024_74#_c_1093_n 0.00253405f $X=5.095 $Y=1.005
+ $X2=0 $Y2=0
cc_520 N_A_418_74#_c_683_p N_A_1024_74#_c_1071_n 2.97785e-19 $X=8.965 $Y=0.665
+ $X2=0 $Y2=0
cc_521 N_A_418_74#_c_581_n N_A_1024_74#_c_1071_n 0.00159647f $X=9.135 $Y=1.485
+ $X2=0 $Y2=0
cc_522 N_A_418_74#_c_583_n N_A_1024_74#_c_1071_n 0.0111329f $X=10.485 $Y=1.542
+ $X2=0 $Y2=0
cc_523 N_A_418_74#_c_599_n N_A_27_392#_M1010_d 0.0112914f $X=1.41 $Y=2.29 $X2=0
+ $Y2=0
cc_524 N_A_418_74#_c_602_n N_A_27_392#_M1010_d 0.0190762f $X=2.21 $Y=2.375 $X2=0
+ $Y2=0
cc_525 N_A_418_74#_c_604_n N_A_27_392#_M1010_d 0.004618f $X=1.495 $Y=2.375 $X2=0
+ $Y2=0
cc_526 N_A_418_74#_c_615_n N_A_27_392#_M1010_d 0.00647549f $X=1.41 $Y=1.83 $X2=0
+ $Y2=0
cc_527 N_A_418_74#_c_599_n N_A_27_392#_c_1232_n 0.0133617f $X=1.41 $Y=2.29 $X2=0
+ $Y2=0
cc_528 N_A_418_74#_c_615_n N_A_27_392#_c_1232_n 0.00714112f $X=1.41 $Y=1.83
+ $X2=0 $Y2=0
cc_529 N_A_418_74#_c_599_n N_A_27_392#_c_1233_n 0.00238695f $X=1.41 $Y=2.29
+ $X2=0 $Y2=0
cc_530 N_A_418_74#_c_604_n N_A_27_392#_c_1233_n 0.0134181f $X=1.495 $Y=2.375
+ $X2=0 $Y2=0
cc_531 N_A_418_74#_c_602_n N_A_27_392#_c_1226_n 0.0389388f $X=2.21 $Y=2.375
+ $X2=0 $Y2=0
cc_532 N_A_418_74#_c_604_n N_A_27_392#_c_1226_n 0.0142344f $X=1.495 $Y=2.375
+ $X2=0 $Y2=0
cc_533 N_A_418_74#_c_590_n N_A_27_392#_c_1226_n 0.00889758f $X=2.375 $Y=2.375
+ $X2=0 $Y2=0
cc_534 N_A_418_74#_c_615_n N_VPWR_M1028_d 0.0027275f $X=1.41 $Y=1.83 $X2=-0.19
+ $Y2=-0.245
cc_535 N_A_418_74#_c_590_n N_VPWR_c_1276_n 0.0117468f $X=2.375 $Y=2.375 $X2=0
+ $Y2=0
cc_536 N_A_418_74#_c_571_n N_VPWR_c_1277_n 5.8697e-19 $X=5.13 $Y=1.66 $X2=0
+ $Y2=0
cc_537 N_A_418_74#_c_585_n N_VPWR_c_1280_n 0.00927148f $X=9.085 $Y=1.765 $X2=0
+ $Y2=0
cc_538 N_A_418_74#_c_581_n N_VPWR_c_1280_n 8.43278e-19 $X=9.135 $Y=1.485 $X2=0
+ $Y2=0
cc_539 N_A_418_74#_c_586_n N_VPWR_c_1281_n 0.00629151f $X=9.535 $Y=1.765 $X2=0
+ $Y2=0
cc_540 N_A_418_74#_c_587_n N_VPWR_c_1281_n 0.00740236f $X=10.035 $Y=1.765 $X2=0
+ $Y2=0
cc_541 N_A_418_74#_c_588_n N_VPWR_c_1283_n 0.00990712f $X=10.485 $Y=1.765 $X2=0
+ $Y2=0
cc_542 N_A_418_74#_c_590_n N_VPWR_c_1284_n 0.00727901f $X=2.375 $Y=2.375 $X2=0
+ $Y2=0
cc_543 N_A_418_74#_c_585_n N_VPWR_c_1290_n 0.00445602f $X=9.085 $Y=1.765 $X2=0
+ $Y2=0
cc_544 N_A_418_74#_c_586_n N_VPWR_c_1290_n 0.00445602f $X=9.535 $Y=1.765 $X2=0
+ $Y2=0
cc_545 N_A_418_74#_c_587_n N_VPWR_c_1291_n 0.00445602f $X=10.035 $Y=1.765 $X2=0
+ $Y2=0
cc_546 N_A_418_74#_c_588_n N_VPWR_c_1291_n 0.00434272f $X=10.485 $Y=1.765 $X2=0
+ $Y2=0
cc_547 N_A_418_74#_c_571_n N_VPWR_c_1274_n 9.39239e-19 $X=5.13 $Y=1.66 $X2=0
+ $Y2=0
cc_548 N_A_418_74#_c_585_n N_VPWR_c_1274_n 0.00857432f $X=9.085 $Y=1.765 $X2=0
+ $Y2=0
cc_549 N_A_418_74#_c_586_n N_VPWR_c_1274_n 0.0085805f $X=9.535 $Y=1.765 $X2=0
+ $Y2=0
cc_550 N_A_418_74#_c_587_n N_VPWR_c_1274_n 0.00857378f $X=10.035 $Y=1.765 $X2=0
+ $Y2=0
cc_551 N_A_418_74#_c_588_n N_VPWR_c_1274_n 0.00824551f $X=10.485 $Y=1.765 $X2=0
+ $Y2=0
cc_552 N_A_418_74#_c_590_n N_VPWR_c_1274_n 0.00889658f $X=2.375 $Y=2.375 $X2=0
+ $Y2=0
cc_553 N_A_418_74#_c_571_n N_A_737_347#_c_1434_n 0.001827f $X=5.13 $Y=1.66 $X2=0
+ $Y2=0
cc_554 N_A_418_74#_c_571_n N_A_737_347#_c_1427_n 0.00554049f $X=5.13 $Y=1.66
+ $X2=0 $Y2=0
cc_555 N_A_418_74#_c_683_p N_SUM_M1020_s 0.00437807f $X=8.965 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_556 N_A_418_74#_c_683_p N_SUM_M1034_s 0.00437412f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_557 N_A_418_74#_c_683_p N_SUM_c_1463_n 0.0576451f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_558 N_A_418_74#_c_683_p N_SUM_c_1464_n 0.0170377f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_559 N_A_418_74#_c_580_n N_SUM_c_1464_n 0.011264f $X=9.05 $Y=1.32 $X2=0 $Y2=0
cc_560 N_A_418_74#_c_585_n N_SUM_c_1465_n 2.56932e-19 $X=9.085 $Y=1.765 $X2=0
+ $Y2=0
cc_561 N_A_418_74#_c_580_n N_SUM_c_1465_n 0.00593841f $X=9.05 $Y=1.32 $X2=0
+ $Y2=0
cc_562 N_A_418_74#_c_581_n N_SUM_c_1465_n 0.0134827f $X=9.135 $Y=1.485 $X2=0
+ $Y2=0
cc_563 N_A_418_74#_c_583_n N_SUM_c_1465_n 8.34232e-19 $X=10.485 $Y=1.542 $X2=0
+ $Y2=0
cc_564 N_A_418_74#_c_585_n N_COUT_c_1530_n 0.00208787f $X=9.085 $Y=1.765 $X2=0
+ $Y2=0
cc_565 N_A_418_74#_c_586_n N_COUT_c_1530_n 6.83942e-19 $X=9.535 $Y=1.765 $X2=0
+ $Y2=0
cc_566 N_A_418_74#_c_764_p N_COUT_c_1530_n 0.0276944f $X=9.84 $Y=1.485 $X2=0
+ $Y2=0
cc_567 N_A_418_74#_c_583_n N_COUT_c_1530_n 0.00808948f $X=10.485 $Y=1.542 $X2=0
+ $Y2=0
cc_568 N_A_418_74#_c_585_n N_COUT_c_1531_n 0.0104444f $X=9.085 $Y=1.765 $X2=0
+ $Y2=0
cc_569 N_A_418_74#_c_586_n N_COUT_c_1531_n 0.0125507f $X=9.535 $Y=1.765 $X2=0
+ $Y2=0
cc_570 N_A_418_74#_c_587_n N_COUT_c_1531_n 7.34595e-19 $X=10.035 $Y=1.765 $X2=0
+ $Y2=0
cc_571 N_A_418_74#_M1013_g N_COUT_c_1526_n 0.00852713f $X=9.255 $Y=0.78 $X2=0
+ $Y2=0
cc_572 N_A_418_74#_M1014_g N_COUT_c_1526_n 3.13308e-19 $X=9.685 $Y=0.78 $X2=0
+ $Y2=0
cc_573 N_A_418_74#_c_586_n N_COUT_c_1532_n 0.0122806f $X=9.535 $Y=1.765 $X2=0
+ $Y2=0
cc_574 N_A_418_74#_c_587_n N_COUT_c_1532_n 0.014256f $X=10.035 $Y=1.765 $X2=0
+ $Y2=0
cc_575 N_A_418_74#_c_764_p N_COUT_c_1532_n 0.0355356f $X=9.84 $Y=1.485 $X2=0
+ $Y2=0
cc_576 N_A_418_74#_c_583_n N_COUT_c_1532_n 0.00898226f $X=10.485 $Y=1.542 $X2=0
+ $Y2=0
cc_577 N_A_418_74#_M1014_g N_COUT_c_1548_n 0.0122129f $X=9.685 $Y=0.78 $X2=0
+ $Y2=0
cc_578 N_A_418_74#_M1022_g N_COUT_c_1548_n 0.0128537f $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_579 N_A_418_74#_c_764_p N_COUT_c_1548_n 0.0250701f $X=9.84 $Y=1.485 $X2=0
+ $Y2=0
cc_580 N_A_418_74#_c_583_n N_COUT_c_1548_n 0.00224919f $X=10.485 $Y=1.542 $X2=0
+ $Y2=0
cc_581 N_A_418_74#_M1013_g N_COUT_c_1527_n 0.00211285f $X=9.255 $Y=0.78 $X2=0
+ $Y2=0
cc_582 N_A_418_74#_c_764_p N_COUT_c_1527_n 0.0178863f $X=9.84 $Y=1.485 $X2=0
+ $Y2=0
cc_583 N_A_418_74#_c_583_n N_COUT_c_1527_n 0.00258765f $X=10.485 $Y=1.542 $X2=0
+ $Y2=0
cc_584 N_A_418_74#_M1014_g N_COUT_c_1528_n 6.05373e-19 $X=9.685 $Y=0.78 $X2=0
+ $Y2=0
cc_585 N_A_418_74#_M1022_g N_COUT_c_1528_n 0.00849808f $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_586 N_A_418_74#_M1035_g N_COUT_c_1528_n 4.03226e-19 $X=10.545 $Y=0.78 $X2=0
+ $Y2=0
cc_587 N_A_418_74#_M1014_g N_COUT_c_1529_n 8.24123e-19 $X=9.685 $Y=0.78 $X2=0
+ $Y2=0
cc_588 N_A_418_74#_M1022_g N_COUT_c_1529_n 0.00456448f $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_589 N_A_418_74#_M1035_g N_COUT_c_1529_n 0.00407331f $X=10.545 $Y=0.78 $X2=0
+ $Y2=0
cc_590 N_A_418_74#_c_764_p N_COUT_c_1529_n 0.0151308f $X=9.84 $Y=1.485 $X2=0
+ $Y2=0
cc_591 N_A_418_74#_c_583_n N_COUT_c_1529_n 0.0208906f $X=10.485 $Y=1.542 $X2=0
+ $Y2=0
cc_592 N_A_418_74#_M1022_g N_COUT_c_1563_n 3.84191e-19 $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_593 N_A_418_74#_c_587_n N_COUT_c_1533_n 0.00234056f $X=10.035 $Y=1.765 $X2=0
+ $Y2=0
cc_594 N_A_418_74#_c_588_n N_COUT_c_1533_n 0.00498446f $X=10.485 $Y=1.765 $X2=0
+ $Y2=0
cc_595 N_A_418_74#_c_764_p N_COUT_c_1533_n 0.0066008f $X=9.84 $Y=1.485 $X2=0
+ $Y2=0
cc_596 N_A_418_74#_c_583_n N_COUT_c_1533_n 0.0258883f $X=10.485 $Y=1.542 $X2=0
+ $Y2=0
cc_597 N_A_418_74#_c_586_n COUT 6.34305e-19 $X=9.535 $Y=1.765 $X2=0 $Y2=0
cc_598 N_A_418_74#_c_587_n COUT 0.0119706f $X=10.035 $Y=1.765 $X2=0 $Y2=0
cc_599 N_A_418_74#_c_588_n COUT 0.0121646f $X=10.485 $Y=1.765 $X2=0 $Y2=0
cc_600 N_A_418_74#_c_638_n N_A_27_74#_M1026_d 0.00228734f $X=2.135 $Y=0.925
+ $X2=0 $Y2=0
cc_601 N_A_418_74#_c_622_n N_A_27_74#_M1026_d 0.00356839f $X=1.835 $Y=0.965
+ $X2=0 $Y2=0
cc_602 N_A_418_74#_c_577_n N_A_27_74#_c_1595_n 0.0140589f $X=2.3 $Y=0.515 $X2=0
+ $Y2=0
cc_603 N_A_418_74#_c_619_n N_A_27_74#_c_1595_n 0.00782456f $X=1.665 $Y=0.965
+ $X2=0 $Y2=0
cc_604 N_A_418_74#_c_622_n N_A_27_74#_c_1595_n 0.0142648f $X=1.835 $Y=0.965
+ $X2=0 $Y2=0
cc_605 N_A_418_74#_c_669_p N_A_27_74#_c_1596_n 0.00503853f $X=1.175 $Y=1.005
+ $X2=0 $Y2=0
cc_606 N_A_418_74#_c_669_p N_A_27_74#_c_1599_n 0.013831f $X=1.175 $Y=1.005 $X2=0
+ $Y2=0
cc_607 N_A_418_74#_c_619_n N_A_27_74#_c_1599_n 0.0207538f $X=1.665 $Y=0.965
+ $X2=0 $Y2=0
cc_608 N_A_418_74#_c_576_n N_VGND_M1032_d 5.28288e-19 $X=1.09 $Y=1.745 $X2=-0.19
+ $Y2=-0.245
cc_609 N_A_418_74#_c_669_p N_VGND_M1032_d 0.00604059f $X=1.175 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_610 N_A_418_74#_c_619_n N_VGND_M1032_d 0.00740987f $X=1.665 $Y=0.965
+ $X2=-0.19 $Y2=-0.245
cc_611 N_A_418_74#_c_626_n N_VGND_M1033_d 0.00278732f $X=3.385 $Y=0.965 $X2=0
+ $Y2=0
cc_612 N_A_418_74#_c_629_n N_VGND_M1033_d 0.00256535f $X=3.555 $Y=0.965 $X2=0
+ $Y2=0
cc_613 N_A_418_74#_c_606_n N_VGND_M1030_d 0.00849548f $X=4.93 $Y=1.005 $X2=0
+ $Y2=0
cc_614 N_A_418_74#_c_683_p N_VGND_M1039_d 0.007557f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_615 N_A_418_74#_c_683_p N_VGND_M1021_d 0.00726636f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_616 N_A_418_74#_c_683_p N_VGND_M1036_d 0.0116153f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_617 N_A_418_74#_c_580_n N_VGND_M1036_d 0.00806651f $X=9.05 $Y=1.32 $X2=0
+ $Y2=0
cc_618 N_A_418_74#_c_626_n N_VGND_c_1627_n 0.0176682f $X=3.385 $Y=0.965 $X2=0
+ $Y2=0
cc_619 N_A_418_74#_M1013_g N_VGND_c_1628_n 4.88565e-19 $X=9.255 $Y=0.78 $X2=0
+ $Y2=0
cc_620 N_A_418_74#_M1014_g N_VGND_c_1628_n 0.00879111f $X=9.685 $Y=0.78 $X2=0
+ $Y2=0
cc_621 N_A_418_74#_M1022_g N_VGND_c_1628_n 0.00176539f $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_622 N_A_418_74#_M1022_g N_VGND_c_1630_n 5.99782e-19 $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_623 N_A_418_74#_M1035_g N_VGND_c_1630_n 0.0157698f $X=10.545 $Y=0.78 $X2=0
+ $Y2=0
cc_624 N_A_418_74#_c_577_n N_VGND_c_1631_n 0.0146038f $X=2.3 $Y=0.515 $X2=0
+ $Y2=0
cc_625 N_A_418_74#_c_579_n N_VGND_c_1633_n 0.00302543f $X=5.255 $Y=0.34 $X2=0
+ $Y2=0
cc_626 N_A_418_74#_c_570_n N_VGND_c_1635_n 0.00418685f $X=5.045 $Y=1.22 $X2=0
+ $Y2=0
cc_627 N_A_418_74#_c_578_n N_VGND_c_1635_n 0.0753865f $X=6.255 $Y=0.34 $X2=0
+ $Y2=0
cc_628 N_A_418_74#_c_579_n N_VGND_c_1635_n 0.0120637f $X=5.255 $Y=0.34 $X2=0
+ $Y2=0
cc_629 N_A_418_74#_c_683_p N_VGND_c_1635_n 0.00540182f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_630 N_A_418_74#_c_683_p N_VGND_c_1636_n 0.0114147f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_631 N_A_418_74#_c_683_p N_VGND_c_1637_n 0.0114147f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_632 N_A_418_74#_M1013_g N_VGND_c_1638_n 0.00523933f $X=9.255 $Y=0.78 $X2=0
+ $Y2=0
cc_633 N_A_418_74#_M1014_g N_VGND_c_1638_n 0.00455951f $X=9.685 $Y=0.78 $X2=0
+ $Y2=0
cc_634 N_A_418_74#_M1022_g N_VGND_c_1639_n 0.00523933f $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_635 N_A_418_74#_M1035_g N_VGND_c_1639_n 0.00455951f $X=10.545 $Y=0.78 $X2=0
+ $Y2=0
cc_636 N_A_418_74#_c_578_n N_VGND_c_1642_n 0.00746752f $X=6.255 $Y=0.34 $X2=0
+ $Y2=0
cc_637 N_A_418_74#_c_683_p N_VGND_c_1642_n 0.0244407f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_638 N_A_418_74#_c_683_p N_VGND_c_1643_n 0.0244835f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_639 N_A_418_74#_M1013_g N_VGND_c_1644_n 0.00192643f $X=9.255 $Y=0.78 $X2=0
+ $Y2=0
cc_640 N_A_418_74#_c_683_p N_VGND_c_1644_n 0.0256831f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_641 N_A_418_74#_c_570_n N_VGND_c_1646_n 0.0078168f $X=5.045 $Y=1.22 $X2=0
+ $Y2=0
cc_642 N_A_418_74#_M1013_g N_VGND_c_1646_n 0.00533081f $X=9.255 $Y=0.78 $X2=0
+ $Y2=0
cc_643 N_A_418_74#_M1014_g N_VGND_c_1646_n 0.00447788f $X=9.685 $Y=0.78 $X2=0
+ $Y2=0
cc_644 N_A_418_74#_M1022_g N_VGND_c_1646_n 0.00533081f $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_645 N_A_418_74#_M1035_g N_VGND_c_1646_n 0.00447788f $X=10.545 $Y=0.78 $X2=0
+ $Y2=0
cc_646 N_A_418_74#_c_577_n N_VGND_c_1646_n 0.0121018f $X=2.3 $Y=0.515 $X2=0
+ $Y2=0
cc_647 N_A_418_74#_c_578_n N_VGND_c_1646_n 0.04278f $X=6.255 $Y=0.34 $X2=0 $Y2=0
cc_648 N_A_418_74#_c_579_n N_VGND_c_1646_n 0.00644906f $X=5.255 $Y=0.34 $X2=0
+ $Y2=0
cc_649 N_A_418_74#_c_683_p N_VGND_c_1646_n 0.0551926f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_650 N_A_418_74#_c_622_n N_VGND_c_1646_n 0.00539663f $X=1.835 $Y=0.965 $X2=0
+ $Y2=0
cc_651 N_A_418_74#_c_626_n N_VGND_c_1646_n 0.0236322f $X=3.385 $Y=0.965 $X2=0
+ $Y2=0
cc_652 N_A_418_74#_c_629_n N_VGND_c_1646_n 0.00156853f $X=3.555 $Y=0.965 $X2=0
+ $Y2=0
cc_653 N_A_418_74#_c_626_n A_532_74# 0.00912043f $X=3.385 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_654 N_A_418_74#_c_606_n N_A_734_74#_M1027_d 0.00443657f $X=4.93 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_655 N_A_418_74#_c_606_n N_A_734_74#_M1015_d 0.00451688f $X=4.93 $Y=1.005
+ $X2=0 $Y2=0
cc_656 N_A_418_74#_c_606_n N_A_734_74#_c_1776_n 0.0390509f $X=4.93 $Y=1.005
+ $X2=0 $Y2=0
cc_657 N_A_418_74#_c_606_n N_A_734_74#_c_1774_n 0.0140929f $X=4.93 $Y=1.005
+ $X2=0 $Y2=0
cc_658 N_A_418_74#_c_606_n N_A_734_74#_c_1775_n 0.0140929f $X=4.93 $Y=1.005
+ $X2=0 $Y2=0
cc_659 N_A_418_74#_c_579_n N_A_734_74#_c_1775_n 0.00392045f $X=5.255 $Y=0.34
+ $X2=0 $Y2=0
cc_660 N_A_418_74#_c_578_n A_1160_74# 0.00206111f $X=6.255 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_661 N_A_418_74#_c_578_n A_1238_74# 8.72382e-19 $X=6.255 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_662 N_A_418_74#_c_613_n A_1238_74# 0.00341292f $X=6.34 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_663 N_A_418_74#_c_683_p A_1238_74# 0.00180488f $X=8.965 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_664 N_A_418_74#_c_614_n A_1238_74# 0.0049852f $X=6.425 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_665 N_A_M1012_g N_A_1024_74#_c_1072_n 0.0191394f $X=6.64 $Y=2.34 $X2=0 $Y2=0
cc_666 N_A_c_897_n N_A_1024_74#_c_1072_n 0.00354341f $X=6.64 $Y=3.15 $X2=0 $Y2=0
cc_667 N_A_M1039_g N_A_1024_74#_M1020_g 0.025914f $X=6.625 $Y=0.74 $X2=0 $Y2=0
cc_668 N_A_M1039_g N_A_1024_74#_c_1084_n 0.0149876f $X=6.625 $Y=0.74 $X2=0 $Y2=0
cc_669 N_A_M1012_g N_A_1024_74#_c_1087_n 0.0185584f $X=6.64 $Y=2.34 $X2=0 $Y2=0
cc_670 N_A_M1039_g N_A_1024_74#_c_1068_n 0.00444019f $X=6.625 $Y=0.74 $X2=0
+ $Y2=0
cc_671 N_A_c_870_n N_A_1024_74#_c_1076_n 7.63821e-19 $X=6.64 $Y=1.765 $X2=0
+ $Y2=0
cc_672 N_A_M1012_g N_A_1024_74#_c_1076_n 0.00372133f $X=6.64 $Y=2.34 $X2=0 $Y2=0
cc_673 N_A_c_891_n N_A_1024_74#_c_1078_n 0.00640339f $X=6.55 $Y=3.15 $X2=0 $Y2=0
cc_674 N_A_M1039_g N_A_1024_74#_c_1093_n 3.84346e-19 $X=6.625 $Y=0.74 $X2=0
+ $Y2=0
cc_675 N_A_M1012_g N_A_1024_74#_c_1095_n 0.00276802f $X=6.64 $Y=2.34 $X2=0 $Y2=0
cc_676 N_A_M1039_g N_A_1024_74#_c_1070_n 0.0031874f $X=6.625 $Y=0.74 $X2=0 $Y2=0
cc_677 N_A_c_870_n N_A_1024_74#_c_1070_n 5.25256e-19 $X=6.64 $Y=1.765 $X2=0
+ $Y2=0
cc_678 N_A_M1039_g N_A_1024_74#_c_1071_n 0.00698694f $X=6.625 $Y=0.74 $X2=0
+ $Y2=0
cc_679 N_A_c_870_n N_A_1024_74#_c_1071_n 0.00393277f $X=6.64 $Y=1.765 $X2=0
+ $Y2=0
cc_680 N_A_c_876_n N_A_27_392#_c_1223_n 4.59984e-19 $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_681 N_A_M1028_g N_A_27_392#_c_1223_n 0.00345041f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_682 A N_A_27_392#_c_1223_n 0.02912f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_683 N_A_c_874_n N_A_27_392#_c_1223_n 0.00143639f $X=0.63 $Y=1.41 $X2=0 $Y2=0
cc_684 N_A_M1028_g N_A_27_392#_c_1224_n 0.00941971f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_685 N_A_c_879_n N_A_27_392#_c_1224_n 3.90045e-19 $X=0.595 $Y=3.15 $X2=0 $Y2=0
cc_686 N_A_M1028_g N_A_27_392#_c_1232_n 0.0135162f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_687 A N_A_27_392#_c_1232_n 0.0184533f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_688 N_A_c_874_n N_A_27_392#_c_1232_n 7.65965e-19 $X=0.63 $Y=1.41 $X2=0 $Y2=0
cc_689 N_A_M1028_g N_A_27_392#_c_1233_n 0.00146175f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_690 N_A_c_878_n N_A_27_392#_c_1225_n 0.00284623f $X=3.02 $Y=3.15 $X2=0 $Y2=0
cc_691 N_A_c_878_n N_A_27_392#_c_1226_n 0.0179795f $X=3.02 $Y=3.15 $X2=0 $Y2=0
cc_692 A N_VPWR_M1028_d 7.01028e-19 $X=0.635 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_693 N_A_M1028_g N_VPWR_c_1275_n 0.00655954f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_694 N_A_c_878_n N_VPWR_c_1275_n 0.0165008f $X=3.02 $Y=3.15 $X2=0 $Y2=0
cc_695 N_A_c_879_n N_VPWR_c_1275_n 0.00159376f $X=0.595 $Y=3.15 $X2=0 $Y2=0
cc_696 N_A_c_881_n N_VPWR_c_1276_n 0.00437861f $X=3.11 $Y=2.9 $X2=0 $Y2=0
cc_697 N_A_c_882_n N_VPWR_c_1276_n 0.0111301f $X=3.11 $Y=3.075 $X2=0 $Y2=0
cc_698 N_A_M1001_g N_VPWR_c_1276_n 0.0149631f $X=3.11 $Y=2.235 $X2=0 $Y2=0
cc_699 N_A_c_885_n N_VPWR_c_1276_n 0.0177656f $X=4.54 $Y=3.15 $X2=0 $Y2=0
cc_700 N_A_c_895_n N_VPWR_c_1276_n 0.00476669f $X=3.11 $Y=3.15 $X2=0 $Y2=0
cc_701 N_A_c_885_n N_VPWR_c_1277_n 0.021565f $X=4.54 $Y=3.15 $X2=0 $Y2=0
cc_702 N_A_c_887_n N_VPWR_c_1277_n 0.004539f $X=4.63 $Y=2.9 $X2=0 $Y2=0
cc_703 N_A_c_888_n N_VPWR_c_1277_n 0.0114653f $X=4.63 $Y=3.075 $X2=0 $Y2=0
cc_704 N_A_M1004_g N_VPWR_c_1277_n 0.00541968f $X=4.63 $Y=2.235 $X2=0 $Y2=0
cc_705 N_A_c_896_n N_VPWR_c_1277_n 0.00477316f $X=4.63 $Y=3.15 $X2=0 $Y2=0
cc_706 N_A_M1012_g N_VPWR_c_1278_n 0.0164201f $X=6.64 $Y=2.34 $X2=0 $Y2=0
cc_707 N_A_c_897_n N_VPWR_c_1278_n 0.00967347f $X=6.64 $Y=3.15 $X2=0 $Y2=0
cc_708 N_A_c_878_n N_VPWR_c_1284_n 0.065989f $X=3.02 $Y=3.15 $X2=0 $Y2=0
cc_709 N_A_c_885_n N_VPWR_c_1286_n 0.0199069f $X=4.54 $Y=3.15 $X2=0 $Y2=0
cc_710 N_A_c_896_n N_VPWR_c_1287_n 0.0699233f $X=4.63 $Y=3.15 $X2=0 $Y2=0
cc_711 N_A_c_879_n N_VPWR_c_1292_n 0.0082546f $X=0.595 $Y=3.15 $X2=0 $Y2=0
cc_712 N_A_c_878_n N_VPWR_c_1274_n 0.0758349f $X=3.02 $Y=3.15 $X2=0 $Y2=0
cc_713 N_A_c_879_n N_VPWR_c_1274_n 0.0116723f $X=0.595 $Y=3.15 $X2=0 $Y2=0
cc_714 N_A_c_885_n N_VPWR_c_1274_n 0.0207512f $X=4.54 $Y=3.15 $X2=0 $Y2=0
cc_715 N_A_c_891_n N_VPWR_c_1274_n 0.071722f $X=6.55 $Y=3.15 $X2=0 $Y2=0
cc_716 N_A_c_895_n N_VPWR_c_1274_n 0.00895426f $X=3.11 $Y=3.15 $X2=0 $Y2=0
cc_717 N_A_c_896_n N_VPWR_c_1274_n 0.00895426f $X=4.63 $Y=3.15 $X2=0 $Y2=0
cc_718 N_A_c_897_n N_VPWR_c_1274_n 0.0131297f $X=6.64 $Y=3.15 $X2=0 $Y2=0
cc_719 N_A_M1004_g N_A_737_347#_c_1431_n 0.0157099f $X=4.63 $Y=2.235 $X2=0 $Y2=0
cc_720 N_A_M1004_g N_A_737_347#_c_1427_n 0.00272481f $X=4.63 $Y=2.235 $X2=0
+ $Y2=0
cc_721 N_A_c_891_n N_A_737_347#_c_1427_n 0.00638811f $X=6.55 $Y=3.15 $X2=0 $Y2=0
cc_722 N_A_c_885_n N_A_737_347#_c_1428_n 0.00614494f $X=4.54 $Y=3.15 $X2=0 $Y2=0
cc_723 N_A_M1004_g N_A_737_347#_c_1428_n 7.61724e-19 $X=4.63 $Y=2.235 $X2=0
+ $Y2=0
cc_724 N_A_M1012_g N_SUM_c_1467_n 9.96836e-19 $X=6.64 $Y=2.34 $X2=0 $Y2=0
cc_725 N_A_M1032_g N_A_27_74#_c_1596_n 0.0205742f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_726 A N_A_27_74#_c_1596_n 0.0246165f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_727 N_A_c_874_n N_A_27_74#_c_1596_n 0.00671505f $X=0.63 $Y=1.41 $X2=0 $Y2=0
cc_728 N_A_M1032_g N_A_27_74#_c_1599_n 0.0120858f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_729 A N_A_27_74#_c_1599_n 0.0119709f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_730 N_A_c_874_n N_A_27_74#_c_1599_n 0.00383117f $X=0.63 $Y=1.41 $X2=0 $Y2=0
cc_731 N_A_c_871_n N_VGND_c_1627_n 0.010869f $X=3.11 $Y=1.185 $X2=0 $Y2=0
cc_732 N_A_c_871_n N_VGND_c_1631_n 0.00383152f $X=3.11 $Y=1.185 $X2=0 $Y2=0
cc_733 N_A_c_872_n N_VGND_c_1633_n 0.0023296f $X=4.63 $Y=1.185 $X2=0 $Y2=0
cc_734 N_A_M1039_g N_VGND_c_1635_n 0.00320129f $X=6.625 $Y=0.74 $X2=0 $Y2=0
cc_735 N_A_c_872_n N_VGND_c_1635_n 0.00316493f $X=4.63 $Y=1.185 $X2=0 $Y2=0
cc_736 N_A_M1032_g N_VGND_c_1640_n 0.00316493f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_737 N_A_M1032_g N_VGND_c_1641_n 0.00608124f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_738 N_A_M1039_g N_VGND_c_1642_n 0.00253998f $X=6.625 $Y=0.74 $X2=0 $Y2=0
cc_739 N_A_M1032_g N_VGND_c_1646_n 0.00400459f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_740 N_A_M1039_g N_VGND_c_1646_n 0.00405511f $X=6.625 $Y=0.74 $X2=0 $Y2=0
cc_741 N_A_c_871_n N_VGND_c_1646_n 0.00384996f $X=3.11 $Y=1.185 $X2=0 $Y2=0
cc_742 N_A_c_872_n N_VGND_c_1646_n 0.00393316f $X=4.63 $Y=1.185 $X2=0 $Y2=0
cc_743 N_A_c_872_n N_A_734_74#_c_1776_n 0.00936301f $X=4.63 $Y=1.185 $X2=0 $Y2=0
cc_744 N_A_c_872_n N_A_734_74#_c_1774_n 8.6409e-19 $X=4.63 $Y=1.185 $X2=0 $Y2=0
cc_745 N_A_c_872_n N_A_734_74#_c_1775_n 0.0057442f $X=4.63 $Y=1.185 $X2=0 $Y2=0
cc_746 N_A_1024_74#_c_1087_n N_VPWR_M1012_d 0.0105098f $X=6.905 $Y=2.035 $X2=0
+ $Y2=0
cc_747 N_A_1024_74#_c_1076_n N_VPWR_M1012_d 0.00209989f $X=6.99 $Y=1.95 $X2=0
+ $Y2=0
cc_748 N_A_1024_74#_c_1072_n N_VPWR_c_1278_n 0.00538964f $X=7.185 $Y=1.765 $X2=0
+ $Y2=0
cc_749 N_A_1024_74#_c_1087_n N_VPWR_c_1278_n 0.021319f $X=6.905 $Y=2.035 $X2=0
+ $Y2=0
cc_750 N_A_1024_74#_c_1073_n N_VPWR_c_1279_n 0.00612247f $X=7.635 $Y=1.765 $X2=0
+ $Y2=0
cc_751 N_A_1024_74#_c_1074_n N_VPWR_c_1279_n 0.00729593f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_752 N_A_1024_74#_c_1075_n N_VPWR_c_1280_n 0.00731086f $X=8.585 $Y=1.765 $X2=0
+ $Y2=0
cc_753 N_A_1024_74#_c_1071_n N_VPWR_c_1280_n 5.712e-19 $X=8.585 $Y=1.552 $X2=0
+ $Y2=0
cc_754 N_A_1024_74#_c_1078_n N_VPWR_c_1287_n 0.00753052f $X=5.405 $Y=2.145 $X2=0
+ $Y2=0
cc_755 N_A_1024_74#_c_1072_n N_VPWR_c_1288_n 0.00445602f $X=7.185 $Y=1.765 $X2=0
+ $Y2=0
cc_756 N_A_1024_74#_c_1073_n N_VPWR_c_1288_n 0.00445602f $X=7.635 $Y=1.765 $X2=0
+ $Y2=0
cc_757 N_A_1024_74#_c_1074_n N_VPWR_c_1289_n 0.00445602f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_758 N_A_1024_74#_c_1075_n N_VPWR_c_1289_n 0.00445602f $X=8.585 $Y=1.765 $X2=0
+ $Y2=0
cc_759 N_A_1024_74#_c_1072_n N_VPWR_c_1274_n 0.00858344f $X=7.185 $Y=1.765 $X2=0
+ $Y2=0
cc_760 N_A_1024_74#_c_1073_n N_VPWR_c_1274_n 0.0085805f $X=7.635 $Y=1.765 $X2=0
+ $Y2=0
cc_761 N_A_1024_74#_c_1074_n N_VPWR_c_1274_n 0.00857378f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_762 N_A_1024_74#_c_1075_n N_VPWR_c_1274_n 0.00858104f $X=8.585 $Y=1.765 $X2=0
+ $Y2=0
cc_763 N_A_1024_74#_c_1078_n N_VPWR_c_1274_n 0.00909433f $X=5.405 $Y=2.145 $X2=0
+ $Y2=0
cc_764 N_A_1024_74#_c_1078_n N_A_737_347#_c_1427_n 0.0195142f $X=5.405 $Y=2.145
+ $X2=0 $Y2=0
cc_765 N_A_1024_74#_c_1081_n A_1141_347# 0.0100099f $X=6.255 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_766 N_A_1024_74#_c_1081_n A_1235_347# 0.00157041f $X=6.255 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_767 N_A_1024_74#_c_1087_n A_1235_347# 0.00446616f $X=6.905 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_768 N_A_1024_74#_c_1095_n A_1235_347# 0.0122459f $X=6.34 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_769 N_A_1024_74#_c_1072_n N_SUM_c_1466_n 0.00183202f $X=7.185 $Y=1.765 $X2=0
+ $Y2=0
cc_770 N_A_1024_74#_c_1073_n N_SUM_c_1466_n 4.27055e-19 $X=7.635 $Y=1.765 $X2=0
+ $Y2=0
cc_771 N_A_1024_74#_c_1069_n N_SUM_c_1466_n 0.0219683f $X=7.94 $Y=1.505 $X2=0
+ $Y2=0
cc_772 N_A_1024_74#_c_1071_n N_SUM_c_1466_n 0.00670438f $X=8.585 $Y=1.552 $X2=0
+ $Y2=0
cc_773 N_A_1024_74#_c_1072_n N_SUM_c_1467_n 0.0121826f $X=7.185 $Y=1.765 $X2=0
+ $Y2=0
cc_774 N_A_1024_74#_c_1073_n N_SUM_c_1467_n 0.0120909f $X=7.635 $Y=1.765 $X2=0
+ $Y2=0
cc_775 N_A_1024_74#_c_1074_n N_SUM_c_1467_n 7.29241e-19 $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_776 N_A_1024_74#_M1020_g N_SUM_c_1463_n 0.0035804f $X=7.215 $Y=0.78 $X2=0
+ $Y2=0
cc_777 N_A_1024_74#_M1021_g N_SUM_c_1463_n 0.0120038f $X=7.645 $Y=0.78 $X2=0
+ $Y2=0
cc_778 N_A_1024_74#_M1034_g N_SUM_c_1463_n 0.0121154f $X=8.235 $Y=0.78 $X2=0
+ $Y2=0
cc_779 N_A_1024_74#_c_1084_n N_SUM_c_1463_n 0.0135437f $X=6.905 $Y=1.005 $X2=0
+ $Y2=0
cc_780 N_A_1024_74#_c_1068_n N_SUM_c_1463_n 0.00568635f $X=6.99 $Y=1.34 $X2=0
+ $Y2=0
cc_781 N_A_1024_74#_c_1069_n N_SUM_c_1463_n 0.064353f $X=7.94 $Y=1.505 $X2=0
+ $Y2=0
cc_782 N_A_1024_74#_c_1071_n N_SUM_c_1463_n 0.0082022f $X=8.585 $Y=1.552 $X2=0
+ $Y2=0
cc_783 N_A_1024_74#_c_1073_n N_SUM_c_1494_n 0.0122806f $X=7.635 $Y=1.765 $X2=0
+ $Y2=0
cc_784 N_A_1024_74#_c_1074_n N_SUM_c_1494_n 0.0135926f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_785 N_A_1024_74#_c_1069_n N_SUM_c_1494_n 0.0345236f $X=7.94 $Y=1.505 $X2=0
+ $Y2=0
cc_786 N_A_1024_74#_c_1071_n N_SUM_c_1494_n 0.00732518f $X=8.585 $Y=1.552 $X2=0
+ $Y2=0
cc_787 N_A_1024_74#_M1034_g N_SUM_c_1464_n 0.00114171f $X=8.235 $Y=0.78 $X2=0
+ $Y2=0
cc_788 N_A_1024_74#_M1036_g N_SUM_c_1464_n 0.00537066f $X=8.665 $Y=0.78 $X2=0
+ $Y2=0
cc_789 N_A_1024_74#_M1021_g N_SUM_c_1465_n 7.63771e-19 $X=7.645 $Y=0.78 $X2=0
+ $Y2=0
cc_790 N_A_1024_74#_c_1074_n N_SUM_c_1465_n 0.00185393f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_791 N_A_1024_74#_M1034_g N_SUM_c_1465_n 0.00486056f $X=8.235 $Y=0.78 $X2=0
+ $Y2=0
cc_792 N_A_1024_74#_c_1075_n N_SUM_c_1465_n 0.00186427f $X=8.585 $Y=1.765 $X2=0
+ $Y2=0
cc_793 N_A_1024_74#_M1036_g N_SUM_c_1465_n 0.00183896f $X=8.665 $Y=0.78 $X2=0
+ $Y2=0
cc_794 N_A_1024_74#_c_1069_n N_SUM_c_1465_n 0.0244401f $X=7.94 $Y=1.505 $X2=0
+ $Y2=0
cc_795 N_A_1024_74#_c_1071_n N_SUM_c_1465_n 0.0298955f $X=8.585 $Y=1.552 $X2=0
+ $Y2=0
cc_796 N_A_1024_74#_c_1074_n SUM 6.21797e-19 $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_797 N_A_1024_74#_c_1075_n SUM 0.00174826f $X=8.585 $Y=1.765 $X2=0 $Y2=0
cc_798 N_A_1024_74#_c_1071_n SUM 0.00163026f $X=8.585 $Y=1.552 $X2=0 $Y2=0
cc_799 N_A_1024_74#_c_1073_n SUM 6.2994e-19 $X=7.635 $Y=1.765 $X2=0 $Y2=0
cc_800 N_A_1024_74#_c_1074_n SUM 0.011525f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_801 N_A_1024_74#_c_1075_n SUM 0.0106842f $X=8.585 $Y=1.765 $X2=0 $Y2=0
cc_802 N_A_1024_74#_M1036_g N_COUT_c_1526_n 9.32329e-19 $X=8.665 $Y=0.78 $X2=0
+ $Y2=0
cc_803 N_A_1024_74#_c_1084_n N_VGND_M1039_d 0.0123197f $X=6.905 $Y=1.005 $X2=0
+ $Y2=0
cc_804 N_A_1024_74#_c_1068_n N_VGND_M1039_d 0.00175048f $X=6.99 $Y=1.34 $X2=0
+ $Y2=0
cc_805 N_A_1024_74#_M1020_g N_VGND_c_1636_n 0.00414982f $X=7.215 $Y=0.78 $X2=0
+ $Y2=0
cc_806 N_A_1024_74#_M1021_g N_VGND_c_1636_n 0.00414982f $X=7.645 $Y=0.78 $X2=0
+ $Y2=0
cc_807 N_A_1024_74#_M1034_g N_VGND_c_1637_n 0.00414982f $X=8.235 $Y=0.78 $X2=0
+ $Y2=0
cc_808 N_A_1024_74#_M1036_g N_VGND_c_1637_n 0.00414982f $X=8.665 $Y=0.78 $X2=0
+ $Y2=0
cc_809 N_A_1024_74#_M1020_g N_VGND_c_1642_n 0.00378066f $X=7.215 $Y=0.78 $X2=0
+ $Y2=0
cc_810 N_A_1024_74#_M1021_g N_VGND_c_1643_n 0.00378066f $X=7.645 $Y=0.78 $X2=0
+ $Y2=0
cc_811 N_A_1024_74#_M1034_g N_VGND_c_1643_n 0.00378066f $X=8.235 $Y=0.78 $X2=0
+ $Y2=0
cc_812 N_A_1024_74#_M1036_g N_VGND_c_1644_n 0.00378066f $X=8.665 $Y=0.78 $X2=0
+ $Y2=0
cc_813 N_A_1024_74#_M1020_g N_VGND_c_1646_n 0.00533081f $X=7.215 $Y=0.78 $X2=0
+ $Y2=0
cc_814 N_A_1024_74#_M1021_g N_VGND_c_1646_n 0.00533081f $X=7.645 $Y=0.78 $X2=0
+ $Y2=0
cc_815 N_A_1024_74#_M1034_g N_VGND_c_1646_n 0.00533081f $X=8.235 $Y=0.78 $X2=0
+ $Y2=0
cc_816 N_A_1024_74#_M1036_g N_VGND_c_1646_n 0.00533081f $X=8.665 $Y=0.78 $X2=0
+ $Y2=0
cc_817 N_A_1024_74#_c_1104_n A_1160_74# 0.00308137f $X=5.915 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_818 N_A_1024_74#_c_1093_n A_1160_74# 0.00302066f $X=6.085 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_819 N_A_1024_74#_c_1084_n A_1238_74# 0.00608853f $X=6.905 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_820 N_A_27_392#_c_1232_n N_VPWR_M1028_d 0.0191384f $X=0.985 $Y=2.17 $X2=-0.19
+ $Y2=1.66
cc_821 N_A_27_392#_c_1233_n N_VPWR_M1028_d 0.00424793f $X=1.07 $Y=2.63 $X2=-0.19
+ $Y2=1.66
cc_822 N_A_27_392#_c_1225_n N_VPWR_M1028_d 0.00100166f $X=1.155 $Y=2.795
+ $X2=-0.19 $Y2=1.66
cc_823 N_A_27_392#_c_1224_n N_VPWR_c_1275_n 0.0361783f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_824 N_A_27_392#_c_1232_n N_VPWR_c_1275_n 0.0136682f $X=0.985 $Y=2.17 $X2=0
+ $Y2=0
cc_825 N_A_27_392#_c_1233_n N_VPWR_c_1275_n 0.0148534f $X=1.07 $Y=2.63 $X2=0
+ $Y2=0
cc_826 N_A_27_392#_c_1225_n N_VPWR_c_1275_n 0.0272461f $X=1.155 $Y=2.795 $X2=0
+ $Y2=0
cc_827 N_A_27_392#_c_1225_n N_VPWR_c_1284_n 0.00701426f $X=1.155 $Y=2.795 $X2=0
+ $Y2=0
cc_828 N_A_27_392#_c_1226_n N_VPWR_c_1284_n 0.0331696f $X=1.84 $Y=2.795 $X2=0
+ $Y2=0
cc_829 N_A_27_392#_c_1224_n N_VPWR_c_1292_n 0.0145932f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_830 N_A_27_392#_c_1224_n N_VPWR_c_1274_n 0.0119865f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_831 N_A_27_392#_c_1225_n N_VPWR_c_1274_n 0.00552059f $X=1.155 $Y=2.795 $X2=0
+ $Y2=0
cc_832 N_A_27_392#_c_1226_n N_VPWR_c_1274_n 0.0268277f $X=1.84 $Y=2.795 $X2=0
+ $Y2=0
cc_833 N_VPWR_M1003_d N_A_737_347#_c_1431_n 0.00696341f $X=4.135 $Y=1.735 $X2=0
+ $Y2=0
cc_834 N_VPWR_c_1277_n N_A_737_347#_c_1431_n 0.02592f $X=4.37 $Y=2.59 $X2=0
+ $Y2=0
cc_835 N_VPWR_c_1277_n N_A_737_347#_c_1427_n 0.0135428f $X=4.37 $Y=2.59 $X2=0
+ $Y2=0
cc_836 N_VPWR_c_1287_n N_A_737_347#_c_1427_n 0.00750989f $X=6.795 $Y=3.33 $X2=0
+ $Y2=0
cc_837 N_VPWR_c_1274_n N_A_737_347#_c_1427_n 0.00907713f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_838 N_VPWR_c_1276_n N_A_737_347#_c_1428_n 0.0195142f $X=3.335 $Y=2.17 $X2=0
+ $Y2=0
cc_839 N_VPWR_c_1277_n N_A_737_347#_c_1428_n 0.0131962f $X=4.37 $Y=2.59 $X2=0
+ $Y2=0
cc_840 N_VPWR_c_1286_n N_A_737_347#_c_1428_n 0.00747692f $X=4.17 $Y=3.33 $X2=0
+ $Y2=0
cc_841 N_VPWR_c_1274_n N_A_737_347#_c_1428_n 0.009061f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_842 N_VPWR_c_1278_n N_SUM_c_1467_n 0.0462948f $X=6.96 $Y=2.455 $X2=0 $Y2=0
cc_843 N_VPWR_c_1279_n N_SUM_c_1467_n 0.0536704f $X=7.86 $Y=2.345 $X2=0 $Y2=0
cc_844 N_VPWR_c_1288_n N_SUM_c_1467_n 0.014552f $X=7.775 $Y=3.33 $X2=0 $Y2=0
cc_845 N_VPWR_c_1274_n N_SUM_c_1467_n 0.0119791f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_846 N_VPWR_M1007_s N_SUM_c_1494_n 0.00473157f $X=7.71 $Y=1.84 $X2=0 $Y2=0
cc_847 N_VPWR_c_1279_n N_SUM_c_1494_n 0.0184684f $X=7.86 $Y=2.345 $X2=0 $Y2=0
cc_848 N_VPWR_c_1280_n N_SUM_c_1465_n 0.00130778f $X=8.81 $Y=1.985 $X2=0 $Y2=0
cc_849 N_VPWR_c_1280_n SUM 0.0121024f $X=8.81 $Y=1.985 $X2=0 $Y2=0
cc_850 N_VPWR_c_1279_n SUM 0.0307758f $X=7.86 $Y=2.345 $X2=0 $Y2=0
cc_851 N_VPWR_c_1280_n SUM 0.0650362f $X=8.81 $Y=1.985 $X2=0 $Y2=0
cc_852 N_VPWR_c_1289_n SUM 0.014552f $X=8.725 $Y=3.33 $X2=0 $Y2=0
cc_853 N_VPWR_c_1274_n SUM 0.0119791f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_854 N_VPWR_c_1280_n N_COUT_c_1530_n 0.00792223f $X=8.81 $Y=1.985 $X2=0 $Y2=0
cc_855 N_VPWR_c_1280_n N_COUT_c_1531_n 0.0378676f $X=8.81 $Y=1.985 $X2=0 $Y2=0
cc_856 N_VPWR_c_1281_n N_COUT_c_1531_n 0.0550114f $X=9.76 $Y=2.325 $X2=0 $Y2=0
cc_857 N_VPWR_c_1290_n N_COUT_c_1531_n 0.014552f $X=9.675 $Y=3.33 $X2=0 $Y2=0
cc_858 N_VPWR_c_1274_n N_COUT_c_1531_n 0.0119791f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_859 N_VPWR_M1009_d N_COUT_c_1532_n 0.00275645f $X=9.61 $Y=1.84 $X2=0 $Y2=0
cc_860 N_VPWR_c_1281_n N_COUT_c_1532_n 0.0184684f $X=9.76 $Y=2.325 $X2=0 $Y2=0
cc_861 N_VPWR_c_1283_n N_COUT_c_1533_n 0.012622f $X=10.71 $Y=1.985 $X2=0 $Y2=0
cc_862 N_VPWR_c_1281_n COUT 0.0316672f $X=9.76 $Y=2.325 $X2=0 $Y2=0
cc_863 N_VPWR_c_1283_n COUT 0.0692f $X=10.71 $Y=1.985 $X2=0 $Y2=0
cc_864 N_VPWR_c_1291_n COUT 0.0149683f $X=10.625 $Y=3.33 $X2=0 $Y2=0
cc_865 N_VPWR_c_1274_n COUT 0.0123002f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_866 N_VPWR_c_1283_n N_VGND_c_1630_n 0.00906267f $X=10.71 $Y=1.985 $X2=0 $Y2=0
cc_867 N_SUM_c_1463_n N_VGND_M1021_d 0.00452945f $X=8.285 $Y=1.045 $X2=0 $Y2=0
cc_868 N_COUT_c_1548_n N_VGND_M1014_s 0.00356752f $X=10.165 $Y=1.065 $X2=0 $Y2=0
cc_869 N_COUT_c_1526_n N_VGND_c_1628_n 0.0151543f $X=9.47 $Y=0.555 $X2=0 $Y2=0
cc_870 N_COUT_c_1548_n N_VGND_c_1628_n 0.0152916f $X=10.165 $Y=1.065 $X2=0 $Y2=0
cc_871 N_COUT_c_1528_n N_VGND_c_1628_n 0.0152413f $X=10.33 $Y=0.555 $X2=0 $Y2=0
cc_872 N_COUT_c_1528_n N_VGND_c_1630_n 0.0229007f $X=10.33 $Y=0.555 $X2=0 $Y2=0
cc_873 N_COUT_c_1529_n N_VGND_c_1630_n 0.00151292f $X=10.295 $Y=1.55 $X2=0 $Y2=0
cc_874 N_COUT_c_1526_n N_VGND_c_1638_n 0.00946322f $X=9.47 $Y=0.555 $X2=0 $Y2=0
cc_875 N_COUT_c_1528_n N_VGND_c_1639_n 0.00984752f $X=10.33 $Y=0.555 $X2=0 $Y2=0
cc_876 N_COUT_c_1526_n N_VGND_c_1644_n 0.00148615f $X=9.47 $Y=0.555 $X2=0 $Y2=0
cc_877 N_COUT_c_1526_n N_VGND_c_1646_n 0.00891381f $X=9.47 $Y=0.555 $X2=0 $Y2=0
cc_878 N_COUT_c_1528_n N_VGND_c_1646_n 0.0092741f $X=10.33 $Y=0.555 $X2=0 $Y2=0
cc_879 N_A_27_74#_c_1599_n N_VGND_M1032_d 0.0262462f $X=1.325 $Y=0.55 $X2=-0.19
+ $Y2=-0.245
cc_880 N_A_27_74#_c_1597_n N_VGND_M1032_d 0.00943635f $X=1.495 $Y=0.55 $X2=-0.19
+ $Y2=-0.245
cc_881 N_A_27_74#_c_1599_n N_VGND_c_1631_n 0.003347f $X=1.325 $Y=0.55 $X2=0
+ $Y2=0
cc_882 N_A_27_74#_c_1597_n N_VGND_c_1631_n 0.0265731f $X=1.495 $Y=0.55 $X2=0
+ $Y2=0
cc_883 N_A_27_74#_c_1596_n N_VGND_c_1640_n 0.0145639f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_884 N_A_27_74#_c_1599_n N_VGND_c_1640_n 0.00294077f $X=1.325 $Y=0.55 $X2=0
+ $Y2=0
cc_885 N_A_27_74#_c_1596_n N_VGND_c_1641_n 0.00294333f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_886 N_A_27_74#_c_1599_n N_VGND_c_1641_n 0.0392999f $X=1.325 $Y=0.55 $X2=0
+ $Y2=0
cc_887 N_A_27_74#_c_1597_n N_VGND_c_1641_n 0.00517613f $X=1.495 $Y=0.55 $X2=0
+ $Y2=0
cc_888 N_A_27_74#_c_1596_n N_VGND_c_1646_n 0.0119984f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_889 N_A_27_74#_c_1599_n N_VGND_c_1646_n 0.0124477f $X=1.325 $Y=0.55 $X2=0
+ $Y2=0
cc_890 N_A_27_74#_c_1597_n N_VGND_c_1646_n 0.022248f $X=1.495 $Y=0.55 $X2=0
+ $Y2=0
cc_891 N_VGND_M1030_d N_A_734_74#_c_1776_n 0.0072679f $X=4.1 $Y=0.37 $X2=0 $Y2=0
cc_892 N_VGND_c_1633_n N_A_734_74#_c_1776_n 0.0243979f $X=4.32 $Y=0 $X2=0 $Y2=0
cc_893 N_VGND_c_1634_n N_A_734_74#_c_1776_n 0.0029521f $X=4.155 $Y=0 $X2=0 $Y2=0
cc_894 N_VGND_c_1635_n N_A_734_74#_c_1776_n 0.0029521f $X=6.755 $Y=0 $X2=0 $Y2=0
cc_895 N_VGND_c_1646_n N_A_734_74#_c_1776_n 0.011204f $X=10.8 $Y=0 $X2=0 $Y2=0
cc_896 N_VGND_c_1627_n N_A_734_74#_c_1774_n 0.00129215f $X=3.34 $Y=0.55 $X2=0
+ $Y2=0
cc_897 N_VGND_c_1633_n N_A_734_74#_c_1774_n 0.00282013f $X=4.32 $Y=0 $X2=0 $Y2=0
cc_898 N_VGND_c_1634_n N_A_734_74#_c_1774_n 0.0105866f $X=4.155 $Y=0 $X2=0 $Y2=0
cc_899 N_VGND_c_1646_n N_A_734_74#_c_1774_n 0.00888607f $X=10.8 $Y=0 $X2=0 $Y2=0
cc_900 N_VGND_c_1633_n N_A_734_74#_c_1775_n 0.00282013f $X=4.32 $Y=0 $X2=0 $Y2=0
cc_901 N_VGND_c_1635_n N_A_734_74#_c_1775_n 0.0105866f $X=6.755 $Y=0 $X2=0 $Y2=0
cc_902 N_VGND_c_1646_n N_A_734_74#_c_1775_n 0.00888607f $X=10.8 $Y=0 $X2=0 $Y2=0
