# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__xor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__xor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.804000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 1.165000 0.915000 1.620000 ;
        RECT 0.585000 1.620000 2.515000 1.790000 ;
        RECT 1.845000 1.350000 2.515000 1.620000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.804000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.155000 1.010000 4.145000 1.180000 ;
        RECT 1.155000 1.180000 1.485000 1.450000 ;
        RECT 3.485000 1.180000 4.145000 1.550000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.754100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.025000 1.850000 4.685000 2.020000 ;
        RECT 3.025000 2.020000 3.195000 2.735000 ;
        RECT 3.330000 0.595000 3.660000 0.670000 ;
        RECT 3.330000 0.670000 4.685000 0.840000 ;
        RECT 4.355000 0.350000 4.685000 0.670000 ;
        RECT 4.355000 0.840000 4.685000 1.850000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.085000 0.710000 0.500000 ;
      RECT 0.115000  2.300000 0.445000 3.245000 ;
      RECT 0.245000  0.670000 1.220000 0.840000 ;
      RECT 0.245000  0.840000 0.415000 1.960000 ;
      RECT 0.245000  1.960000 2.855000 2.130000 ;
      RECT 0.890000  0.350000 1.220000 0.670000 ;
      RECT 1.065000  2.130000 1.315000 2.980000 ;
      RECT 1.390000  0.085000 1.720000 0.840000 ;
      RECT 1.545000  2.300000 2.825000 2.470000 ;
      RECT 1.545000  2.470000 1.795000 2.980000 ;
      RECT 1.970000  0.350000 2.300000 0.670000 ;
      RECT 1.970000  0.670000 3.160000 0.840000 ;
      RECT 1.995000  2.640000 2.325000 3.245000 ;
      RECT 2.480000  0.085000 2.820000 0.500000 ;
      RECT 2.495000  2.470000 2.825000 2.905000 ;
      RECT 2.495000  2.905000 3.675000 3.075000 ;
      RECT 2.685000  1.350000 3.125000 1.680000 ;
      RECT 2.685000  1.680000 2.855000 1.960000 ;
      RECT 2.990000  0.255000 4.175000 0.425000 ;
      RECT 2.990000  0.425000 3.160000 0.670000 ;
      RECT 3.395000  2.190000 4.685000 2.360000 ;
      RECT 3.395000  2.360000 3.675000 2.905000 ;
      RECT 3.840000  0.425000 4.175000 0.500000 ;
      RECT 3.845000  2.530000 4.175000 3.245000 ;
      RECT 4.345000  2.360000 4.685000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_ls__xor2_2
END LIBRARY
