* File: sky130_fd_sc_ls__xnor2_4.spice
* Created: Wed Sep  2 11:30:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__xnor2_4.pex.spice"
.subckt sky130_fd_sc_ls__xnor2_4  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1012 N_A_27_74#_M1012_d N_A_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1824 AS=0.112 PD=1.85 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1027 N_A_27_74#_M1027_d N_A_M1027_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75000.7
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1018 N_A_27_74#_M1027_d N_B_M1018_g N_A_116_368#_M1018_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75001.1 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1022 N_A_27_74#_M1022_d N_B_M1022_g N_A_116_368#_M1018_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1824 AS=0.112 PD=1.85 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_A_511_74#_M1005_d N_A_116_368#_M1005_g N_Y_M1005_s VNB NSHORT L=0.15
+ W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.2 SB=75005.9 A=0.111 P=1.78 MULT=1
MM1008 N_A_511_74#_M1008_d N_A_116_368#_M1008_g N_Y_M1005_s VNB NSHORT L=0.15
+ W=0.74 AD=0.16465 AS=0.1295 PD=1.185 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75005.4 A=0.111 P=1.78 MULT=1
MM1011 N_A_511_74#_M1008_d N_A_116_368#_M1011_g N_Y_M1011_s VNB NSHORT L=0.15
+ W=0.74 AD=0.16465 AS=0.1036 PD=1.185 PS=1.02 NRD=15.396 NRS=0 M=1 R=4.93333
+ SA=75001.3 SB=75004.8 A=0.111 P=1.78 MULT=1
MM1028 N_A_511_74#_M1028_d N_A_116_368#_M1028_g N_Y_M1011_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001.7 SB=75004.4 A=0.111 P=1.78 MULT=1
MM1002 N_A_511_74#_M1028_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1889 PD=1.09 PS=1.36 NRD=0 NRS=32.472 M=1 R=4.93333 SA=75002.2
+ SB=75003.9 A=0.111 P=1.78 MULT=1
MM1006 N_A_511_74#_M1006_d N_A_M1006_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1889 PD=1.02 PS=1.36 NRD=0 NRS=32.472 M=1 R=4.93333 SA=75002.8
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1017 N_A_511_74#_M1006_d N_A_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1889 PD=1.02 PS=1.36 NRD=0 NRS=32.472 M=1 R=4.93333 SA=75003.3
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1019 N_A_511_74#_M1019_d N_A_M1019_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1889 PD=1.02 PS=1.36 NRD=0 NRS=32.472 M=1 R=4.93333 SA=75003.8
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1009 N_A_511_74#_M1019_d N_B_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.205 PD=1.02 PS=1.395 NRD=0 NRS=36 M=1 R=4.93333 SA=75004.3
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1010 N_A_511_74#_M1010_d N_B_M1010_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.205 PD=1.02 PS=1.395 NRD=0 NRS=36 M=1 R=4.93333 SA=75004.9
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1020 N_A_511_74#_M1010_d N_B_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1889 PD=1.02 PS=1.36 NRD=0 NRS=32.472 M=1 R=4.93333 SA=75005.3
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1029 N_A_511_74#_M1029_d N_B_M1029_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1889 PD=2.05 PS=1.36 NRD=0 NRS=32.472 M=1 R=4.93333 SA=75005.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_A_116_368#_M1015_d N_A_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.2478 PD=1.14 PS=2.27 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75002.7 A=0.126 P=1.98 MULT=1
MM1016 N_A_116_368#_M1015_d N_A_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.126 PD=1.14 PS=1.14 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75000.7
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1016_s N_B_M1003_g N_A_116_368#_M1003_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.126 AS=0.126 PD=1.14 PS=1.14 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75001.1
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1026 N_VPWR_M1026_d N_B_M1026_g N_A_116_368#_M1003_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.249814 AS=0.126 PD=1.57286 PS=1.14 NRD=56.8345 NRS=2.3443 M=1 R=5.6
+ SA=75001.6 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1014 N_Y_M1014_d N_A_116_368#_M1014_g N_VPWR_M1026_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.333086 PD=1.42 PS=2.09714 NRD=1.7533 NRS=42.6308 M=1 R=7.46667
+ SA=75001.7 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1024 N_Y_M1014_d N_A_116_368#_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.49375 PD=1.42 PS=3.47 NRD=1.7533 NRS=67.8665 M=1 R=7.46667
+ SA=75002.2 SB=75000.3 A=0.168 P=2.54 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_950_368#_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.300662 AS=0.3304 PD=1.83 PS=2.83 NRD=37.5285 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.7 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1000_d N_A_M1004_g N_A_950_368#_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.300662 AS=0.168 PD=1.83 PS=1.42 NRD=37.5285 NRS=1.7533 M=1 R=7.46667
+ SA=75000.8 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1023 N_VPWR_M1023_d N_A_M1023_g N_A_950_368#_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.297275 AS=0.168 PD=1.825 PS=1.42 NRD=36.9966 NRS=1.7533 M=1 R=7.46667
+ SA=75001.3 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1025 N_VPWR_M1023_d N_A_M1025_g N_A_950_368#_M1025_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.297275 AS=0.168 PD=1.825 PS=1.42 NRD=36.9966 NRS=1.7533 M=1 R=7.46667
+ SA=75001.9 SB=75002 A=0.168 P=2.54 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g N_A_950_368#_M1025_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.4 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1001_d N_B_M1007_g N_A_950_368#_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.8 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1013 N_Y_M1013_d N_B_M1013_g N_A_950_368#_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.3 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1021 N_Y_M1013_d N_B_M1021_g N_A_950_368#_M1021_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX30_noxref VNB VPB NWDIODE A=17.67 P=22.72
c_77 VNB 0 1.57454e-19 $X=0 $Y=0
c_143 VPB 0 3.00577e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__xnor2_4.pxi.spice"
*
.ends
*
*
