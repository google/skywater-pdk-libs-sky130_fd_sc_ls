* NGSPICE file created from sky130_fd_sc_ls__decaphe_18.ext - technology: sky130A

.subckt sky130_fd_sc_ls__decaphe_18 VGND VNB VPB VPWR
M1000 VGND VPWR VGND VNB nshort w=775000u l=7.85e+06u
+  ad=4.03e+11p pd=4.14e+06u as=0p ps=0u
M1001 VPWR VGND VPWR VPB pshort w=1.255e+06u l=7.85e+06u
+  ad=6.526e+11p pd=6.06e+06u as=0p ps=0u
.ends

