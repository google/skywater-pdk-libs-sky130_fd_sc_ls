* File: sky130_fd_sc_ls__xnor3_1.spice
* Created: Fri Aug 28 14:09:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__xnor3_1.pex.spice"
.subckt sky130_fd_sc_ls__xnor3_1  VNB VPB C B A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_81_268#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.74
+ AD=0.24975 AS=0.2109 PD=1.90103 PS=2.05 NRD=45.804 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1014 N_A_232_162#_M1014_d N_C_M1014_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1575 AS=0.14175 PD=1.59 PS=1.07897 NRD=0 NRS=80.712 M=1 R=2.8 SA=75000.8
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1011 N_A_81_268#_M1011_d N_C_M1011_g N_A_371_74#_M1011_s VNB NSHORT L=0.15
+ W=0.64 AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1008 N_A_363_394#_M1008_d N_A_232_162#_M1008_g N_A_81_268#_M1011_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.2272 AS=0.112 PD=1.99 PS=0.99 NRD=6.552 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1021 N_A_786_100#_M1021_d N_B_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.36 PD=2.05 PS=2.83 NRD=0 NRS=69.96 M=1 R=4.93333 SA=75000.3
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_A_371_74#_M1010_d N_A_786_100#_M1010_g N_A_897_54#_M1010_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.1328 AS=0.374625 PD=1.055 PS=2.77 NRD=12.18 NRS=99.432 M=1
+ R=4.26667 SA=75000.3 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1001 N_A_1113_383#_M1001_d N_B_M1001_g N_A_371_74#_M1010_d VNB NSHORT L=0.15
+ W=0.64 AD=0.137177 AS=0.1328 PD=1.26792 PS=1.055 NRD=20.616 NRS=13.116 M=1
+ R=4.26667 SA=75000.9 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1020 N_A_363_394#_M1020_d N_A_786_100#_M1020_g N_A_1113_383#_M1001_d VNB
+ NSHORT L=0.15 W=0.42 AD=0.0792057 AS=0.0900226 PD=0.780566 PS=0.832075
+ NRD=18.564 NRS=5.712 M=1 R=2.8 SA=75001.5 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1015 N_A_897_54#_M1015_d N_B_M1015_g N_A_363_394#_M1020_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1104 AS=0.120694 PD=0.985 PS=1.18943 NRD=12.18 NRS=0 M=1 R=4.26667
+ SA=75001.3 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1017 N_VGND_M1017_d N_A_M1017_g N_A_897_54#_M1015_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1376 AS=0.1104 PD=1.07 PS=0.985 NRD=20.616 NRS=0 M=1 R=4.26667 SA=75001.8
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1006 N_A_1113_383#_M1006_d N_A_897_54#_M1006_g N_VGND_M1017_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.1376 PD=1.85 PS=1.07 NRD=0 NRS=7.488 M=1
+ R=4.26667 SA=75002.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 N_VPWR_M1018_d N_A_81_268#_M1018_g N_X_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.305964 AS=0.3192 PD=2.1 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1013 N_A_232_162#_M1013_d N_C_M1013_g N_VPWR_M1018_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1888 AS=0.174836 PD=1.87 PS=1.2 NRD=3.0732 NRS=75.4116 M=1 R=4.26667
+ SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_A_81_268#_M1007_d N_C_M1007_g N_A_363_394#_M1007_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.208975 AS=0.2478 PD=1.425 PS=2.27 NRD=22.261 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1009 N_A_371_74#_M1009_d N_A_232_162#_M1009_g N_A_81_268#_M1007_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2436 AS=0.208975 PD=2.26 PS=1.425 NRD=2.3443 NRS=21.0987
+ M=1 R=5.6 SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1019 N_A_786_100#_M1019_d N_B_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3192 AS=0.4194 PD=2.81 PS=3.08 NRD=1.7533 NRS=15.8191 M=1 R=7.46667
+ SA=75000.3 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1002 N_A_363_394#_M1002_d N_A_786_100#_M1002_g N_A_897_54#_M1002_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.173335 AS=0.36585 PD=1.39054 PS=2.87 NRD=2.3443 NRS=89.241
+ M=1 R=5.6 SA=75000.3 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1003 N_A_1113_383#_M1003_d N_B_M1003_g N_A_363_394#_M1002_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.096 AS=0.132065 PD=0.94 PS=1.05946 NRD=3.0732 NRS=29.2348 M=1
+ R=4.26667 SA=75000.8 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1012 N_A_371_74#_M1012_d N_A_786_100#_M1012_g N_A_1113_383#_M1003_d VPB
+ PHIGHVT L=0.15 W=0.64 AD=0.160173 AS=0.096 PD=1.14595 PS=0.94 NRD=3.0732
+ NRS=3.0732 M=1 R=4.26667 SA=75001.3 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1005 N_A_897_54#_M1005_d N_B_M1005_g N_A_371_74#_M1012_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.169643 AS=0.210227 PD=1.26913 PS=1.50405 NRD=22.261 NRS=45.7237
+ M=1 R=5.6 SA=75001.5 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1016 N_VPWR_M1016_d N_A_M1016_g N_A_897_54#_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1925 AS=0.201957 PD=1.385 PS=1.51087 NRD=18.715 NRS=2.9353 M=1 R=6.66667
+ SA=75001.7 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1004 N_A_1113_383#_M1004_d N_A_897_54#_M1004_g N_VPWR_M1016_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.3 AS=0.1925 PD=2.6 PS=1.385 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75002.3 SB=75000.2 A=0.15 P=2.3 MULT=1
DX22_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ls__xnor3_1.pxi.spice"
*
.ends
*
*
