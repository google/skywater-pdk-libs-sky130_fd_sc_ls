* File: sky130_fd_sc_ls__sdfrtp_2.pxi.spice
* Created: Wed Sep  2 11:27:23 2020
* 
x_PM_SKY130_FD_SC_LS__SDFRTP_2%A_27_74# N_A_27_74#_M1031_s N_A_27_74#_M1022_s
+ N_A_27_74#_c_283_n N_A_27_74#_c_284_n N_A_27_74#_M1005_g N_A_27_74#_c_290_n
+ N_A_27_74#_M1017_g N_A_27_74#_c_285_n N_A_27_74#_c_286_n N_A_27_74#_c_292_n
+ N_A_27_74#_c_287_n N_A_27_74#_c_293_n N_A_27_74#_c_288_n N_A_27_74#_c_294_n
+ N_A_27_74#_c_295_n N_A_27_74#_c_289_n PM_SKY130_FD_SC_LS__SDFRTP_2%A_27_74#
x_PM_SKY130_FD_SC_LS__SDFRTP_2%SCE N_SCE_c_371_n N_SCE_M1031_g N_SCE_c_372_n
+ N_SCE_M1022_g N_SCE_c_373_n N_SCE_c_374_n N_SCE_M1025_g N_SCE_M1026_g
+ N_SCE_c_364_n N_SCE_c_365_n N_SCE_c_366_n N_SCE_c_367_n N_SCE_c_368_n
+ N_SCE_c_369_n SCE SCE SCE N_SCE_c_370_n PM_SKY130_FD_SC_LS__SDFRTP_2%SCE
x_PM_SKY130_FD_SC_LS__SDFRTP_2%D N_D_M1006_g N_D_c_442_n N_D_M1004_g N_D_c_447_n
+ D N_D_c_444_n N_D_c_445_n PM_SKY130_FD_SC_LS__SDFRTP_2%D
x_PM_SKY130_FD_SC_LS__SDFRTP_2%SCD N_SCD_M1027_g N_SCD_M1011_g N_SCD_c_487_n
+ N_SCD_c_491_n SCD SCD N_SCD_c_489_n SCD PM_SKY130_FD_SC_LS__SDFRTP_2%SCD
x_PM_SKY130_FD_SC_LS__SDFRTP_2%CLK N_CLK_c_529_n N_CLK_c_530_n N_CLK_c_531_n
+ N_CLK_M1029_g N_CLK_c_532_n N_CLK_M1028_g N_CLK_c_533_n N_CLK_c_537_n CLK
+ N_CLK_c_535_n PM_SKY130_FD_SC_LS__SDFRTP_2%CLK
x_PM_SKY130_FD_SC_LS__SDFRTP_2%A_1034_392# N_A_1034_392#_M1032_d
+ N_A_1034_392#_M1030_d N_A_1034_392#_c_603_n N_A_1034_392#_c_604_n
+ N_A_1034_392#_M1040_g N_A_1034_392#_c_583_n N_A_1034_392#_M1000_g
+ N_A_1034_392#_c_585_n N_A_1034_392#_M1016_g N_A_1034_392#_c_586_n
+ N_A_1034_392#_c_587_n N_A_1034_392#_c_606_n N_A_1034_392#_M1037_g
+ N_A_1034_392#_c_607_n N_A_1034_392#_c_588_n N_A_1034_392#_c_589_n
+ N_A_1034_392#_c_590_n N_A_1034_392#_c_591_n N_A_1034_392#_c_608_n
+ N_A_1034_392#_c_592_n N_A_1034_392#_c_593_n N_A_1034_392#_c_594_n
+ N_A_1034_392#_c_618_p N_A_1034_392#_c_641_p N_A_1034_392#_c_595_n
+ N_A_1034_392#_c_596_n N_A_1034_392#_c_656_p N_A_1034_392#_c_597_n
+ N_A_1034_392#_c_598_n N_A_1034_392#_c_599_n N_A_1034_392#_c_600_n
+ N_A_1034_392#_c_601_n N_A_1034_392#_c_602_n
+ PM_SKY130_FD_SC_LS__SDFRTP_2%A_1034_392#
x_PM_SKY130_FD_SC_LS__SDFRTP_2%A_1367_93# N_A_1367_93#_M1035_d
+ N_A_1367_93#_M1015_d N_A_1367_93#_M1019_g N_A_1367_93#_M1033_g
+ N_A_1367_93#_c_791_n N_A_1367_93#_c_792_n N_A_1367_93#_c_793_n
+ N_A_1367_93#_c_799_n N_A_1367_93#_c_794_n N_A_1367_93#_c_816_n
+ N_A_1367_93#_c_800_n N_A_1367_93#_c_795_n
+ PM_SKY130_FD_SC_LS__SDFRTP_2%A_1367_93#
x_PM_SKY130_FD_SC_LS__SDFRTP_2%RESET_B N_RESET_B_M1036_g N_RESET_B_M1039_g
+ N_RESET_B_c_891_n N_RESET_B_c_892_n N_RESET_B_c_898_n N_RESET_B_c_899_n
+ N_RESET_B_M1009_g N_RESET_B_c_900_n N_RESET_B_M1001_g N_RESET_B_c_894_n
+ N_RESET_B_M1014_g N_RESET_B_c_903_n N_RESET_B_c_904_n N_RESET_B_M1013_g
+ N_RESET_B_c_905_n N_RESET_B_c_896_n N_RESET_B_c_906_n N_RESET_B_c_907_n
+ N_RESET_B_c_908_n N_RESET_B_c_966_n N_RESET_B_c_909_n RESET_B
+ N_RESET_B_c_910_n N_RESET_B_c_911_n N_RESET_B_c_912_n N_RESET_B_c_1027_p
+ PM_SKY130_FD_SC_LS__SDFRTP_2%RESET_B
x_PM_SKY130_FD_SC_LS__SDFRTP_2%A_1234_119# N_A_1234_119#_M1034_d
+ N_A_1234_119#_M1040_d N_A_1234_119#_M1001_d N_A_1234_119#_M1035_g
+ N_A_1234_119#_c_1111_n N_A_1234_119#_M1015_g N_A_1234_119#_c_1112_n
+ N_A_1234_119#_c_1121_n N_A_1234_119#_c_1113_n N_A_1234_119#_c_1114_n
+ N_A_1234_119#_c_1123_n N_A_1234_119#_c_1124_n N_A_1234_119#_c_1115_n
+ N_A_1234_119#_c_1116_n N_A_1234_119#_c_1117_n N_A_1234_119#_c_1118_n
+ N_A_1234_119#_c_1126_n N_A_1234_119#_c_1194_n N_A_1234_119#_c_1127_n
+ N_A_1234_119#_c_1128_n PM_SKY130_FD_SC_LS__SDFRTP_2%A_1234_119#
x_PM_SKY130_FD_SC_LS__SDFRTP_2%A_835_98# N_A_835_98#_M1029_s N_A_835_98#_M1028_s
+ N_A_835_98#_c_1247_n N_A_835_98#_M1030_g N_A_835_98#_c_1236_n
+ N_A_835_98#_M1032_g N_A_835_98#_c_1248_n N_A_835_98#_c_1249_n
+ N_A_835_98#_c_1250_n N_A_835_98#_c_1237_n N_A_835_98#_c_1238_n
+ N_A_835_98#_M1034_g N_A_835_98#_M1008_g N_A_835_98#_c_1252_n
+ N_A_835_98#_M1018_g N_A_835_98#_c_1239_n N_A_835_98#_c_1255_n
+ N_A_835_98#_c_1240_n N_A_835_98#_M1002_g N_A_835_98#_c_1256_n
+ N_A_835_98#_c_1257_n N_A_835_98#_c_1242_n N_A_835_98#_c_1243_n
+ N_A_835_98#_c_1244_n N_A_835_98#_c_1245_n N_A_835_98#_c_1246_n
+ PM_SKY130_FD_SC_LS__SDFRTP_2%A_835_98#
x_PM_SKY130_FD_SC_LS__SDFRTP_2%A_2082_446# N_A_2082_446#_M1007_d
+ N_A_2082_446#_M1013_d N_A_2082_446#_c_1425_n N_A_2082_446#_M1038_g
+ N_A_2082_446#_M1003_g N_A_2082_446#_c_1426_n N_A_2082_446#_c_1439_n
+ N_A_2082_446#_c_1417_n N_A_2082_446#_c_1418_n N_A_2082_446#_c_1429_n
+ N_A_2082_446#_c_1486_p N_A_2082_446#_c_1430_n N_A_2082_446#_c_1419_n
+ N_A_2082_446#_c_1420_n N_A_2082_446#_c_1421_n N_A_2082_446#_c_1422_n
+ N_A_2082_446#_c_1423_n N_A_2082_446#_c_1424_n
+ PM_SKY130_FD_SC_LS__SDFRTP_2%A_2082_446#
x_PM_SKY130_FD_SC_LS__SDFRTP_2%A_1824_74# N_A_1824_74#_M1016_d
+ N_A_1824_74#_M1018_d N_A_1824_74#_M1007_g N_A_1824_74#_c_1552_n
+ N_A_1824_74#_c_1553_n N_A_1824_74#_c_1554_n N_A_1824_74#_M1024_g
+ N_A_1824_74#_c_1539_n N_A_1824_74#_c_1540_n N_A_1824_74#_c_1541_n
+ N_A_1824_74#_c_1556_n N_A_1824_74#_M1010_g N_A_1824_74#_c_1542_n
+ N_A_1824_74#_M1021_g N_A_1824_74#_c_1543_n N_A_1824_74#_c_1544_n
+ N_A_1824_74#_c_1563_n N_A_1824_74#_c_1545_n N_A_1824_74#_c_1557_n
+ N_A_1824_74#_c_1558_n N_A_1824_74#_c_1546_n N_A_1824_74#_c_1547_n
+ N_A_1824_74#_c_1548_n N_A_1824_74#_c_1549_n N_A_1824_74#_c_1550_n
+ N_A_1824_74#_c_1551_n PM_SKY130_FD_SC_LS__SDFRTP_2%A_1824_74#
x_PM_SKY130_FD_SC_LS__SDFRTP_2%A_2492_392# N_A_2492_392#_M1021_d
+ N_A_2492_392#_M1010_d N_A_2492_392#_c_1689_n N_A_2492_392#_M1012_g
+ N_A_2492_392#_M1023_g N_A_2492_392#_c_1690_n N_A_2492_392#_M1020_g
+ N_A_2492_392#_M1041_g N_A_2492_392#_c_1691_n N_A_2492_392#_c_1692_n
+ N_A_2492_392#_c_1684_n N_A_2492_392#_c_1685_n N_A_2492_392#_c_1686_n
+ N_A_2492_392#_c_1687_n N_A_2492_392#_c_1688_n
+ PM_SKY130_FD_SC_LS__SDFRTP_2%A_2492_392#
x_PM_SKY130_FD_SC_LS__SDFRTP_2%VPWR N_VPWR_M1022_d N_VPWR_M1027_d N_VPWR_M1028_d
+ N_VPWR_M1033_d N_VPWR_M1015_s N_VPWR_M1038_d N_VPWR_M1024_d N_VPWR_M1012_s
+ N_VPWR_M1020_s N_VPWR_c_1745_n N_VPWR_c_1746_n N_VPWR_c_1747_n N_VPWR_c_1748_n
+ N_VPWR_c_1749_n N_VPWR_c_1750_n N_VPWR_c_1751_n N_VPWR_c_1752_n
+ N_VPWR_c_1753_n N_VPWR_c_1754_n N_VPWR_c_1755_n N_VPWR_c_1756_n
+ N_VPWR_c_1757_n N_VPWR_c_1758_n VPWR N_VPWR_c_1759_n N_VPWR_c_1760_n
+ N_VPWR_c_1761_n N_VPWR_c_1762_n N_VPWR_c_1763_n N_VPWR_c_1764_n
+ N_VPWR_c_1765_n N_VPWR_c_1766_n N_VPWR_c_1767_n N_VPWR_c_1768_n
+ N_VPWR_c_1769_n N_VPWR_c_1744_n PM_SKY130_FD_SC_LS__SDFRTP_2%VPWR
x_PM_SKY130_FD_SC_LS__SDFRTP_2%A_390_81# N_A_390_81#_M1006_d N_A_390_81#_M1034_s
+ N_A_390_81#_M1004_d N_A_390_81#_M1039_d N_A_390_81#_M1040_s
+ N_A_390_81#_c_1916_n N_A_390_81#_c_1932_n N_A_390_81#_c_1917_n
+ N_A_390_81#_c_1924_n N_A_390_81#_c_1925_n N_A_390_81#_c_1926_n
+ N_A_390_81#_c_1918_n N_A_390_81#_c_1919_n N_A_390_81#_c_1927_n
+ N_A_390_81#_c_1920_n N_A_390_81#_c_1921_n N_A_390_81#_c_1928_n
+ N_A_390_81#_c_1929_n N_A_390_81#_c_1922_n N_A_390_81#_c_1931_n
+ PM_SKY130_FD_SC_LS__SDFRTP_2%A_390_81#
x_PM_SKY130_FD_SC_LS__SDFRTP_2%Q N_Q_M1023_s N_Q_M1012_d N_Q_c_2074_n Q Q Q Q
+ PM_SKY130_FD_SC_LS__SDFRTP_2%Q
x_PM_SKY130_FD_SC_LS__SDFRTP_2%VGND N_VGND_M1031_d N_VGND_M1036_d N_VGND_M1029_d
+ N_VGND_M1009_d N_VGND_M1003_d N_VGND_M1021_s N_VGND_M1023_d N_VGND_M1041_d
+ N_VGND_c_2095_n N_VGND_c_2096_n N_VGND_c_2097_n N_VGND_c_2098_n
+ N_VGND_c_2099_n N_VGND_c_2100_n N_VGND_c_2101_n N_VGND_c_2102_n
+ N_VGND_c_2103_n N_VGND_c_2104_n N_VGND_c_2105_n N_VGND_c_2106_n VGND
+ N_VGND_c_2107_n N_VGND_c_2108_n N_VGND_c_2109_n N_VGND_c_2110_n
+ N_VGND_c_2111_n N_VGND_c_2112_n N_VGND_c_2113_n N_VGND_c_2114_n
+ N_VGND_c_2115_n N_VGND_c_2116_n N_VGND_c_2117_n N_VGND_c_2118_n
+ PM_SKY130_FD_SC_LS__SDFRTP_2%VGND
x_PM_SKY130_FD_SC_LS__SDFRTP_2%noxref_24 N_noxref_24_M1005_s N_noxref_24_M1011_d
+ N_noxref_24_c_2234_n N_noxref_24_c_2248_n N_noxref_24_c_2235_n
+ PM_SKY130_FD_SC_LS__SDFRTP_2%noxref_24
cc_1 VNB N_A_27_74#_c_283_n 0.0258189f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_2 VNB N_A_27_74#_c_284_n 0.0202565f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_3 VNB N_A_27_74#_c_285_n 0.0257773f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_4 VNB N_A_27_74#_c_286_n 0.018732f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_5 VNB N_A_27_74#_c_287_n 0.00973186f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_6 VNB N_A_27_74#_c_288_n 0.018224f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_7 VNB N_A_27_74#_c_289_n 0.0395906f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.01
cc_8 VNB N_SCE_M1031_g 0.0669677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_SCE_c_364_n 0.00778437f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_10 VNB N_SCE_c_365_n 0.0421461f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_11 VNB N_SCE_c_366_n 0.0150893f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_12 VNB N_SCE_c_367_n 0.0126529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_SCE_c_368_n 0.0258818f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_14 VNB N_SCE_c_369_n 0.0297017f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_15 VNB N_SCE_c_370_n 0.0121586f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_16 VNB N_D_c_442_n 0.0268599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB D 0.00947517f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_18 VNB N_D_c_444_n 0.0371634f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_19 VNB N_D_c_445_n 0.0161524f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.935
cc_20 VNB N_SCD_M1011_g 0.0386753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_SCD_c_487_n 0.00375249f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_22 VNB SCD 0.00299368f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.245
cc_23 VNB N_SCD_c_489_n 0.015301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_CLK_c_529_n 0.0269111f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_25 VNB N_CLK_c_530_n 0.0128563f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=2.32
cc_26 VNB N_CLK_c_531_n 0.0155002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_CLK_c_532_n 0.00452949f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_28 VNB N_CLK_c_533_n 0.00964253f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.245
cc_29 VNB CLK 0.017894f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_30 VNB N_CLK_c_535_n 0.0381944f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_31 VNB N_A_1034_392#_c_583_n 0.0113969f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.245
cc_32 VNB N_A_1034_392#_M1000_g 0.0378998f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_33 VNB N_A_1034_392#_c_585_n 0.0171555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_1034_392#_c_586_n 0.0222225f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_35 VNB N_A_1034_392#_c_587_n 0.0102361f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_36 VNB N_A_1034_392#_c_588_n 0.00991314f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.09
cc_37 VNB N_A_1034_392#_c_589_n 6.30651e-19 $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_38 VNB N_A_1034_392#_c_590_n 0.0329865f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_39 VNB N_A_1034_392#_c_591_n 0.00321642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1034_392#_c_592_n 0.00171326f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.01
cc_41 VNB N_A_1034_392#_c_593_n 0.00375765f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_42 VNB N_A_1034_392#_c_594_n 8.50976e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1034_392#_c_595_n 0.011598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1034_392#_c_596_n 0.00281818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1034_392#_c_597_n 0.00595338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1034_392#_c_598_n 0.00363165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1034_392#_c_599_n 0.0322548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1034_392#_c_600_n 0.0101868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1034_392#_c_601_n 4.42537e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1034_392#_c_602_n 0.0114218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1367_93#_M1019_g 0.030989f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_52 VNB N_A_1367_93#_c_791_n 0.00389529f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_53 VNB N_A_1367_93#_c_792_n 0.0235983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1367_93#_c_793_n 4.58327e-19 $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_55 VNB N_A_1367_93#_c_794_n 0.00811998f $X=-0.19 $Y=-0.245 $X2=2.375 $Y2=2.09
cc_56 VNB N_A_1367_93#_c_795_n 0.0146516f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_57 VNB N_RESET_B_M1036_g 0.0458723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_RESET_B_c_891_n 0.27239f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.01
cc_59 VNB N_RESET_B_c_892_n 0.012806f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_60 VNB N_RESET_B_M1009_g 0.0265319f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.935
cc_61 VNB N_RESET_B_c_894_n 0.0204626f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_62 VNB N_RESET_B_M1014_g 0.0531601f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_63 VNB N_RESET_B_c_896_n 0.0328935f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_64 VNB N_A_1234_119#_M1035_g 0.0245433f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.245
cc_65 VNB N_A_1234_119#_c_1111_n 0.0172777f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.64
cc_66 VNB N_A_1234_119#_c_1112_n 0.0274717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1234_119#_c_1113_n 0.0028857f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.465
cc_68 VNB N_A_1234_119#_c_1114_n 0.00422204f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.1
cc_69 VNB N_A_1234_119#_c_1115_n 6.72487e-19 $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_70 VNB N_A_1234_119#_c_1116_n 0.00192123f $X=-0.19 $Y=-0.245 $X2=2.5
+ $Y2=1.995
cc_71 VNB N_A_1234_119#_c_1117_n 0.00723053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1234_119#_c_1118_n 0.00301796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_835_98#_c_1236_n 0.0155098f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_74 VNB N_A_835_98#_c_1237_n 0.0316811f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_75 VNB N_A_835_98#_c_1238_n 0.0159407f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_76 VNB N_A_835_98#_c_1239_n 0.012531f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_77 VNB N_A_835_98#_c_1240_n 0.0236403f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_78 VNB N_A_835_98#_M1002_g 0.027022f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=2.09
cc_79 VNB N_A_835_98#_c_1242_n 0.0209137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_835_98#_c_1243_n 0.00128593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_835_98#_c_1244_n 0.00398883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_835_98#_c_1245_n 0.00150962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_835_98#_c_1246_n 0.0545089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_2082_446#_M1003_g 0.0407896f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.245
cc_85 VNB N_A_2082_446#_c_1417_n 0.00604102f $X=-0.19 $Y=-0.245 $X2=0.2
+ $Y2=1.265
cc_86 VNB N_A_2082_446#_c_1418_n 0.00978233f $X=-0.19 $Y=-0.245 $X2=0.2
+ $Y2=2.005
cc_87 VNB N_A_2082_446#_c_1419_n 0.00743589f $X=-0.19 $Y=-0.245 $X2=2.375
+ $Y2=2.09
cc_88 VNB N_A_2082_446#_c_1420_n 0.00688415f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_89 VNB N_A_2082_446#_c_1421_n 0.00281201f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.09
cc_90 VNB N_A_2082_446#_c_1422_n 0.00528256f $X=-0.19 $Y=-0.245 $X2=2.5
+ $Y2=1.995
cc_91 VNB N_A_2082_446#_c_1423_n 0.00129589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2082_446#_c_1424_n 0.0231274f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=2.09
cc_93 VNB N_A_1824_74#_M1007_g 0.0313995f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_94 VNB N_A_1824_74#_c_1539_n 0.0313227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1824_74#_c_1540_n 0.0323107f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_96 VNB N_A_1824_74#_c_1541_n 0.0156535f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_97 VNB N_A_1824_74#_c_1542_n 0.0193338f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_98 VNB N_A_1824_74#_c_1543_n 0.0143534f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_99 VNB N_A_1824_74#_c_1544_n 0.0203145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1824_74#_c_1545_n 0.00728448f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_101 VNB N_A_1824_74#_c_1546_n 0.00580575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1824_74#_c_1547_n 0.00783827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1824_74#_c_1548_n 0.0103967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1824_74#_c_1549_n 4.11765e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1824_74#_c_1550_n 0.0164314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1824_74#_c_1551_n 0.00253069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_2492_392#_M1023_g 0.0229518f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.245
cc_108 VNB N_A_2492_392#_M1041_g 0.0260209f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_109 VNB N_A_2492_392#_c_1684_n 0.0162202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_2492_392#_c_1685_n 0.0113264f $X=-0.19 $Y=-0.245 $X2=2.5
+ $Y2=1.995
cc_111 VNB N_A_2492_392#_c_1686_n 7.87382e-19 $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=2.09
cc_112 VNB N_A_2492_392#_c_1687_n 0.00922601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2492_392#_c_1688_n 0.0953071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VPWR_c_1744_n 0.601534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_390_81#_c_1916_n 0.0297923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_390_81#_c_1917_n 0.00321538f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_117 VNB N_A_390_81#_c_1918_n 9.90482e-19 $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_118 VNB N_A_390_81#_c_1919_n 0.00159941f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_119 VNB N_A_390_81#_c_1920_n 0.00510468f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=2.09
cc_120 VNB N_A_390_81#_c_1921_n 0.00161453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_390_81#_c_1922_n 0.0025068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_Q_c_2074_n 2.86109e-19 $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_123 VNB Q 0.00240191f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_124 VNB N_VGND_c_2095_n 0.0110567f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_125 VNB N_VGND_c_2096_n 0.00699239f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=2.09
cc_126 VNB N_VGND_c_2097_n 0.0125052f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_127 VNB N_VGND_c_2098_n 0.0067048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2099_n 0.00861345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2100_n 0.0169646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2101_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2102_n 0.0505973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2103_n 0.0640331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2104_n 0.00359556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2105_n 0.0217694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2106_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2107_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2108_n 0.0552549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2109_n 0.0756669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2110_n 0.0296745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2111_n 0.0187654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2112_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2113_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2114_n 0.0146197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2115_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2116_n 0.00613227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2117_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2118_n 0.749906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_noxref_24_c_2234_n 0.0156963f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_149 VNB N_noxref_24_c_2235_n 0.00655627f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.64
cc_150 VPB N_A_27_74#_c_290_n 0.0503982f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.245
cc_151 VPB N_A_27_74#_c_286_n 0.0161943f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_152 VPB N_A_27_74#_c_292_n 0.0338402f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_153 VPB N_A_27_74#_c_293_n 0.0338778f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_154 VPB N_A_27_74#_c_294_n 0.0129728f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_155 VPB N_A_27_74#_c_295_n 0.00577366f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_156 VPB N_SCE_c_371_n 0.0264922f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=2.32
cc_157 VPB N_SCE_c_372_n 0.0318721f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.01
cc_158 VPB N_SCE_c_373_n 0.0231924f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_159 VPB N_SCE_c_374_n 0.0275748f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.245
cc_160 VPB N_SCE_c_364_n 0.00782879f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_161 VPB N_SCE_c_365_n 0.0410982f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_162 VPB N_SCE_c_368_n 0.0100126f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_163 VPB N_D_c_442_n 0.0251089f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_D_c_447_n 0.0214007f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_165 VPB N_SCD_c_487_n 0.0284918f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_166 VPB N_SCD_c_491_n 0.032062f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_167 VPB SCD 0.00204244f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.245
cc_168 VPB SCD 0.00309096f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_169 VPB N_CLK_c_532_n 0.00946373f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.01
cc_170 VPB N_CLK_c_537_n 0.0260159f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_171 VPB N_A_1034_392#_c_603_n 0.0152883f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.01
cc_172 VPB N_A_1034_392#_c_604_n 0.0194827f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_173 VPB N_A_1034_392#_c_583_n 0.012785f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.245
cc_174 VPB N_A_1034_392#_c_606_n 0.0670682f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_175 VPB N_A_1034_392#_c_607_n 0.00243629f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_176 VPB N_A_1034_392#_c_608_n 0.00144418f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_177 VPB N_A_1034_392#_c_592_n 0.0019321f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.01
cc_178 VPB N_A_1034_392#_c_600_n 0.00643236f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_1034_392#_c_602_n 0.0175819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_1367_93#_M1033_g 0.0381305f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_181 VPB N_A_1367_93#_c_791_n 0.00183672f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_182 VPB N_A_1367_93#_c_792_n 0.0212319f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_1367_93#_c_799_n 5.83952e-19 $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_184 VPB N_A_1367_93#_c_800_n 0.00552703f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_185 VPB N_A_1367_93#_c_795_n 0.00452983f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_186 VPB N_RESET_B_M1036_g 0.00778474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_RESET_B_c_898_n 0.0402856f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_188 VPB N_RESET_B_c_899_n 0.0302301f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_189 VPB N_RESET_B_c_900_n 0.017445f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.58
cc_190 VPB N_RESET_B_c_894_n 0.0098094f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_191 VPB N_RESET_B_M1014_g 0.0132171f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_192 VPB N_RESET_B_c_903_n 0.00850302f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_193 VPB N_RESET_B_c_904_n 0.0233033f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_194 VPB N_RESET_B_c_905_n 0.0216256f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.1
cc_195 VPB N_RESET_B_c_906_n 0.0180958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_RESET_B_c_907_n 0.00158906f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_197 VPB N_RESET_B_c_908_n 0.0135889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_RESET_B_c_909_n 0.0206686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_RESET_B_c_910_n 0.00811747f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_RESET_B_c_911_n 0.0706585f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_RESET_B_c_912_n 0.035184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_1234_119#_c_1111_n 0.0299658f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_203 VPB N_A_1234_119#_c_1112_n 0.0106164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_1234_119#_c_1121_n 0.00449915f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_205 VPB N_A_1234_119#_c_1114_n 0.00354403f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_206 VPB N_A_1234_119#_c_1123_n 0.00182206f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_207 VPB N_A_1234_119#_c_1124_n 0.00814204f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_1234_119#_c_1115_n 0.00255881f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.1
cc_209 VPB N_A_1234_119#_c_1126_n 8.22498e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_1234_119#_c_1127_n 0.00316701f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_1234_119#_c_1128_n 0.00257652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_835_98#_c_1247_n 0.0162235f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.01
cc_213 VPB N_A_835_98#_c_1248_n 0.0722913f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_214 VPB N_A_835_98#_c_1249_n 0.0567222f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.935
cc_215 VPB N_A_835_98#_c_1250_n 0.0123764f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.58
cc_216 VPB N_A_835_98#_M1008_g 0.0386451f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_835_98#_c_1252_n 0.196972f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_218 VPB N_A_835_98#_M1018_g 0.010423f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=2.09
cc_219 VPB N_A_835_98#_c_1239_n 0.03645f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.1
cc_220 VPB N_A_835_98#_c_1255_n 0.0129219f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_221 VPB N_A_835_98#_c_1256_n 0.00749069f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.01
cc_222 VPB N_A_835_98#_c_1257_n 0.0289165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_835_98#_c_1245_n 0.00811881f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_835_98#_c_1246_n 0.028132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_2082_446#_c_1425_n 0.0165865f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.01
cc_226 VPB N_A_2082_446#_c_1426_n 0.0276144f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_227 VPB N_A_2082_446#_c_1417_n 0.0447354f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_228 VPB N_A_2082_446#_c_1418_n 0.0137444f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_229 VPB N_A_2082_446#_c_1429_n 0.00779622f $X=-0.19 $Y=1.66 $X2=0.28
+ $Y2=2.465
cc_230 VPB N_A_2082_446#_c_1430_n 0.00256678f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_231 VPB N_A_1824_74#_c_1552_n 0.00554553f $X=-0.19 $Y=1.66 $X2=1.485
+ $Y2=0.615
cc_232 VPB N_A_1824_74#_c_1553_n 0.0382574f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.245
cc_233 VPB N_A_1824_74#_c_1554_n 0.0224017f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_234 VPB N_A_1824_74#_c_1541_n 0.00845967f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_235 VPB N_A_1824_74#_c_1556_n 0.0253471f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_236 VPB N_A_1824_74#_c_1557_n 0.0061417f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_237 VPB N_A_1824_74#_c_1558_n 0.00281397f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_1824_74#_c_1547_n 0.0144635f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_2492_392#_c_1689_n 0.0177177f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.01
cc_240 VPB N_A_2492_392#_c_1690_n 0.0174134f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_241 VPB N_A_2492_392#_c_1691_n 0.00506653f $X=-0.19 $Y=1.66 $X2=0.28
+ $Y2=2.465
cc_242 VPB N_A_2492_392#_c_1692_n 0.0105448f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_243 VPB N_A_2492_392#_c_1686_n 0.00706142f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_244 VPB N_A_2492_392#_c_1688_n 0.0176866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1745_n 0.0066123f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_246 VPB N_VPWR_c_1746_n 0.00396467f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_247 VPB N_VPWR_c_1747_n 0.0157581f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_248 VPB N_VPWR_c_1748_n 0.0233377f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_249 VPB N_VPWR_c_1749_n 0.0194601f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1750_n 0.0187962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1751_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1752_n 0.0688105f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1753_n 0.0348441f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1754_n 0.00601569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1755_n 0.0551755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1756_n 0.00317016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1757_n 0.0198404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1758_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1759_n 0.0191816f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1760_n 0.0457766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1761_n 0.0274158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1762_n 0.0534696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1763_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1764_n 0.0174925f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1765_n 0.0312859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1766_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1767_n 0.00443527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1768_n 0.0232464f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1769_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1744_n 0.117041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_390_81#_c_1917_n 0.00666589f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_272 VPB N_A_390_81#_c_1924_n 8.30015e-19 $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_273 VPB N_A_390_81#_c_1925_n 0.016932f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_274 VPB N_A_390_81#_c_1926_n 0.00361747f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_275 VPB N_A_390_81#_c_1927_n 0.00289353f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_390_81#_c_1928_n 0.00543975f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.01
cc_277 VPB N_A_390_81#_c_1929_n 0.001897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_A_390_81#_c_1922_n 0.00484787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_390_81#_c_1931_n 0.00248457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_Q_c_2074_n 0.00395156f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_281 N_A_27_74#_c_293_n N_SCE_c_371_n 0.00797393f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_282 N_A_27_74#_c_294_n N_SCE_c_371_n 0.00496169f $X=0.28 $Y=2.09 $X2=0 $Y2=0
cc_283 N_A_27_74#_c_285_n N_SCE_M1031_g 0.00686809f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_284 N_A_27_74#_c_286_n N_SCE_M1031_g 0.00827951f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_285 N_A_27_74#_c_287_n N_SCE_M1031_g 0.0245034f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_286 N_A_27_74#_c_289_n N_SCE_M1031_g 0.0181297f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_287 N_A_27_74#_c_292_n N_SCE_c_372_n 0.0173713f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_288 N_A_27_74#_c_293_n N_SCE_c_372_n 0.00721429f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_289 N_A_27_74#_c_294_n N_SCE_c_372_n 4.59028e-19 $X=0.28 $Y=2.09 $X2=0 $Y2=0
cc_290 N_A_27_74#_c_293_n N_SCE_c_373_n 0.0100663f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_291 N_A_27_74#_c_293_n N_SCE_c_374_n 0.00784761f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_292 N_A_27_74#_c_286_n N_SCE_c_364_n 0.0152937f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_293 N_A_27_74#_c_287_n N_SCE_c_364_n 0.00183089f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_294 N_A_27_74#_c_283_n N_SCE_c_365_n 0.0106974f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_295 N_A_27_74#_c_287_n N_SCE_c_365_n 4.10759e-19 $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_296 N_A_27_74#_c_293_n N_SCE_c_365_n 0.0170396f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_297 N_A_27_74#_c_289_n N_SCE_c_365_n 0.0175645f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_298 N_A_27_74#_c_283_n N_SCE_c_368_n 0.00818136f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_290_n N_SCE_c_368_n 0.00153728f $X=2.485 $Y=2.245 $X2=0
+ $Y2=0
cc_300 N_A_27_74#_c_286_n N_SCE_c_368_n 0.0273677f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_301 N_A_27_74#_c_287_n N_SCE_c_368_n 0.0446621f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_302 N_A_27_74#_c_293_n N_SCE_c_368_n 0.139132f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_303 N_A_27_74#_c_295_n N_SCE_c_368_n 0.0272862f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_304 N_A_27_74#_c_289_n N_SCE_c_368_n 0.00202099f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_305 N_A_27_74#_c_290_n N_SCE_c_369_n 0.0175948f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_306 N_A_27_74#_c_295_n N_SCE_c_369_n 3.7877e-19 $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_307 N_A_27_74#_c_290_n N_D_c_442_n 0.0213701f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_308 N_A_27_74#_c_293_n N_D_c_442_n 0.00770606f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_309 N_A_27_74#_c_295_n N_D_c_442_n 0.00113412f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_310 N_A_27_74#_c_290_n N_D_c_447_n 0.0143856f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_311 N_A_27_74#_c_293_n N_D_c_447_n 0.00696286f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_312 N_A_27_74#_c_284_n D 0.00559191f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_313 N_A_27_74#_c_287_n D 0.0143876f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_314 N_A_27_74#_c_289_n D 8.79717e-19 $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_315 N_A_27_74#_c_283_n N_D_c_444_n 0.00979672f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_316 N_A_27_74#_c_287_n N_D_c_444_n 2.46837e-19 $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_317 N_A_27_74#_c_289_n N_D_c_444_n 0.00222688f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_318 N_A_27_74#_c_284_n N_D_c_445_n 0.0338541f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_319 N_A_27_74#_c_290_n N_SCD_c_487_n 0.0198002f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_320 N_A_27_74#_c_295_n N_SCD_c_487_n 0.00169063f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_321 N_A_27_74#_c_290_n N_SCD_c_491_n 0.0292143f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_322 N_A_27_74#_c_295_n SCD 0.0103734f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_323 N_A_27_74#_c_290_n SCD 5.41362e-19 $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_324 N_A_27_74#_c_295_n SCD 0.014782f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_325 N_A_27_74#_c_290_n N_VPWR_c_1745_n 0.00141701f $X=2.485 $Y=2.245 $X2=0
+ $Y2=0
cc_326 N_A_27_74#_c_292_n N_VPWR_c_1759_n 0.0145938f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_327 N_A_27_74#_c_290_n N_VPWR_c_1760_n 0.00445602f $X=2.485 $Y=2.245 $X2=0
+ $Y2=0
cc_328 N_A_27_74#_c_292_n N_VPWR_c_1765_n 0.0247088f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_329 N_A_27_74#_c_293_n N_VPWR_c_1765_n 0.0746993f $X=2.375 $Y=2.09 $X2=0
+ $Y2=0
cc_330 N_A_27_74#_c_290_n N_VPWR_c_1744_n 0.00448766f $X=2.485 $Y=2.245 $X2=0
+ $Y2=0
cc_331 N_A_27_74#_c_292_n N_VPWR_c_1744_n 0.0120466f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_332 N_A_27_74#_c_290_n N_A_390_81#_c_1932_n 0.0100562f $X=2.485 $Y=2.245
+ $X2=0 $Y2=0
cc_333 N_A_27_74#_c_295_n N_A_390_81#_c_1932_n 0.0188695f $X=2.5 $Y=1.995 $X2=0
+ $Y2=0
cc_334 N_A_27_74#_c_290_n N_A_390_81#_c_1931_n 0.0100573f $X=2.485 $Y=2.245
+ $X2=0 $Y2=0
cc_335 N_A_27_74#_c_293_n N_A_390_81#_c_1931_n 0.0192938f $X=2.375 $Y=2.09 $X2=0
+ $Y2=0
cc_336 N_A_27_74#_c_295_n N_A_390_81#_c_1931_n 0.00253584f $X=2.5 $Y=1.995 $X2=0
+ $Y2=0
cc_337 N_A_27_74#_c_284_n N_VGND_c_2095_n 0.00287309f $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_338 N_A_27_74#_c_285_n N_VGND_c_2095_n 0.0156021f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_339 N_A_27_74#_c_287_n N_VGND_c_2095_n 0.0254818f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_340 N_A_27_74#_c_289_n N_VGND_c_2095_n 0.00149092f $X=0.975 $Y=1.01 $X2=0
+ $Y2=0
cc_341 N_A_27_74#_c_284_n N_VGND_c_2103_n 9.09582e-19 $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_342 N_A_27_74#_c_285_n N_VGND_c_2107_n 0.011066f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_343 N_A_27_74#_c_285_n N_VGND_c_2118_n 0.00915947f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_344 N_A_27_74#_c_284_n N_noxref_24_c_2234_n 0.0108727f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_345 N_A_27_74#_c_284_n N_noxref_24_c_2235_n 0.00824832f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_346 N_A_27_74#_c_287_n N_noxref_24_c_2235_n 0.00178881f $X=0.975 $Y=1.1 $X2=0
+ $Y2=0
cc_347 N_A_27_74#_c_289_n N_noxref_24_c_2235_n 0.00859402f $X=0.975 $Y=1.01
+ $X2=0 $Y2=0
cc_348 N_SCE_c_365_n N_D_c_442_n 0.020652f $X=1.535 $Y=1.67 $X2=0 $Y2=0
cc_349 N_SCE_c_368_n N_D_c_442_n 0.0203012f $X=2.033 $Y=1.662 $X2=0 $Y2=0
cc_350 N_SCE_c_373_n N_D_c_447_n 0.020652f $X=1.625 $Y=2.155 $X2=0 $Y2=0
cc_351 N_SCE_c_374_n N_D_c_447_n 0.0372975f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_352 N_SCE_c_365_n D 0.00107772f $X=1.535 $Y=1.67 $X2=0 $Y2=0
cc_353 N_SCE_c_366_n D 0.00153875f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_354 N_SCE_c_367_n D 0.00254389f $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_355 N_SCE_c_368_n D 0.036943f $X=2.033 $Y=1.662 $X2=0 $Y2=0
cc_356 N_SCE_c_367_n N_D_c_444_n 0.0109066f $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_357 N_SCE_c_368_n N_D_c_444_n 0.00271432f $X=2.033 $Y=1.662 $X2=0 $Y2=0
cc_358 N_SCE_c_369_n N_D_c_444_n 0.0203067f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_359 N_SCE_c_366_n N_D_c_445_n 0.00703815f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_360 N_SCE_c_367_n N_D_c_445_n 5.13516e-19 $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_361 N_SCE_c_366_n N_SCD_M1011_g 0.0413189f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_362 N_SCE_c_368_n N_SCD_M1011_g 0.00364537f $X=2.033 $Y=1.662 $X2=0 $Y2=0
cc_363 N_SCE_c_370_n N_SCD_M1011_g 0.0152935f $X=2.51 $Y=1.26 $X2=0 $Y2=0
cc_364 N_SCE_c_368_n N_SCD_c_487_n 0.00446886f $X=2.033 $Y=1.662 $X2=0 $Y2=0
cc_365 N_SCE_c_368_n SCD 0.0141219f $X=2.033 $Y=1.662 $X2=0 $Y2=0
cc_366 N_SCE_c_368_n N_SCD_c_489_n 0.00270439f $X=2.033 $Y=1.662 $X2=0 $Y2=0
cc_367 N_SCE_c_369_n N_SCD_c_489_n 0.00938989f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_368 N_SCE_c_372_n N_VPWR_c_1759_n 0.00445602f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_369 N_SCE_c_374_n N_VPWR_c_1760_n 0.00415318f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_370 N_SCE_c_372_n N_VPWR_c_1765_n 0.017697f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_371 N_SCE_c_374_n N_VPWR_c_1765_n 0.0162868f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_372 N_SCE_c_372_n N_VPWR_c_1744_n 0.00865213f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_373 N_SCE_c_374_n N_VPWR_c_1744_n 0.00817532f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_374 N_SCE_c_366_n N_A_390_81#_c_1916_n 0.0135725f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_375 N_SCE_c_367_n N_A_390_81#_c_1916_n 0.00561864f $X=2.625 $Y=1.05 $X2=0
+ $Y2=0
cc_376 N_SCE_c_368_n N_A_390_81#_c_1916_n 0.0169341f $X=2.033 $Y=1.662 $X2=0
+ $Y2=0
cc_377 N_SCE_c_369_n N_A_390_81#_c_1916_n 0.00156175f $X=2.51 $Y=1.425 $X2=0
+ $Y2=0
cc_378 N_SCE_c_370_n N_A_390_81#_c_1916_n 0.00559641f $X=2.51 $Y=1.26 $X2=0
+ $Y2=0
cc_379 N_SCE_c_374_n N_A_390_81#_c_1931_n 0.0018587f $X=1.625 $Y=2.245 $X2=0
+ $Y2=0
cc_380 N_SCE_M1031_g N_VGND_c_2095_n 0.0129468f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_381 N_SCE_c_366_n N_VGND_c_2103_n 9.15902e-19 $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_382 N_SCE_M1031_g N_VGND_c_2107_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_383 N_SCE_M1031_g N_VGND_c_2118_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_384 N_SCE_c_366_n N_noxref_24_c_2234_n 0.0107418f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_385 N_SCE_M1031_g N_noxref_24_c_2235_n 9.19966e-19 $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_386 N_D_c_447_n N_VPWR_c_1760_n 0.00434272f $X=2.04 $Y=2.245 $X2=0 $Y2=0
cc_387 N_D_c_447_n N_VPWR_c_1765_n 0.00235425f $X=2.04 $Y=2.245 $X2=0 $Y2=0
cc_388 N_D_c_447_n N_VPWR_c_1744_n 0.00821463f $X=2.04 $Y=2.245 $X2=0 $Y2=0
cc_389 D N_A_390_81#_M1006_d 0.00319564f $X=1.595 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_390 D N_A_390_81#_c_1916_n 0.0219281f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_391 N_D_c_445_n N_A_390_81#_c_1916_n 8.49892e-19 $X=1.947 $Y=0.935 $X2=0
+ $Y2=0
cc_392 N_D_c_447_n N_A_390_81#_c_1931_n 0.0118376f $X=2.04 $Y=2.245 $X2=0 $Y2=0
cc_393 N_D_c_445_n N_VGND_c_2103_n 9.15902e-19 $X=1.947 $Y=0.935 $X2=0 $Y2=0
cc_394 D N_noxref_24_c_2234_n 0.0273249f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_395 N_D_c_444_n N_noxref_24_c_2234_n 0.00116484f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_396 N_D_c_445_n N_noxref_24_c_2234_n 0.0107356f $X=1.947 $Y=0.935 $X2=0 $Y2=0
cc_397 N_D_c_445_n N_noxref_24_c_2235_n 9.47434e-19 $X=1.947 $Y=0.935 $X2=0
+ $Y2=0
cc_398 D noxref_25 0.00135662f $X=1.595 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_399 N_SCD_M1011_g N_RESET_B_M1036_g 0.0322467f $X=3.04 $Y=0.615 $X2=0 $Y2=0
cc_400 SCD N_RESET_B_M1036_g 0.00220695f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_401 N_SCD_c_489_n N_RESET_B_M1036_g 0.0254311f $X=3.05 $Y=1.605 $X2=0 $Y2=0
cc_402 N_SCD_c_487_n N_RESET_B_c_899_n 0.0254311f $X=3.05 $Y=2.08 $X2=0 $Y2=0
cc_403 SCD N_RESET_B_c_899_n 0.00220695f $X=3.12 $Y=2.035 $X2=0 $Y2=0
cc_404 N_SCD_c_491_n N_RESET_B_c_905_n 0.016608f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_405 N_SCD_c_491_n N_VPWR_c_1745_n 0.0101332f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_406 N_SCD_c_491_n N_VPWR_c_1760_n 0.00413917f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_407 N_SCD_c_491_n N_VPWR_c_1744_n 0.00409757f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_408 N_SCD_M1011_g N_A_390_81#_c_1916_n 0.0257675f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_409 SCD N_A_390_81#_c_1916_n 0.0278904f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_410 N_SCD_c_489_n N_A_390_81#_c_1916_n 0.00381702f $X=3.05 $Y=1.605 $X2=0
+ $Y2=0
cc_411 N_SCD_c_491_n N_A_390_81#_c_1932_n 0.0177595f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_412 SCD N_A_390_81#_c_1932_n 0.0265196f $X=3.12 $Y=2.035 $X2=0 $Y2=0
cc_413 N_SCD_M1011_g N_A_390_81#_c_1917_n 0.0010027f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_414 N_SCD_c_491_n N_A_390_81#_c_1917_n 0.00199663f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_415 SCD N_A_390_81#_c_1917_n 0.0556356f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_416 N_SCD_c_489_n N_A_390_81#_c_1917_n 7.93612e-19 $X=3.05 $Y=1.605 $X2=0
+ $Y2=0
cc_417 N_SCD_c_491_n N_A_390_81#_c_1925_n 0.00104585f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_418 N_SCD_c_491_n N_A_390_81#_c_1931_n 0.00167743f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_419 N_SCD_M1011_g N_VGND_c_2103_n 9.15902e-19 $X=3.04 $Y=0.615 $X2=0 $Y2=0
cc_420 N_SCD_M1011_g N_noxref_24_c_2234_n 0.0101767f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_421 N_CLK_c_537_n N_A_1034_392#_c_607_n 2.73677e-19 $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_422 N_CLK_c_531_n N_A_1034_392#_c_588_n 8.03717e-19 $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_423 CLK N_RESET_B_M1036_g 0.00105038f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_424 N_CLK_c_535_n N_RESET_B_M1036_g 0.0433156f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_425 N_CLK_c_531_n N_RESET_B_c_891_n 0.0100076f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_426 CLK N_RESET_B_c_891_n 0.00336855f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_427 N_CLK_c_535_n N_RESET_B_c_891_n 0.00432122f $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_428 N_CLK_c_530_n N_RESET_B_c_898_n 0.0213192f $X=4.115 $Y=1.515 $X2=0 $Y2=0
cc_429 N_CLK_c_537_n N_RESET_B_c_898_n 0.00545707f $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_430 CLK N_RESET_B_c_898_n 0.00128901f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_431 CLK N_RESET_B_c_906_n 0.00634387f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_432 CLK N_RESET_B_c_907_n 0.00430124f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_433 N_CLK_c_530_n N_RESET_B_c_910_n 7.94102e-19 $X=4.115 $Y=1.515 $X2=0 $Y2=0
cc_434 N_CLK_c_537_n N_RESET_B_c_910_n 4.10028e-19 $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_435 CLK N_RESET_B_c_910_n 0.0269243f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_436 CLK N_A_835_98#_M1029_s 0.00349248f $X=3.995 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_437 N_CLK_c_537_n N_A_835_98#_c_1247_n 0.0374488f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_438 N_CLK_c_531_n N_A_835_98#_c_1236_n 0.0211616f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_439 N_CLK_c_531_n N_A_835_98#_c_1243_n 0.00445277f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_440 N_CLK_c_533_n N_A_835_98#_c_1243_n 3.29111e-19 $X=4.62 $Y=1.515 $X2=0
+ $Y2=0
cc_441 CLK N_A_835_98#_c_1243_n 0.0181996f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_442 N_CLK_c_529_n N_A_835_98#_c_1244_n 0.00113381f $X=4.52 $Y=1.515 $X2=0
+ $Y2=0
cc_443 N_CLK_c_531_n N_A_835_98#_c_1244_n 0.0264704f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_444 CLK N_A_835_98#_c_1244_n 0.0339329f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_445 N_CLK_c_535_n N_A_835_98#_c_1244_n 0.00116798f $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_446 N_CLK_c_529_n N_A_835_98#_c_1245_n 0.00133487f $X=4.52 $Y=1.515 $X2=0
+ $Y2=0
cc_447 N_CLK_c_533_n N_A_835_98#_c_1245_n 0.00633166f $X=4.62 $Y=1.515 $X2=0
+ $Y2=0
cc_448 N_CLK_c_537_n N_A_835_98#_c_1245_n 0.0196714f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_449 CLK N_A_835_98#_c_1245_n 0.036729f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_450 N_CLK_c_533_n N_A_835_98#_c_1246_n 0.0261328f $X=4.62 $Y=1.515 $X2=0
+ $Y2=0
cc_451 N_CLK_c_537_n N_VPWR_c_1746_n 0.0164315f $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_452 N_CLK_c_537_n N_VPWR_c_1753_n 0.00302783f $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_453 N_CLK_c_537_n N_VPWR_c_1744_n 0.00396658f $X=4.62 $Y=1.885 $X2=0 $Y2=0
cc_454 CLK N_A_390_81#_c_1916_n 0.0296573f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_455 N_CLK_c_535_n N_A_390_81#_c_1916_n 0.00120791f $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_456 CLK N_A_390_81#_c_1917_n 0.0287351f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_457 N_CLK_c_535_n N_A_390_81#_c_1917_n 0.00101712f $X=3.95 $Y=1.115 $X2=0
+ $Y2=0
cc_458 N_CLK_c_537_n N_A_390_81#_c_1924_n 0.0102356f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_459 N_CLK_c_537_n N_A_390_81#_c_1925_n 0.0094743f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_460 N_CLK_c_537_n N_A_390_81#_c_1926_n 0.00644616f $X=4.62 $Y=1.885 $X2=0
+ $Y2=0
cc_461 N_CLK_c_531_n N_VGND_c_2096_n 0.00155538f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_462 CLK N_VGND_c_2096_n 0.00799287f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_463 N_CLK_c_535_n N_VGND_c_2096_n 4.43186e-19 $X=3.95 $Y=1.115 $X2=0 $Y2=0
cc_464 N_CLK_c_531_n N_VGND_c_2097_n 0.00259354f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_465 N_CLK_c_531_n N_VGND_c_2118_n 9.39239e-19 $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_466 N_A_1034_392#_c_595_n N_A_1367_93#_M1035_d 0.00256812f $X=9.09 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_467 N_A_1034_392#_M1000_g N_A_1367_93#_M1019_g 0.0333609f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_468 N_A_1034_392#_c_590_n N_A_1367_93#_M1019_g 0.00344795f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_469 N_A_1034_392#_c_593_n N_A_1367_93#_M1019_g 0.00262964f $X=7.135 $Y=0.58
+ $X2=0 $Y2=0
cc_470 N_A_1034_392#_c_618_p N_A_1367_93#_M1019_g 0.0026982f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_471 N_A_1034_392#_c_603_n N_A_1367_93#_M1033_g 0.00334209f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_472 N_A_1034_392#_c_602_n N_A_1367_93#_M1033_g 7.41525e-19 $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_473 N_A_1034_392#_c_583_n N_A_1367_93#_c_792_n 0.0333609f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_474 N_A_1034_392#_c_602_n N_A_1367_93#_c_792_n 0.00108114f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_475 N_A_1034_392#_c_590_n N_A_1367_93#_c_793_n 5.94333e-19 $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_476 N_A_1034_392#_c_594_n N_A_1367_93#_c_793_n 0.00304701f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_477 N_A_1034_392#_c_618_p N_A_1367_93#_c_793_n 0.0103944f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_478 N_A_1034_392#_c_594_n N_A_1367_93#_c_794_n 0.0570369f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_479 N_A_1034_392#_c_595_n N_A_1367_93#_c_794_n 0.0055642f $X=9.09 $Y=0.34
+ $X2=0 $Y2=0
cc_480 N_A_1034_392#_c_594_n N_A_1367_93#_c_816_n 0.0138386f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_481 N_A_1034_392#_c_595_n N_A_1367_93#_c_816_n 0.0383715f $X=9.09 $Y=0.34
+ $X2=0 $Y2=0
cc_482 N_A_1034_392#_c_587_n N_A_1367_93#_c_800_n 0.00481612f $X=9.12 $Y=1.26
+ $X2=0 $Y2=0
cc_483 N_A_1034_392#_c_598_n N_A_1367_93#_c_800_n 0.0011706f $X=9.26 $Y=1.17
+ $X2=0 $Y2=0
cc_484 N_A_1034_392#_c_600_n N_A_1367_93#_c_800_n 0.00385352f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_485 N_A_1034_392#_c_585_n N_A_1367_93#_c_795_n 0.00223701f $X=9.045 $Y=1.185
+ $X2=0 $Y2=0
cc_486 N_A_1034_392#_c_598_n N_A_1367_93#_c_795_n 0.0187413f $X=9.26 $Y=1.17
+ $X2=0 $Y2=0
cc_487 N_A_1034_392#_M1000_g N_RESET_B_c_891_n 0.00882199f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_488 N_A_1034_392#_c_590_n N_RESET_B_c_891_n 0.0294278f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_489 N_A_1034_392#_c_591_n N_RESET_B_c_891_n 0.00992957f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_490 N_A_1034_392#_c_590_n N_RESET_B_M1009_g 0.00466687f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_491 N_A_1034_392#_c_593_n N_RESET_B_M1009_g 0.00445709f $X=7.135 $Y=0.58
+ $X2=0 $Y2=0
cc_492 N_A_1034_392#_c_594_n N_RESET_B_M1009_g 0.0128168f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_493 N_A_1034_392#_c_641_p N_RESET_B_M1009_g 0.0035287f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_494 N_A_1034_392#_c_596_n N_RESET_B_M1009_g 6.46496e-19 $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_495 N_A_1034_392#_c_603_n N_RESET_B_c_906_n 0.00315542f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_496 N_A_1034_392#_c_583_n N_RESET_B_c_906_n 0.00325193f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_497 N_A_1034_392#_c_607_n N_RESET_B_c_906_n 0.0144304f $X=5.45 $Y=2.085 $X2=0
+ $Y2=0
cc_498 N_A_1034_392#_c_608_n N_RESET_B_c_906_n 0.017308f $X=5.63 $Y=1.71 $X2=0
+ $Y2=0
cc_499 N_A_1034_392#_c_592_n N_RESET_B_c_906_n 0.0155597f $X=6.085 $Y=1.71 $X2=0
+ $Y2=0
cc_500 N_A_1034_392#_c_602_n N_RESET_B_c_906_n 0.00379596f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_501 N_A_1034_392#_c_586_n N_RESET_B_c_908_n 3.77242e-19 $X=9.48 $Y=1.26 $X2=0
+ $Y2=0
cc_502 N_A_1034_392#_c_606_n N_RESET_B_c_908_n 0.00339815f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_503 N_A_1034_392#_c_600_n N_RESET_B_c_908_n 0.0178906f $X=9.95 $Y=2.165 $X2=0
+ $Y2=0
cc_504 N_A_1034_392#_c_585_n N_A_1234_119#_M1035_g 0.0134624f $X=9.045 $Y=1.185
+ $X2=0 $Y2=0
cc_505 N_A_1034_392#_c_594_n N_A_1234_119#_M1035_g 0.00131978f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_506 N_A_1034_392#_c_641_p N_A_1234_119#_M1035_g 0.00428575f $X=8.015 $Y=0.58
+ $X2=0 $Y2=0
cc_507 N_A_1034_392#_c_595_n N_A_1234_119#_M1035_g 0.0113704f $X=9.09 $Y=0.34
+ $X2=0 $Y2=0
cc_508 N_A_1034_392#_c_656_p N_A_1234_119#_M1035_g 9.4741e-19 $X=9.175 $Y=1.005
+ $X2=0 $Y2=0
cc_509 N_A_1034_392#_c_587_n N_A_1234_119#_c_1111_n 0.0134624f $X=9.12 $Y=1.26
+ $X2=0 $Y2=0
cc_510 N_A_1034_392#_c_583_n N_A_1234_119#_c_1121_n 9.01642e-19 $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_511 N_A_1034_392#_M1000_g N_A_1234_119#_c_1113_n 0.0110407f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_512 N_A_1034_392#_c_590_n N_A_1234_119#_c_1113_n 0.0110883f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_513 N_A_1034_392#_M1000_g N_A_1234_119#_c_1114_n 0.0071804f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_514 N_A_1034_392#_c_583_n N_A_1234_119#_c_1118_n 6.46907e-19 $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_515 N_A_1034_392#_M1000_g N_A_1234_119#_c_1118_n 0.00636651f $X=6.525
+ $Y=0.805 $X2=0 $Y2=0
cc_516 N_A_1034_392#_c_590_n N_A_1234_119#_c_1118_n 0.019863f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_517 N_A_1034_392#_c_618_p N_A_1234_119#_c_1118_n 0.00486547f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_518 N_A_1034_392#_c_603_n N_A_1234_119#_c_1126_n 2.99618e-19 $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_519 N_A_1034_392#_c_607_n N_A_835_98#_c_1247_n 0.00258584f $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_520 N_A_1034_392#_c_608_n N_A_835_98#_c_1247_n 6.39872e-19 $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_521 N_A_1034_392#_c_588_n N_A_835_98#_c_1236_n 0.00987138f $X=5.36 $Y=0.78
+ $X2=0 $Y2=0
cc_522 N_A_1034_392#_c_589_n N_A_835_98#_c_1236_n 8.65367e-19 $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_523 N_A_1034_392#_c_601_n N_A_835_98#_c_1236_n 0.00191523f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_524 N_A_1034_392#_c_603_n N_A_835_98#_c_1248_n 0.0111007f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_525 N_A_1034_392#_c_604_n N_A_835_98#_c_1248_n 0.0130881f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_526 N_A_1034_392#_c_607_n N_A_835_98#_c_1248_n 4.97235e-19 $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_527 N_A_1034_392#_c_608_n N_A_835_98#_c_1248_n 0.0104193f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_528 N_A_1034_392#_c_604_n N_A_835_98#_c_1249_n 0.00899632f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_529 N_A_1034_392#_c_590_n N_A_835_98#_c_1237_n 0.00139627f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_530 N_A_1034_392#_c_592_n N_A_835_98#_c_1237_n 0.00441445f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_531 N_A_1034_392#_c_602_n N_A_835_98#_c_1237_n 0.0160947f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_532 N_A_1034_392#_M1000_g N_A_835_98#_c_1238_n 0.0223151f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_533 N_A_1034_392#_c_588_n N_A_835_98#_c_1238_n 0.00472785f $X=5.36 $Y=0.78
+ $X2=0 $Y2=0
cc_534 N_A_1034_392#_c_590_n N_A_835_98#_c_1238_n 0.00330666f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_535 N_A_1034_392#_c_604_n N_A_835_98#_M1008_g 0.0140799f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_536 N_A_1034_392#_c_583_n N_A_835_98#_M1008_g 0.00296839f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_537 N_A_1034_392#_c_606_n N_A_835_98#_M1018_g 0.001338f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_538 N_A_1034_392#_c_600_n N_A_835_98#_M1018_g 0.00134374f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_539 N_A_1034_392#_c_606_n N_A_835_98#_c_1239_n 0.0207729f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_540 N_A_1034_392#_c_599_n N_A_835_98#_c_1239_n 0.0169827f $X=9.645 $Y=1.17
+ $X2=0 $Y2=0
cc_541 N_A_1034_392#_c_600_n N_A_835_98#_c_1239_n 0.0202931f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_542 N_A_1034_392#_c_586_n N_A_835_98#_c_1255_n 0.0169827f $X=9.48 $Y=1.26
+ $X2=0 $Y2=0
cc_543 N_A_1034_392#_c_597_n N_A_835_98#_c_1255_n 0.00271869f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_544 N_A_1034_392#_c_598_n N_A_835_98#_c_1255_n 6.613e-19 $X=9.26 $Y=1.17
+ $X2=0 $Y2=0
cc_545 N_A_1034_392#_c_600_n N_A_835_98#_c_1255_n 5.48883e-19 $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_546 N_A_1034_392#_c_600_n N_A_835_98#_c_1240_n 0.00569302f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_547 N_A_1034_392#_c_606_n N_A_835_98#_c_1257_n 0.00415106f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_548 N_A_1034_392#_c_597_n N_A_835_98#_c_1242_n 0.00289132f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_549 N_A_1034_392#_c_599_n N_A_835_98#_c_1242_n 0.0181127f $X=9.645 $Y=1.17
+ $X2=0 $Y2=0
cc_550 N_A_1034_392#_c_589_n N_A_835_98#_c_1243_n 0.00563685f $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_551 N_A_1034_392#_c_588_n N_A_835_98#_c_1244_n 0.00231034f $X=5.36 $Y=0.78
+ $X2=0 $Y2=0
cc_552 N_A_1034_392#_c_607_n N_A_835_98#_c_1245_n 0.0199151f $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_553 N_A_1034_392#_c_589_n N_A_835_98#_c_1245_n 0.0236806f $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_554 N_A_1034_392#_c_608_n N_A_835_98#_c_1245_n 0.00658609f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_555 N_A_1034_392#_c_601_n N_A_835_98#_c_1245_n 0.00267749f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_556 N_A_1034_392#_c_607_n N_A_835_98#_c_1246_n 0.00634613f $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_557 N_A_1034_392#_c_589_n N_A_835_98#_c_1246_n 0.0141907f $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_558 N_A_1034_392#_c_590_n N_A_835_98#_c_1246_n 0.00385788f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_559 N_A_1034_392#_c_608_n N_A_835_98#_c_1246_n 0.0120306f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_560 N_A_1034_392#_c_592_n N_A_835_98#_c_1246_n 0.0116804f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_561 N_A_1034_392#_c_601_n N_A_835_98#_c_1246_n 0.0122529f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_562 N_A_1034_392#_c_602_n N_A_835_98#_c_1246_n 0.021574f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_563 N_A_1034_392#_c_606_n N_A_2082_446#_c_1425_n 0.0313578f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_564 N_A_1034_392#_c_606_n N_A_2082_446#_c_1426_n 0.0134605f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_565 N_A_1034_392#_c_606_n N_A_2082_446#_c_1417_n 0.0127423f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_566 N_A_1034_392#_c_595_n N_A_1824_74#_M1016_d 0.00248108f $X=9.09 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_567 N_A_1034_392#_c_656_p N_A_1824_74#_M1016_d 0.0130256f $X=9.175 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_568 N_A_1034_392#_c_597_n N_A_1824_74#_M1016_d 0.00450592f $X=9.785 $Y=1.17
+ $X2=-0.19 $Y2=-0.245
cc_569 N_A_1034_392#_c_606_n N_A_1824_74#_c_1563_n 0.004427f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_570 N_A_1034_392#_c_597_n N_A_1824_74#_c_1563_n 0.00861974f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_571 N_A_1034_392#_c_600_n N_A_1824_74#_c_1563_n 0.0339543f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_572 N_A_1034_392#_c_585_n N_A_1824_74#_c_1545_n 0.0018748f $X=9.045 $Y=1.185
+ $X2=0 $Y2=0
cc_573 N_A_1034_392#_c_586_n N_A_1824_74#_c_1545_n 2.42458e-19 $X=9.48 $Y=1.26
+ $X2=0 $Y2=0
cc_574 N_A_1034_392#_c_656_p N_A_1824_74#_c_1545_n 0.026719f $X=9.175 $Y=1.005
+ $X2=0 $Y2=0
cc_575 N_A_1034_392#_c_597_n N_A_1824_74#_c_1545_n 0.0466861f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_576 N_A_1034_392#_c_599_n N_A_1824_74#_c_1545_n 0.0070276f $X=9.645 $Y=1.17
+ $X2=0 $Y2=0
cc_577 N_A_1034_392#_c_606_n N_A_1824_74#_c_1557_n 0.0157095f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_578 N_A_1034_392#_c_600_n N_A_1824_74#_c_1557_n 0.019012f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_579 N_A_1034_392#_c_597_n N_A_1824_74#_c_1546_n 0.00187033f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_580 N_A_1034_392#_c_606_n N_A_1824_74#_c_1547_n 0.00479636f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_581 N_A_1034_392#_c_597_n N_A_1824_74#_c_1547_n 0.0107493f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_582 N_A_1034_392#_c_600_n N_A_1824_74#_c_1547_n 0.0746733f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_583 N_A_1034_392#_c_597_n N_A_1824_74#_c_1549_n 0.0146626f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_584 N_A_1034_392#_c_606_n N_VPWR_c_1762_n 0.00308386f $X=10.11 $Y=2.465 $X2=0
+ $Y2=0
cc_585 N_A_1034_392#_c_606_n N_VPWR_c_1768_n 0.0012612f $X=10.11 $Y=2.465 $X2=0
+ $Y2=0
cc_586 N_A_1034_392#_c_604_n N_VPWR_c_1744_n 9.49986e-19 $X=6.135 $Y=2.21 $X2=0
+ $Y2=0
cc_587 N_A_1034_392#_c_606_n N_VPWR_c_1744_n 0.00381714f $X=10.11 $Y=2.465 $X2=0
+ $Y2=0
cc_588 N_A_1034_392#_M1030_d N_A_390_81#_c_1926_n 0.00695361f $X=5.17 $Y=1.96
+ $X2=0 $Y2=0
cc_589 N_A_1034_392#_c_607_n N_A_390_81#_c_1926_n 0.016647f $X=5.45 $Y=2.085
+ $X2=0 $Y2=0
cc_590 N_A_1034_392#_c_608_n N_A_390_81#_c_1926_n 0.0134529f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_591 N_A_1034_392#_c_592_n N_A_390_81#_c_1926_n 0.0029069f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_592 N_A_1034_392#_c_588_n N_A_390_81#_c_1918_n 0.0311322f $X=5.36 $Y=0.78
+ $X2=0 $Y2=0
cc_593 N_A_1034_392#_c_590_n N_A_390_81#_c_1918_n 0.013349f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_594 N_A_1034_392#_M1000_g N_A_390_81#_c_1919_n 3.66002e-19 $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_595 N_A_1034_392#_c_588_n N_A_390_81#_c_1919_n 0.00571418f $X=5.36 $Y=0.78
+ $X2=0 $Y2=0
cc_596 N_A_1034_392#_c_601_n N_A_390_81#_c_1919_n 0.00980399f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_597 N_A_1034_392#_c_604_n N_A_390_81#_c_1927_n 0.00783906f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_598 N_A_1034_392#_M1000_g N_A_390_81#_c_1920_n 0.00551398f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_599 N_A_1034_392#_c_592_n N_A_390_81#_c_1920_n 0.0142722f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_600 N_A_1034_392#_c_602_n N_A_390_81#_c_1920_n 0.00577594f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_601 N_A_1034_392#_c_592_n N_A_390_81#_c_1921_n 0.0145081f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_602 N_A_1034_392#_c_601_n N_A_390_81#_c_1921_n 0.013579f $X=5.422 $Y=1.285
+ $X2=0 $Y2=0
cc_603 N_A_1034_392#_c_602_n N_A_390_81#_c_1921_n 3.38485e-19 $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_604 N_A_1034_392#_c_603_n N_A_390_81#_c_1928_n 0.00390532f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_605 N_A_1034_392#_c_604_n N_A_390_81#_c_1928_n 0.00843492f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_606 N_A_1034_392#_c_583_n N_A_390_81#_c_1928_n 0.00177679f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_607 N_A_1034_392#_c_592_n N_A_390_81#_c_1928_n 0.00615957f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_608 N_A_1034_392#_c_602_n N_A_390_81#_c_1928_n 6.46491e-19 $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_609 N_A_1034_392#_c_603_n N_A_390_81#_c_1929_n 0.00121768f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_610 N_A_1034_392#_c_604_n N_A_390_81#_c_1929_n 0.00154832f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_611 N_A_1034_392#_c_608_n N_A_390_81#_c_1929_n 0.0116706f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_612 N_A_1034_392#_c_592_n N_A_390_81#_c_1929_n 0.016874f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_613 N_A_1034_392#_c_602_n N_A_390_81#_c_1929_n 0.00278662f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_614 N_A_1034_392#_c_603_n N_A_390_81#_c_1922_n 0.00400586f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_615 N_A_1034_392#_c_583_n N_A_390_81#_c_1922_n 0.0122247f $X=6.45 $Y=1.635
+ $X2=0 $Y2=0
cc_616 N_A_1034_392#_M1000_g N_A_390_81#_c_1922_n 0.00504469f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_617 N_A_1034_392#_c_592_n N_A_390_81#_c_1922_n 0.0250842f $X=6.085 $Y=1.71
+ $X2=0 $Y2=0
cc_618 N_A_1034_392#_c_602_n N_A_390_81#_c_1922_n 0.00171299f $X=6.085 $Y=1.635
+ $X2=0 $Y2=0
cc_619 N_A_1034_392#_c_594_n N_VGND_M1009_d 0.0193371f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_620 N_A_1034_392#_c_641_p N_VGND_M1009_d 0.00598032f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_621 N_A_1034_392#_c_595_n N_VGND_M1009_d 0.00505669f $X=9.09 $Y=0.34 $X2=0
+ $Y2=0
cc_622 N_A_1034_392#_c_596_n N_VGND_M1009_d 0.00120457f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_623 N_A_1034_392#_c_588_n N_VGND_c_2097_n 0.0174236f $X=5.36 $Y=0.78 $X2=0
+ $Y2=0
cc_624 N_A_1034_392#_c_591_n N_VGND_c_2097_n 0.0144411f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_625 N_A_1034_392#_c_590_n N_VGND_c_2108_n 0.103356f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_626 N_A_1034_392#_c_591_n N_VGND_c_2108_n 0.0276098f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_627 N_A_1034_392#_c_594_n N_VGND_c_2108_n 0.00402072f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_628 N_A_1034_392#_c_585_n N_VGND_c_2109_n 0.00278242f $X=9.045 $Y=1.185 $X2=0
+ $Y2=0
cc_629 N_A_1034_392#_c_594_n N_VGND_c_2109_n 0.00335833f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_630 N_A_1034_392#_c_595_n N_VGND_c_2109_n 0.0750141f $X=9.09 $Y=0.34 $X2=0
+ $Y2=0
cc_631 N_A_1034_392#_c_596_n N_VGND_c_2109_n 0.0118998f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_632 N_A_1034_392#_c_590_n N_VGND_c_2114_n 0.0118008f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_633 N_A_1034_392#_c_594_n N_VGND_c_2114_n 0.0246154f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_634 N_A_1034_392#_c_596_n N_VGND_c_2114_n 0.0135796f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_635 N_A_1034_392#_c_585_n N_VGND_c_2118_n 0.00359177f $X=9.045 $Y=1.185 $X2=0
+ $Y2=0
cc_636 N_A_1034_392#_c_590_n N_VGND_c_2118_n 0.0538367f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_637 N_A_1034_392#_c_591_n N_VGND_c_2118_n 0.0138923f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_638 N_A_1034_392#_c_594_n N_VGND_c_2118_n 0.0122484f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_639 N_A_1034_392#_c_595_n N_VGND_c_2118_n 0.0424576f $X=9.09 $Y=0.34 $X2=0
+ $Y2=0
cc_640 N_A_1034_392#_c_596_n N_VGND_c_2118_n 0.00655543f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_641 N_A_1034_392#_c_618_p A_1397_119# 0.00349303f $X=7.22 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_642 N_A_1367_93#_M1019_g N_RESET_B_c_891_n 0.00882199f $X=6.91 $Y=0.805 $X2=0
+ $Y2=0
cc_643 N_A_1367_93#_c_793_n N_RESET_B_c_891_n 2.57602e-19 $X=7.265 $Y=1.005
+ $X2=0 $Y2=0
cc_644 N_A_1367_93#_M1019_g N_RESET_B_M1009_g 0.0398547f $X=6.91 $Y=0.805 $X2=0
+ $Y2=0
cc_645 N_A_1367_93#_c_791_n N_RESET_B_M1009_g 0.00116633f $X=7.145 $Y=1.64 $X2=0
+ $Y2=0
cc_646 N_A_1367_93#_c_793_n N_RESET_B_M1009_g 0.00250892f $X=7.265 $Y=1.005
+ $X2=0 $Y2=0
cc_647 N_A_1367_93#_c_794_n N_RESET_B_M1009_g 0.0104334f $X=8.27 $Y=0.842 $X2=0
+ $Y2=0
cc_648 N_A_1367_93#_M1019_g N_RESET_B_c_894_n 0.00178049f $X=6.91 $Y=0.805 $X2=0
+ $Y2=0
cc_649 N_A_1367_93#_c_791_n N_RESET_B_c_894_n 7.18471e-19 $X=7.145 $Y=1.64 $X2=0
+ $Y2=0
cc_650 N_A_1367_93#_c_792_n N_RESET_B_c_894_n 0.0209381f $X=7.145 $Y=1.64 $X2=0
+ $Y2=0
cc_651 N_A_1367_93#_c_791_n N_RESET_B_c_896_n 0.00822559f $X=7.145 $Y=1.64 $X2=0
+ $Y2=0
cc_652 N_A_1367_93#_c_792_n N_RESET_B_c_896_n 0.0059618f $X=7.145 $Y=1.64 $X2=0
+ $Y2=0
cc_653 N_A_1367_93#_c_794_n N_RESET_B_c_896_n 0.00903119f $X=8.27 $Y=0.842 $X2=0
+ $Y2=0
cc_654 N_A_1367_93#_M1033_g N_RESET_B_c_906_n 0.0065779f $X=6.945 $Y=2.495 $X2=0
+ $Y2=0
cc_655 N_A_1367_93#_c_791_n N_RESET_B_c_906_n 0.00621585f $X=7.145 $Y=1.64 $X2=0
+ $Y2=0
cc_656 N_A_1367_93#_c_792_n N_RESET_B_c_906_n 0.00171088f $X=7.145 $Y=1.64 $X2=0
+ $Y2=0
cc_657 N_A_1367_93#_M1015_d N_RESET_B_c_908_n 0.00622796f $X=8.715 $Y=1.735
+ $X2=0 $Y2=0
cc_658 N_A_1367_93#_c_799_n N_RESET_B_c_908_n 0.0432512f $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_659 N_A_1367_93#_c_799_n N_RESET_B_c_966_n 6.64095e-19 $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_660 N_A_1367_93#_c_799_n N_RESET_B_c_909_n 0.0153091f $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_661 N_A_1367_93#_M1033_g N_RESET_B_c_911_n 0.0207015f $X=6.945 $Y=2.495 $X2=0
+ $Y2=0
cc_662 N_A_1367_93#_c_816_n N_A_1234_119#_M1035_g 0.0268444f $X=8.835 $Y=0.842
+ $X2=0 $Y2=0
cc_663 N_A_1367_93#_c_795_n N_A_1234_119#_M1035_g 0.00696321f $X=8.932 $Y=1.715
+ $X2=0 $Y2=0
cc_664 N_A_1367_93#_c_816_n N_A_1234_119#_c_1111_n 0.00334118f $X=8.835 $Y=0.842
+ $X2=0 $Y2=0
cc_665 N_A_1367_93#_c_795_n N_A_1234_119#_c_1111_n 0.0167422f $X=8.932 $Y=1.715
+ $X2=0 $Y2=0
cc_666 N_A_1367_93#_c_794_n N_A_1234_119#_c_1112_n 0.00849203f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_667 N_A_1367_93#_M1033_g N_A_1234_119#_c_1121_n 0.00128347f $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_668 N_A_1367_93#_M1019_g N_A_1234_119#_c_1113_n 0.00419324f $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_669 N_A_1367_93#_c_793_n N_A_1234_119#_c_1113_n 0.00492865f $X=7.265 $Y=1.005
+ $X2=0 $Y2=0
cc_670 N_A_1367_93#_M1019_g N_A_1234_119#_c_1114_n 0.00722399f $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_671 N_A_1367_93#_M1033_g N_A_1234_119#_c_1114_n 0.00308621f $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_672 N_A_1367_93#_c_791_n N_A_1234_119#_c_1114_n 0.0512142f $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_673 N_A_1367_93#_c_792_n N_A_1234_119#_c_1114_n 0.00805995f $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_674 N_A_1367_93#_c_793_n N_A_1234_119#_c_1114_n 0.00480618f $X=7.265 $Y=1.005
+ $X2=0 $Y2=0
cc_675 N_A_1367_93#_M1033_g N_A_1234_119#_c_1123_n 0.00178971f $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_676 N_A_1367_93#_M1033_g N_A_1234_119#_c_1124_n 0.0175598f $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_677 N_A_1367_93#_c_791_n N_A_1234_119#_c_1124_n 0.0155534f $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_678 N_A_1367_93#_c_792_n N_A_1234_119#_c_1124_n 0.00383298f $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_679 N_A_1367_93#_M1033_g N_A_1234_119#_c_1115_n 0.00183154f $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_680 N_A_1367_93#_c_791_n N_A_1234_119#_c_1115_n 0.0190372f $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_681 N_A_1367_93#_c_792_n N_A_1234_119#_c_1115_n 0.00157419f $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_682 N_A_1367_93#_c_791_n N_A_1234_119#_c_1116_n 0.0243296f $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_683 N_A_1367_93#_c_792_n N_A_1234_119#_c_1116_n 4.90401e-19 $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_684 N_A_1367_93#_c_794_n N_A_1234_119#_c_1116_n 0.0135838f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_685 N_A_1367_93#_c_794_n N_A_1234_119#_c_1117_n 0.0655079f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_686 N_A_1367_93#_c_795_n N_A_1234_119#_c_1117_n 0.0161785f $X=8.932 $Y=1.715
+ $X2=0 $Y2=0
cc_687 N_A_1367_93#_M1019_g N_A_1234_119#_c_1118_n 0.00107025f $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_688 N_A_1367_93#_M1033_g N_A_1234_119#_c_1128_n 6.64763e-19 $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_689 N_A_1367_93#_M1033_g N_A_835_98#_M1008_g 0.0385033f $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_690 N_A_1367_93#_M1033_g N_A_835_98#_c_1252_n 0.00907339f $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_691 N_A_1367_93#_c_799_n N_A_835_98#_c_1252_n 0.00737375f $X=8.95 $Y=2.235
+ $X2=0 $Y2=0
cc_692 N_A_1367_93#_c_800_n N_A_835_98#_M1018_g 0.0104192f $X=8.95 $Y=1.88 $X2=0
+ $Y2=0
cc_693 N_A_1367_93#_c_800_n N_A_835_98#_c_1255_n 7.1022e-19 $X=8.95 $Y=1.88
+ $X2=0 $Y2=0
cc_694 N_A_1367_93#_c_795_n N_A_835_98#_c_1255_n 0.00307401f $X=8.932 $Y=1.715
+ $X2=0 $Y2=0
cc_695 N_A_1367_93#_c_800_n N_A_1824_74#_c_1563_n 0.0438134f $X=8.95 $Y=1.88
+ $X2=0 $Y2=0
cc_696 N_A_1367_93#_c_799_n N_A_1824_74#_c_1558_n 0.0168727f $X=8.95 $Y=2.235
+ $X2=0 $Y2=0
cc_697 N_A_1367_93#_M1033_g N_VPWR_c_1747_n 0.0033811f $X=6.945 $Y=2.495 $X2=0
+ $Y2=0
cc_698 N_A_1367_93#_c_799_n N_VPWR_c_1748_n 0.0167864f $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_699 N_A_1367_93#_c_799_n N_VPWR_c_1762_n 0.00805754f $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_700 N_A_1367_93#_M1033_g N_VPWR_c_1744_n 9.49986e-19 $X=6.945 $Y=2.495 $X2=0
+ $Y2=0
cc_701 N_A_1367_93#_c_799_n N_VPWR_c_1744_n 0.0100713f $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_702 N_A_1367_93#_M1033_g N_A_390_81#_c_1928_n 3.2345e-19 $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_703 N_A_1367_93#_M1019_g N_A_390_81#_c_1922_n 3.00253e-19 $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_704 N_A_1367_93#_M1033_g N_A_390_81#_c_1922_n 3.97102e-19 $X=6.945 $Y=2.495
+ $X2=0 $Y2=0
cc_705 N_A_1367_93#_c_792_n N_A_390_81#_c_1922_n 2.16488e-19 $X=7.145 $Y=1.64
+ $X2=0 $Y2=0
cc_706 N_A_1367_93#_c_794_n N_VGND_M1009_d 0.0145119f $X=8.27 $Y=0.842 $X2=0
+ $Y2=0
cc_707 N_A_1367_93#_c_816_n N_VGND_M1009_d 0.0123681f $X=8.835 $Y=0.842 $X2=0
+ $Y2=0
cc_708 N_A_1367_93#_c_793_n A_1397_119# 0.00138862f $X=7.265 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_709 N_RESET_B_c_908_n N_A_1234_119#_c_1111_n 0.012888f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_710 N_RESET_B_c_909_n N_A_1234_119#_c_1111_n 0.00953577f $X=8.4 $Y=2.035
+ $X2=0 $Y2=0
cc_711 N_RESET_B_c_911_n N_A_1234_119#_c_1111_n 0.00589904f $X=7.595 $Y=2.002
+ $X2=0 $Y2=0
cc_712 N_RESET_B_c_896_n N_A_1234_119#_c_1112_n 0.00901141f $X=7.595 $Y=1.19
+ $X2=0 $Y2=0
cc_713 N_RESET_B_c_909_n N_A_1234_119#_c_1112_n 0.0108866f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_714 N_RESET_B_c_906_n N_A_1234_119#_c_1121_n 0.00849024f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_715 N_RESET_B_M1009_g N_A_1234_119#_c_1113_n 3.7607e-19 $X=7.3 $Y=0.805 $X2=0
+ $Y2=0
cc_716 N_RESET_B_c_906_n N_A_1234_119#_c_1114_n 0.00946491f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_717 N_RESET_B_c_906_n N_A_1234_119#_c_1124_n 0.0312549f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_718 N_RESET_B_c_911_n N_A_1234_119#_c_1124_n 0.0100553f $X=7.595 $Y=2.002
+ $X2=0 $Y2=0
cc_719 N_RESET_B_c_894_n N_A_1234_119#_c_1115_n 0.0115547f $X=7.595 $Y=1.795
+ $X2=0 $Y2=0
cc_720 N_RESET_B_c_906_n N_A_1234_119#_c_1115_n 0.00996661f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_721 N_RESET_B_c_909_n N_A_1234_119#_c_1115_n 0.014155f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_722 N_RESET_B_c_911_n N_A_1234_119#_c_1115_n 0.00515774f $X=7.595 $Y=2.002
+ $X2=0 $Y2=0
cc_723 N_RESET_B_c_894_n N_A_1234_119#_c_1116_n 0.00374691f $X=7.595 $Y=1.795
+ $X2=0 $Y2=0
cc_724 N_RESET_B_c_896_n N_A_1234_119#_c_1116_n 0.00371515f $X=7.595 $Y=1.19
+ $X2=0 $Y2=0
cc_725 N_RESET_B_c_894_n N_A_1234_119#_c_1117_n 0.00744469f $X=7.595 $Y=1.795
+ $X2=0 $Y2=0
cc_726 N_RESET_B_c_896_n N_A_1234_119#_c_1117_n 5.9918e-19 $X=7.595 $Y=1.19
+ $X2=0 $Y2=0
cc_727 N_RESET_B_c_906_n N_A_1234_119#_c_1117_n 0.00811442f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_728 N_RESET_B_c_966_n N_A_1234_119#_c_1117_n 0.00122923f $X=8.545 $Y=2.035
+ $X2=0 $Y2=0
cc_729 N_RESET_B_c_909_n N_A_1234_119#_c_1117_n 0.0376394f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_730 N_RESET_B_c_911_n N_A_1234_119#_c_1117_n 0.00934295f $X=7.595 $Y=2.002
+ $X2=0 $Y2=0
cc_731 N_RESET_B_c_906_n N_A_1234_119#_c_1126_n 0.0126021f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_732 N_RESET_B_c_906_n N_A_1234_119#_c_1194_n 0.0124953f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_733 N_RESET_B_c_909_n N_A_1234_119#_c_1194_n 0.0117249f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_734 N_RESET_B_c_911_n N_A_1234_119#_c_1194_n 0.00691511f $X=7.595 $Y=2.002
+ $X2=0 $Y2=0
cc_735 N_RESET_B_c_900_n N_A_1234_119#_c_1127_n 0.00633065f $X=7.395 $Y=2.21
+ $X2=0 $Y2=0
cc_736 N_RESET_B_c_906_n N_A_1234_119#_c_1127_n 0.00702421f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_737 N_RESET_B_c_911_n N_A_1234_119#_c_1127_n 0.00724773f $X=7.595 $Y=2.002
+ $X2=0 $Y2=0
cc_738 N_RESET_B_c_900_n N_A_1234_119#_c_1128_n 0.00390298f $X=7.395 $Y=2.21
+ $X2=0 $Y2=0
cc_739 N_RESET_B_c_911_n N_A_1234_119#_c_1128_n 0.00611895f $X=7.595 $Y=2.002
+ $X2=0 $Y2=0
cc_740 N_RESET_B_c_906_n N_A_835_98#_M1028_s 0.00114217f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_741 N_RESET_B_c_906_n N_A_835_98#_c_1247_n 0.00350083f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_742 N_RESET_B_c_891_n N_A_835_98#_c_1236_n 0.0103973f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_743 N_RESET_B_c_906_n N_A_835_98#_c_1248_n 0.00218847f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_744 N_RESET_B_c_891_n N_A_835_98#_c_1238_n 0.00882199f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_745 N_RESET_B_c_906_n N_A_835_98#_M1008_g 0.00325607f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_746 N_RESET_B_c_900_n N_A_835_98#_c_1252_n 0.00889176f $X=7.395 $Y=2.21 $X2=0
+ $Y2=0
cc_747 N_RESET_B_c_908_n N_A_835_98#_M1018_g 0.00944311f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_748 N_RESET_B_c_908_n N_A_835_98#_c_1239_n 0.00577012f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_749 N_RESET_B_c_908_n N_A_835_98#_c_1255_n 3.19444e-19 $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_750 N_RESET_B_M1036_g N_A_835_98#_c_1244_n 0.00203097f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_751 N_RESET_B_c_891_n N_A_835_98#_c_1244_n 0.00943182f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_752 N_RESET_B_c_898_n N_A_835_98#_c_1245_n 0.0011403f $X=3.93 $Y=1.995 $X2=0
+ $Y2=0
cc_753 N_RESET_B_c_899_n N_A_835_98#_c_1245_n 0.00130059f $X=3.695 $Y=1.995
+ $X2=0 $Y2=0
cc_754 N_RESET_B_c_906_n N_A_835_98#_c_1245_n 0.046775f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_755 N_RESET_B_c_907_n N_A_835_98#_c_1245_n 0.00284227f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_756 N_RESET_B_c_910_n N_A_835_98#_c_1245_n 0.0281559f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_757 N_RESET_B_c_906_n N_A_835_98#_c_1246_n 0.00151487f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_758 N_RESET_B_c_904_n N_A_2082_446#_c_1425_n 0.00549853f $X=11.35 $Y=2.465
+ $X2=0 $Y2=0
cc_759 N_RESET_B_M1014_g N_A_2082_446#_M1003_g 0.0332604f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_760 N_RESET_B_c_903_n N_A_2082_446#_c_1426_n 0.00482347f $X=11.35 $Y=2.375
+ $X2=0 $Y2=0
cc_761 N_RESET_B_c_904_n N_A_2082_446#_c_1426_n 9.24257e-19 $X=11.35 $Y=2.465
+ $X2=0 $Y2=0
cc_762 N_RESET_B_c_908_n N_A_2082_446#_c_1426_n 7.79989e-19 $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_763 N_RESET_B_c_903_n N_A_2082_446#_c_1439_n 8.40443e-19 $X=11.35 $Y=2.375
+ $X2=0 $Y2=0
cc_764 N_RESET_B_c_908_n N_A_2082_446#_c_1439_n 0.0371304f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_765 RESET_B N_A_2082_446#_c_1439_n 5.86564e-19 $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_766 N_RESET_B_c_912_n N_A_2082_446#_c_1439_n 0.00153537f $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_767 N_RESET_B_c_1027_p N_A_2082_446#_c_1439_n 0.0134652f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_768 N_RESET_B_c_908_n N_A_2082_446#_c_1417_n 0.0118555f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_769 N_RESET_B_c_912_n N_A_2082_446#_c_1417_n 0.031607f $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_770 N_RESET_B_c_1027_p N_A_2082_446#_c_1417_n 0.00107974f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_771 N_RESET_B_M1014_g N_A_2082_446#_c_1418_n 0.0112646f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_772 N_RESET_B_c_908_n N_A_2082_446#_c_1418_n 0.00766736f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_773 RESET_B N_A_2082_446#_c_1418_n 0.0021857f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_774 N_RESET_B_c_912_n N_A_2082_446#_c_1418_n 0.00565198f $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_775 N_RESET_B_c_1027_p N_A_2082_446#_c_1418_n 0.0208148f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_776 N_RESET_B_c_904_n N_A_2082_446#_c_1429_n 0.0137666f $X=11.35 $Y=2.465
+ $X2=0 $Y2=0
cc_777 N_RESET_B_c_908_n N_A_2082_446#_c_1429_n 0.00726729f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_778 RESET_B N_A_2082_446#_c_1429_n 0.00176886f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_779 N_RESET_B_c_912_n N_A_2082_446#_c_1429_n 0.00469264f $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_780 N_RESET_B_c_1027_p N_A_2082_446#_c_1429_n 0.0223172f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_781 N_RESET_B_c_904_n N_A_2082_446#_c_1430_n 0.0102517f $X=11.35 $Y=2.465
+ $X2=0 $Y2=0
cc_782 N_RESET_B_M1014_g N_A_2082_446#_c_1419_n 0.00114233f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_783 N_RESET_B_M1014_g N_A_2082_446#_c_1421_n 7.54334e-19 $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_784 N_RESET_B_M1014_g N_A_2082_446#_c_1423_n 0.00211977f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_785 N_RESET_B_M1014_g N_A_2082_446#_c_1424_n 0.0225188f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_786 N_RESET_B_c_908_n N_A_1824_74#_M1018_d 6.85563e-19 $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_787 N_RESET_B_M1014_g N_A_1824_74#_M1007_g 0.0603983f $X=11.135 $Y=0.58 $X2=0
+ $Y2=0
cc_788 N_RESET_B_M1014_g N_A_1824_74#_c_1552_n 0.00632307f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_789 N_RESET_B_c_912_n N_A_1824_74#_c_1553_n 0.013294f $X=11.275 $Y=2.07 $X2=0
+ $Y2=0
cc_790 N_RESET_B_c_1027_p N_A_1824_74#_c_1553_n 0.00121903f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_791 N_RESET_B_c_903_n N_A_1824_74#_c_1554_n 0.013294f $X=11.35 $Y=2.375 $X2=0
+ $Y2=0
cc_792 N_RESET_B_c_904_n N_A_1824_74#_c_1554_n 0.00940262f $X=11.35 $Y=2.465
+ $X2=0 $Y2=0
cc_793 N_RESET_B_M1014_g N_A_1824_74#_c_1540_n 0.00629822f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_794 N_RESET_B_c_912_n N_A_1824_74#_c_1540_n 2.27226e-19 $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_795 N_RESET_B_M1014_g N_A_1824_74#_c_1543_n 0.00585373f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_796 N_RESET_B_c_908_n N_A_1824_74#_c_1563_n 0.0283424f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_797 N_RESET_B_c_908_n N_A_1824_74#_c_1557_n 0.0138963f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_798 N_RESET_B_c_908_n N_A_1824_74#_c_1547_n 0.023417f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_799 N_RESET_B_M1014_g N_A_1824_74#_c_1548_n 0.00517953f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_800 N_RESET_B_M1014_g N_A_1824_74#_c_1551_n 0.0159185f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_801 N_RESET_B_c_906_n N_VPWR_M1028_d 5.797e-19 $X=8.255 $Y=2.035 $X2=0 $Y2=0
cc_802 N_RESET_B_c_966_n N_VPWR_M1015_s 0.00198868f $X=8.545 $Y=2.035 $X2=0
+ $Y2=0
cc_803 N_RESET_B_c_909_n N_VPWR_M1015_s 0.00592726f $X=8.4 $Y=2.035 $X2=0 $Y2=0
cc_804 N_RESET_B_c_905_n N_VPWR_c_1745_n 0.0054851f $X=3.56 $Y=2.245 $X2=0 $Y2=0
cc_805 N_RESET_B_c_900_n N_VPWR_c_1747_n 0.00279283f $X=7.395 $Y=2.21 $X2=0
+ $Y2=0
cc_806 N_RESET_B_c_906_n N_VPWR_c_1747_n 0.00177009f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_807 N_RESET_B_c_908_n N_VPWR_c_1748_n 5.59089e-19 $X=11.135 $Y=2.035 $X2=0
+ $Y2=0
cc_808 N_RESET_B_c_966_n N_VPWR_c_1748_n 0.00820672f $X=8.545 $Y=2.035 $X2=0
+ $Y2=0
cc_809 N_RESET_B_c_909_n N_VPWR_c_1748_n 0.0187314f $X=8.4 $Y=2.035 $X2=0 $Y2=0
cc_810 RESET_B N_VPWR_c_1749_n 0.00143958f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_811 N_RESET_B_c_1027_p N_VPWR_c_1749_n 0.00812957f $X=11.28 $Y=2.035 $X2=0
+ $Y2=0
cc_812 N_RESET_B_c_905_n N_VPWR_c_1753_n 0.00387819f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_813 N_RESET_B_c_904_n N_VPWR_c_1757_n 0.00445602f $X=11.35 $Y=2.465 $X2=0
+ $Y2=0
cc_814 N_RESET_B_c_904_n N_VPWR_c_1768_n 0.00638397f $X=11.35 $Y=2.465 $X2=0
+ $Y2=0
cc_815 N_RESET_B_c_900_n N_VPWR_c_1744_n 9.49986e-19 $X=7.395 $Y=2.21 $X2=0
+ $Y2=0
cc_816 N_RESET_B_c_904_n N_VPWR_c_1744_n 0.00439026f $X=11.35 $Y=2.465 $X2=0
+ $Y2=0
cc_817 N_RESET_B_c_905_n N_VPWR_c_1744_n 0.00421415f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_818 N_RESET_B_M1036_g N_A_390_81#_c_1916_n 0.0207344f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_819 N_RESET_B_c_899_n N_A_390_81#_c_1932_n 8.77027e-19 $X=3.695 $Y=1.995
+ $X2=0 $Y2=0
cc_820 N_RESET_B_M1036_g N_A_390_81#_c_1917_n 0.0135694f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_821 N_RESET_B_c_899_n N_A_390_81#_c_1917_n 0.0185734f $X=3.695 $Y=1.995 $X2=0
+ $Y2=0
cc_822 N_RESET_B_c_905_n N_A_390_81#_c_1917_n 0.00445911f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_823 N_RESET_B_c_907_n N_A_390_81#_c_1917_n 0.00108729f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_824 N_RESET_B_c_910_n N_A_390_81#_c_1917_n 0.0243953f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_825 N_RESET_B_c_906_n N_A_390_81#_c_1924_n 0.00515092f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_826 N_RESET_B_c_898_n N_A_390_81#_c_1925_n 0.00525694f $X=3.93 $Y=1.995 $X2=0
+ $Y2=0
cc_827 N_RESET_B_c_905_n N_A_390_81#_c_1925_n 0.0198966f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_828 N_RESET_B_c_906_n N_A_390_81#_c_1925_n 0.00101627f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_829 N_RESET_B_c_907_n N_A_390_81#_c_1925_n 0.00440614f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_830 N_RESET_B_c_910_n N_A_390_81#_c_1925_n 0.0258211f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_831 N_RESET_B_c_906_n N_A_390_81#_c_1926_n 0.0137461f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_832 N_RESET_B_c_906_n N_A_390_81#_c_1920_n 0.00348472f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_833 N_RESET_B_c_906_n N_A_390_81#_c_1928_n 0.0172886f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_834 N_RESET_B_c_906_n N_A_390_81#_c_1929_n 0.0167671f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_835 N_RESET_B_c_906_n N_A_390_81#_c_1922_n 0.00940891f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_836 N_RESET_B_M1036_g N_VGND_c_2096_n 0.0013744f $X=3.5 $Y=0.615 $X2=0 $Y2=0
cc_837 N_RESET_B_c_891_n N_VGND_c_2096_n 0.0201841f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_838 N_RESET_B_c_891_n N_VGND_c_2097_n 0.0255051f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_839 N_RESET_B_M1014_g N_VGND_c_2098_n 0.0122528f $X=11.135 $Y=0.58 $X2=0
+ $Y2=0
cc_840 N_RESET_B_c_892_n N_VGND_c_2103_n 0.00710481f $X=3.575 $Y=0.18 $X2=0
+ $Y2=0
cc_841 N_RESET_B_c_891_n N_VGND_c_2105_n 0.0242408f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_842 N_RESET_B_c_891_n N_VGND_c_2108_n 0.0512939f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_843 N_RESET_B_M1014_g N_VGND_c_2110_n 0.00383152f $X=11.135 $Y=0.58 $X2=0
+ $Y2=0
cc_844 N_RESET_B_c_891_n N_VGND_c_2114_n 0.00939536f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_845 N_RESET_B_c_891_n N_VGND_c_2118_n 0.0912414f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_846 N_RESET_B_c_892_n N_VGND_c_2118_n 0.0112438f $X=3.575 $Y=0.18 $X2=0 $Y2=0
cc_847 N_RESET_B_M1014_g N_VGND_c_2118_n 0.0075694f $X=11.135 $Y=0.58 $X2=0
+ $Y2=0
cc_848 N_RESET_B_M1036_g N_noxref_24_c_2234_n 0.00427839f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_849 N_RESET_B_M1036_g N_noxref_24_c_2248_n 0.00289613f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_850 N_A_1234_119#_c_1121_n N_A_835_98#_c_1249_n 0.00321336f $X=6.685 $Y=2.555
+ $X2=0 $Y2=0
cc_851 N_A_1234_119#_c_1118_n N_A_835_98#_c_1238_n 0.00566398f $X=6.31 $Y=0.81
+ $X2=0 $Y2=0
cc_852 N_A_1234_119#_c_1121_n N_A_835_98#_M1008_g 0.0121868f $X=6.685 $Y=2.555
+ $X2=0 $Y2=0
cc_853 N_A_1234_119#_c_1123_n N_A_835_98#_M1008_g 0.00150864f $X=6.77 $Y=2.385
+ $X2=0 $Y2=0
cc_854 N_A_1234_119#_c_1111_n N_A_835_98#_c_1252_n 0.0103562f $X=8.64 $Y=1.66
+ $X2=0 $Y2=0
cc_855 N_A_1234_119#_c_1121_n N_A_835_98#_c_1252_n 0.00382216f $X=6.685 $Y=2.555
+ $X2=0 $Y2=0
cc_856 N_A_1234_119#_c_1127_n N_A_835_98#_c_1252_n 0.00592408f $X=7.62 $Y=2.53
+ $X2=0 $Y2=0
cc_857 N_A_1234_119#_c_1111_n N_A_835_98#_M1018_g 0.0199663f $X=8.64 $Y=1.66
+ $X2=0 $Y2=0
cc_858 N_A_1234_119#_c_1111_n N_A_835_98#_c_1255_n 0.00359436f $X=8.64 $Y=1.66
+ $X2=0 $Y2=0
cc_859 N_A_1234_119#_c_1111_n N_A_1824_74#_c_1558_n 4.59845e-19 $X=8.64 $Y=1.66
+ $X2=0 $Y2=0
cc_860 N_A_1234_119#_c_1121_n N_VPWR_c_1747_n 0.00162755f $X=6.685 $Y=2.555
+ $X2=0 $Y2=0
cc_861 N_A_1234_119#_c_1124_n N_VPWR_c_1747_n 0.0152964f $X=7.435 $Y=2.075 $X2=0
+ $Y2=0
cc_862 N_A_1234_119#_c_1127_n N_VPWR_c_1747_n 0.0165552f $X=7.62 $Y=2.53 $X2=0
+ $Y2=0
cc_863 N_A_1234_119#_c_1111_n N_VPWR_c_1748_n 0.0116888f $X=8.64 $Y=1.66 $X2=0
+ $Y2=0
cc_864 N_A_1234_119#_c_1127_n N_VPWR_c_1748_n 0.0162421f $X=7.62 $Y=2.53 $X2=0
+ $Y2=0
cc_865 N_A_1234_119#_c_1121_n N_VPWR_c_1755_n 0.0122075f $X=6.685 $Y=2.555 $X2=0
+ $Y2=0
cc_866 N_A_1234_119#_c_1127_n N_VPWR_c_1761_n 0.00718093f $X=7.62 $Y=2.53 $X2=0
+ $Y2=0
cc_867 N_A_1234_119#_c_1111_n N_VPWR_c_1744_n 8.51577e-19 $X=8.64 $Y=1.66 $X2=0
+ $Y2=0
cc_868 N_A_1234_119#_c_1121_n N_VPWR_c_1744_n 0.0157408f $X=6.685 $Y=2.555 $X2=0
+ $Y2=0
cc_869 N_A_1234_119#_c_1127_n N_VPWR_c_1744_n 0.00888445f $X=7.62 $Y=2.53 $X2=0
+ $Y2=0
cc_870 N_A_1234_119#_c_1118_n N_A_390_81#_c_1919_n 0.0168132f $X=6.31 $Y=0.81
+ $X2=0 $Y2=0
cc_871 N_A_1234_119#_c_1121_n N_A_390_81#_c_1927_n 0.0139433f $X=6.685 $Y=2.555
+ $X2=0 $Y2=0
cc_872 N_A_1234_119#_c_1123_n N_A_390_81#_c_1927_n 0.00314452f $X=6.77 $Y=2.385
+ $X2=0 $Y2=0
cc_873 N_A_1234_119#_c_1113_n N_A_390_81#_c_1920_n 0.00342789f $X=6.685 $Y=0.945
+ $X2=0 $Y2=0
cc_874 N_A_1234_119#_c_1114_n N_A_390_81#_c_1920_n 0.0136392f $X=6.77 $Y=1.985
+ $X2=0 $Y2=0
cc_875 N_A_1234_119#_c_1118_n N_A_390_81#_c_1920_n 0.0270482f $X=6.31 $Y=0.81
+ $X2=0 $Y2=0
cc_876 N_A_1234_119#_c_1121_n N_A_390_81#_c_1928_n 0.0180051f $X=6.685 $Y=2.555
+ $X2=0 $Y2=0
cc_877 N_A_1234_119#_c_1123_n N_A_390_81#_c_1928_n 0.00396213f $X=6.77 $Y=2.385
+ $X2=0 $Y2=0
cc_878 N_A_1234_119#_c_1126_n N_A_390_81#_c_1928_n 0.0100574f $X=6.77 $Y=2.075
+ $X2=0 $Y2=0
cc_879 N_A_1234_119#_c_1114_n N_A_390_81#_c_1922_n 0.0447672f $X=6.77 $Y=1.985
+ $X2=0 $Y2=0
cc_880 N_A_1234_119#_c_1126_n N_A_390_81#_c_1922_n 0.00431721f $X=6.77 $Y=2.075
+ $X2=0 $Y2=0
cc_881 N_A_1234_119#_M1035_g N_VGND_c_2109_n 0.00278271f $X=8.54 $Y=0.74 $X2=0
+ $Y2=0
cc_882 N_A_1234_119#_M1035_g N_VGND_c_2118_n 0.0035918f $X=8.54 $Y=0.74 $X2=0
+ $Y2=0
cc_883 N_A_1234_119#_c_1113_n A_1320_119# 0.00179335f $X=6.685 $Y=0.945
+ $X2=-0.19 $Y2=-0.245
cc_884 N_A_835_98#_c_1240_n N_A_2082_446#_M1003_g 0.00472321f $X=10.125 $Y=1.575
+ $X2=0 $Y2=0
cc_885 N_A_835_98#_M1002_g N_A_2082_446#_M1003_g 0.0465564f $X=10.315 $Y=0.58
+ $X2=0 $Y2=0
cc_886 N_A_835_98#_c_1239_n N_A_2082_446#_c_1417_n 0.00873113f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_887 N_A_835_98#_c_1240_n N_A_2082_446#_c_1424_n 0.00873113f $X=10.125
+ $Y=1.575 $X2=0 $Y2=0
cc_888 N_A_835_98#_M1018_g N_A_1824_74#_c_1563_n 0.00686632f $X=9.26 $Y=2.33
+ $X2=0 $Y2=0
cc_889 N_A_835_98#_c_1239_n N_A_1824_74#_c_1563_n 0.00627973f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_890 N_A_835_98#_M1002_g N_A_1824_74#_c_1545_n 0.0085841f $X=10.315 $Y=0.58
+ $X2=0 $Y2=0
cc_891 N_A_835_98#_c_1242_n N_A_1824_74#_c_1545_n 0.0073765f $X=10.315 $Y=1.055
+ $X2=0 $Y2=0
cc_892 N_A_835_98#_M1018_g N_A_1824_74#_c_1558_n 0.00525155f $X=9.26 $Y=2.33
+ $X2=0 $Y2=0
cc_893 N_A_835_98#_c_1257_n N_A_1824_74#_c_1558_n 4.63769e-19 $X=9.26 $Y=3.15
+ $X2=0 $Y2=0
cc_894 N_A_835_98#_M1002_g N_A_1824_74#_c_1546_n 0.00682018f $X=10.315 $Y=0.58
+ $X2=0 $Y2=0
cc_895 N_A_835_98#_c_1242_n N_A_1824_74#_c_1546_n 0.00308052f $X=10.315 $Y=1.055
+ $X2=0 $Y2=0
cc_896 N_A_835_98#_c_1240_n N_A_1824_74#_c_1547_n 0.00432791f $X=10.125 $Y=1.575
+ $X2=0 $Y2=0
cc_897 N_A_835_98#_c_1240_n N_A_1824_74#_c_1549_n 7.4004e-19 $X=10.125 $Y=1.575
+ $X2=0 $Y2=0
cc_898 N_A_835_98#_c_1242_n N_A_1824_74#_c_1549_n 0.00823777f $X=10.315 $Y=1.055
+ $X2=0 $Y2=0
cc_899 N_A_835_98#_c_1245_n N_VPWR_M1028_d 0.00264396f $X=4.93 $Y=1.852 $X2=0
+ $Y2=0
cc_900 N_A_835_98#_c_1247_n N_VPWR_c_1746_n 0.00850453f $X=5.095 $Y=1.875 $X2=0
+ $Y2=0
cc_901 N_A_835_98#_c_1248_n N_VPWR_c_1746_n 0.00158412f $X=5.615 $Y=3.075 $X2=0
+ $Y2=0
cc_902 N_A_835_98#_c_1250_n N_VPWR_c_1746_n 0.00232909f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_903 N_A_835_98#_M1008_g N_VPWR_c_1747_n 0.00714317f $X=6.585 $Y=2.495 $X2=0
+ $Y2=0
cc_904 N_A_835_98#_c_1252_n N_VPWR_c_1747_n 0.0210626f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_905 N_A_835_98#_c_1252_n N_VPWR_c_1748_n 0.0262303f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_906 N_A_835_98#_M1018_g N_VPWR_c_1748_n 0.00149025f $X=9.26 $Y=2.33 $X2=0
+ $Y2=0
cc_907 N_A_835_98#_c_1257_n N_VPWR_c_1748_n 0.00416255f $X=9.26 $Y=3.15 $X2=0
+ $Y2=0
cc_908 N_A_835_98#_c_1247_n N_VPWR_c_1755_n 0.00303678f $X=5.095 $Y=1.875 $X2=0
+ $Y2=0
cc_909 N_A_835_98#_c_1250_n N_VPWR_c_1755_n 0.0419935f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_910 N_A_835_98#_c_1252_n N_VPWR_c_1761_n 0.0308835f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_911 N_A_835_98#_c_1252_n N_VPWR_c_1762_n 0.0232816f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_912 N_A_835_98#_c_1247_n N_VPWR_c_1744_n 0.00394737f $X=5.095 $Y=1.875 $X2=0
+ $Y2=0
cc_913 N_A_835_98#_c_1249_n N_VPWR_c_1744_n 0.0241704f $X=6.51 $Y=3.15 $X2=0
+ $Y2=0
cc_914 N_A_835_98#_c_1250_n N_VPWR_c_1744_n 0.00688721f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_915 N_A_835_98#_c_1252_n N_VPWR_c_1744_n 0.0705408f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_916 N_A_835_98#_c_1256_n N_VPWR_c_1744_n 0.00423956f $X=6.585 $Y=3.15 $X2=0
+ $Y2=0
cc_917 N_A_835_98#_c_1257_n N_VPWR_c_1744_n 0.0122553f $X=9.26 $Y=3.15 $X2=0
+ $Y2=0
cc_918 N_A_835_98#_M1028_s N_A_390_81#_c_1924_n 0.00851724f $X=4.275 $Y=1.96
+ $X2=0 $Y2=0
cc_919 N_A_835_98#_c_1245_n N_A_390_81#_c_1924_n 0.017483f $X=4.93 $Y=1.852
+ $X2=0 $Y2=0
cc_920 N_A_835_98#_c_1247_n N_A_390_81#_c_1926_n 0.0151931f $X=5.095 $Y=1.875
+ $X2=0 $Y2=0
cc_921 N_A_835_98#_c_1248_n N_A_390_81#_c_1926_n 0.0148953f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_922 N_A_835_98#_c_1249_n N_A_390_81#_c_1926_n 7.24606e-19 $X=6.51 $Y=3.15
+ $X2=0 $Y2=0
cc_923 N_A_835_98#_c_1245_n N_A_390_81#_c_1926_n 0.0189376f $X=4.93 $Y=1.852
+ $X2=0 $Y2=0
cc_924 N_A_835_98#_c_1246_n N_A_390_81#_c_1926_n 4.98991e-19 $X=5.115 $Y=1.635
+ $X2=0 $Y2=0
cc_925 N_A_835_98#_c_1237_n N_A_390_81#_c_1919_n 0.00777044f $X=6.02 $Y=1.225
+ $X2=0 $Y2=0
cc_926 N_A_835_98#_c_1238_n N_A_390_81#_c_1919_n 0.00423903f $X=6.095 $Y=1.115
+ $X2=0 $Y2=0
cc_927 N_A_835_98#_c_1248_n N_A_390_81#_c_1927_n 0.00760865f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_928 N_A_835_98#_c_1249_n N_A_390_81#_c_1927_n 0.00469098f $X=6.51 $Y=3.15
+ $X2=0 $Y2=0
cc_929 N_A_835_98#_M1008_g N_A_390_81#_c_1927_n 5.52147e-19 $X=6.585 $Y=2.495
+ $X2=0 $Y2=0
cc_930 N_A_835_98#_c_1237_n N_A_390_81#_c_1920_n 0.0119917f $X=6.02 $Y=1.225
+ $X2=0 $Y2=0
cc_931 N_A_835_98#_c_1237_n N_A_390_81#_c_1921_n 0.00600188f $X=6.02 $Y=1.225
+ $X2=0 $Y2=0
cc_932 N_A_835_98#_c_1246_n N_A_390_81#_c_1921_n 7.71188e-19 $X=5.115 $Y=1.635
+ $X2=0 $Y2=0
cc_933 N_A_835_98#_M1008_g N_A_390_81#_c_1928_n 0.00138335f $X=6.585 $Y=2.495
+ $X2=0 $Y2=0
cc_934 N_A_835_98#_c_1248_n N_A_390_81#_c_1929_n 0.00126f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_935 N_A_835_98#_c_1246_n N_A_390_81#_c_1922_n 0.00436361f $X=5.115 $Y=1.635
+ $X2=0 $Y2=0
cc_936 N_A_835_98#_c_1243_n N_VGND_M1029_d 0.00428321f $X=4.93 $Y=1.455 $X2=0
+ $Y2=0
cc_937 N_A_835_98#_c_1244_n N_VGND_M1029_d 0.00811195f $X=4.32 $Y=0.665 $X2=0
+ $Y2=0
cc_938 N_A_835_98#_c_1244_n N_VGND_c_2096_n 0.0141187f $X=4.32 $Y=0.665 $X2=0
+ $Y2=0
cc_939 N_A_835_98#_c_1236_n N_VGND_c_2097_n 0.00191749f $X=5.145 $Y=1.41 $X2=0
+ $Y2=0
cc_940 N_A_835_98#_c_1244_n N_VGND_c_2097_n 0.0372149f $X=4.32 $Y=0.665 $X2=0
+ $Y2=0
cc_941 N_A_835_98#_c_1246_n N_VGND_c_2097_n 2.12055e-19 $X=5.115 $Y=1.635 $X2=0
+ $Y2=0
cc_942 N_A_835_98#_M1002_g N_VGND_c_2098_n 0.00155929f $X=10.315 $Y=0.58 $X2=0
+ $Y2=0
cc_943 N_A_835_98#_c_1244_n N_VGND_c_2105_n 0.0103545f $X=4.32 $Y=0.665 $X2=0
+ $Y2=0
cc_944 N_A_835_98#_M1002_g N_VGND_c_2109_n 0.00308264f $X=10.315 $Y=0.58 $X2=0
+ $Y2=0
cc_945 N_A_835_98#_c_1236_n N_VGND_c_2118_n 9.10391e-19 $X=5.145 $Y=1.41 $X2=0
+ $Y2=0
cc_946 N_A_835_98#_M1002_g N_VGND_c_2118_n 0.00383744f $X=10.315 $Y=0.58 $X2=0
+ $Y2=0
cc_947 N_A_835_98#_c_1244_n N_VGND_c_2118_n 0.0140767f $X=4.32 $Y=0.665 $X2=0
+ $Y2=0
cc_948 N_A_2082_446#_c_1419_n N_A_1824_74#_M1007_g 0.00761651f $X=11.71 $Y=0.58
+ $X2=0 $Y2=0
cc_949 N_A_2082_446#_c_1421_n N_A_1824_74#_M1007_g 0.00732912f $X=11.875
+ $Y=0.855 $X2=0 $Y2=0
cc_950 N_A_2082_446#_c_1422_n N_A_1824_74#_M1007_g 0.00376832f $X=12.145 $Y=1.58
+ $X2=0 $Y2=0
cc_951 N_A_2082_446#_c_1418_n N_A_1824_74#_c_1552_n 0.0116511f $X=12.06 $Y=1.665
+ $X2=0 $Y2=0
cc_952 N_A_2082_446#_c_1429_n N_A_1824_74#_c_1554_n 0.00502098f $X=11.41
+ $Y=2.475 $X2=0 $Y2=0
cc_953 N_A_2082_446#_c_1430_n N_A_1824_74#_c_1554_n 0.00496874f $X=11.575
+ $Y=2.75 $X2=0 $Y2=0
cc_954 N_A_2082_446#_c_1418_n N_A_1824_74#_c_1539_n 0.00220284f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_955 N_A_2082_446#_c_1422_n N_A_1824_74#_c_1539_n 0.022644f $X=12.145 $Y=1.58
+ $X2=0 $Y2=0
cc_956 N_A_2082_446#_c_1418_n N_A_1824_74#_c_1540_n 0.00461365f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_957 N_A_2082_446#_c_1420_n N_A_1824_74#_c_1540_n 0.0054249f $X=12.06 $Y=0.855
+ $X2=0 $Y2=0
cc_958 N_A_2082_446#_c_1421_n N_A_1824_74#_c_1540_n 0.00561111f $X=11.875
+ $Y=0.855 $X2=0 $Y2=0
cc_959 N_A_2082_446#_c_1418_n N_A_1824_74#_c_1541_n 0.00230014f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_960 N_A_2082_446#_c_1422_n N_A_1824_74#_c_1541_n 0.0017493f $X=12.145 $Y=1.58
+ $X2=0 $Y2=0
cc_961 N_A_2082_446#_c_1419_n N_A_1824_74#_c_1542_n 0.00350124f $X=11.71 $Y=0.58
+ $X2=0 $Y2=0
cc_962 N_A_2082_446#_c_1420_n N_A_1824_74#_c_1542_n 0.00386679f $X=12.06
+ $Y=0.855 $X2=0 $Y2=0
cc_963 N_A_2082_446#_c_1422_n N_A_1824_74#_c_1542_n 0.00324637f $X=12.145
+ $Y=1.58 $X2=0 $Y2=0
cc_964 N_A_2082_446#_c_1418_n N_A_1824_74#_c_1543_n 0.00573299f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_965 N_A_2082_446#_c_1422_n N_A_1824_74#_c_1543_n 0.00338011f $X=12.145
+ $Y=1.58 $X2=0 $Y2=0
cc_966 N_A_2082_446#_M1003_g N_A_1824_74#_c_1545_n 0.00114145f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_967 N_A_2082_446#_c_1425_n N_A_1824_74#_c_1557_n 0.00134164f $X=10.5 $Y=2.465
+ $X2=0 $Y2=0
cc_968 N_A_2082_446#_c_1486_p N_A_1824_74#_c_1557_n 0.00258251f $X=10.85
+ $Y=2.475 $X2=0 $Y2=0
cc_969 N_A_2082_446#_M1003_g N_A_1824_74#_c_1546_n 0.00142814f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_970 N_A_2082_446#_c_1425_n N_A_1824_74#_c_1547_n 3.62386e-19 $X=10.5 $Y=2.465
+ $X2=0 $Y2=0
cc_971 N_A_2082_446#_M1003_g N_A_1824_74#_c_1547_n 0.00172861f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_972 N_A_2082_446#_c_1426_n N_A_1824_74#_c_1547_n 0.00168467f $X=10.645
+ $Y=2.23 $X2=0 $Y2=0
cc_973 N_A_2082_446#_c_1486_p N_A_1824_74#_c_1547_n 0.0103077f $X=10.85 $Y=2.475
+ $X2=0 $Y2=0
cc_974 N_A_2082_446#_c_1423_n N_A_1824_74#_c_1547_n 0.074835f $X=10.685 $Y=1.535
+ $X2=0 $Y2=0
cc_975 N_A_2082_446#_c_1424_n N_A_1824_74#_c_1547_n 0.0114396f $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_976 N_A_2082_446#_c_1420_n N_A_1824_74#_c_1548_n 0.00108154f $X=12.06
+ $Y=0.855 $X2=0 $Y2=0
cc_977 N_A_2082_446#_c_1421_n N_A_1824_74#_c_1548_n 0.0272174f $X=11.875
+ $Y=0.855 $X2=0 $Y2=0
cc_978 N_A_2082_446#_c_1422_n N_A_1824_74#_c_1548_n 0.0227002f $X=12.145 $Y=1.58
+ $X2=0 $Y2=0
cc_979 N_A_2082_446#_M1003_g N_A_1824_74#_c_1550_n 0.0143673f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_980 N_A_2082_446#_c_1418_n N_A_1824_74#_c_1550_n 0.00732151f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_981 N_A_2082_446#_c_1423_n N_A_1824_74#_c_1550_n 0.0224547f $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_982 N_A_2082_446#_c_1424_n N_A_1824_74#_c_1550_n 0.00598209f $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_983 N_A_2082_446#_M1003_g N_A_1824_74#_c_1551_n 0.0019127f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_984 N_A_2082_446#_c_1418_n N_A_1824_74#_c_1551_n 0.06452f $X=12.06 $Y=1.665
+ $X2=0 $Y2=0
cc_985 N_A_2082_446#_c_1423_n N_A_1824_74#_c_1551_n 0.00326018f $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_986 N_A_2082_446#_c_1424_n N_A_1824_74#_c_1551_n 2.45278e-19 $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_987 N_A_2082_446#_c_1422_n N_A_2492_392#_c_1684_n 0.0135871f $X=12.145
+ $Y=1.58 $X2=0 $Y2=0
cc_988 N_A_2082_446#_c_1418_n N_A_2492_392#_c_1686_n 0.0058056f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_989 N_A_2082_446#_c_1418_n N_A_2492_392#_c_1687_n 0.00268745f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_990 N_A_2082_446#_c_1422_n N_A_2492_392#_c_1687_n 0.0131081f $X=12.145
+ $Y=1.58 $X2=0 $Y2=0
cc_991 N_A_2082_446#_c_1429_n N_VPWR_M1038_d 0.00387797f $X=11.41 $Y=2.475 $X2=0
+ $Y2=0
cc_992 N_A_2082_446#_c_1486_p N_VPWR_M1038_d 0.00236476f $X=10.85 $Y=2.475 $X2=0
+ $Y2=0
cc_993 N_A_2082_446#_c_1418_n N_VPWR_c_1749_n 0.0235807f $X=12.06 $Y=1.665 $X2=0
+ $Y2=0
cc_994 N_A_2082_446#_c_1429_n N_VPWR_c_1749_n 0.012314f $X=11.41 $Y=2.475 $X2=0
+ $Y2=0
cc_995 N_A_2082_446#_c_1430_n N_VPWR_c_1749_n 0.0282274f $X=11.575 $Y=2.75 $X2=0
+ $Y2=0
cc_996 N_A_2082_446#_c_1430_n N_VPWR_c_1757_n 0.0144033f $X=11.575 $Y=2.75 $X2=0
+ $Y2=0
cc_997 N_A_2082_446#_c_1425_n N_VPWR_c_1762_n 0.00415318f $X=10.5 $Y=2.465 $X2=0
+ $Y2=0
cc_998 N_A_2082_446#_c_1425_n N_VPWR_c_1768_n 0.00864935f $X=10.5 $Y=2.465 $X2=0
+ $Y2=0
cc_999 N_A_2082_446#_c_1426_n N_VPWR_c_1768_n 0.00123389f $X=10.645 $Y=2.23
+ $X2=0 $Y2=0
cc_1000 N_A_2082_446#_c_1429_n N_VPWR_c_1768_n 0.0288765f $X=11.41 $Y=2.475
+ $X2=0 $Y2=0
cc_1001 N_A_2082_446#_c_1486_p N_VPWR_c_1768_n 0.0201549f $X=10.85 $Y=2.475
+ $X2=0 $Y2=0
cc_1002 N_A_2082_446#_c_1430_n N_VPWR_c_1768_n 0.0102623f $X=11.575 $Y=2.75
+ $X2=0 $Y2=0
cc_1003 N_A_2082_446#_c_1425_n N_VPWR_c_1744_n 0.00817239f $X=10.5 $Y=2.465
+ $X2=0 $Y2=0
cc_1004 N_A_2082_446#_c_1426_n N_VPWR_c_1744_n 3.19707e-19 $X=10.645 $Y=2.23
+ $X2=0 $Y2=0
cc_1005 N_A_2082_446#_c_1429_n N_VPWR_c_1744_n 0.00667547f $X=11.41 $Y=2.475
+ $X2=0 $Y2=0
cc_1006 N_A_2082_446#_c_1486_p N_VPWR_c_1744_n 0.00116499f $X=10.85 $Y=2.475
+ $X2=0 $Y2=0
cc_1007 N_A_2082_446#_c_1430_n N_VPWR_c_1744_n 0.0119211f $X=11.575 $Y=2.75
+ $X2=0 $Y2=0
cc_1008 N_A_2082_446#_c_1420_n N_VGND_M1021_s 0.00405314f $X=12.06 $Y=0.855
+ $X2=0 $Y2=0
cc_1009 N_A_2082_446#_c_1422_n N_VGND_M1021_s 8.04296e-19 $X=12.145 $Y=1.58
+ $X2=0 $Y2=0
cc_1010 N_A_2082_446#_M1003_g N_VGND_c_2098_n 0.0119771f $X=10.705 $Y=0.58 $X2=0
+ $Y2=0
cc_1011 N_A_2082_446#_c_1419_n N_VGND_c_2098_n 0.0140354f $X=11.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1012 N_A_2082_446#_c_1421_n N_VGND_c_2098_n 0.00142029f $X=11.875 $Y=0.855
+ $X2=0 $Y2=0
cc_1013 N_A_2082_446#_c_1419_n N_VGND_c_2099_n 0.0168546f $X=11.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1014 N_A_2082_446#_c_1420_n N_VGND_c_2099_n 0.0109002f $X=12.06 $Y=0.855
+ $X2=0 $Y2=0
cc_1015 N_A_2082_446#_M1003_g N_VGND_c_2109_n 0.00383152f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_1016 N_A_2082_446#_c_1419_n N_VGND_c_2110_n 0.014415f $X=11.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1017 N_A_2082_446#_M1003_g N_VGND_c_2118_n 0.0075725f $X=10.705 $Y=0.58 $X2=0
+ $Y2=0
cc_1018 N_A_2082_446#_c_1419_n N_VGND_c_2118_n 0.0119404f $X=11.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1019 N_A_2082_446#_c_1420_n N_VGND_c_2118_n 0.0092009f $X=12.06 $Y=0.855
+ $X2=0 $Y2=0
cc_1020 N_A_1824_74#_c_1556_n N_A_2492_392#_c_1691_n 0.00352637f $X=12.385
+ $Y=1.885 $X2=0 $Y2=0
cc_1021 N_A_1824_74#_c_1544_n N_A_2492_392#_c_1691_n 0.00239754f $X=12.295
+ $Y=1.095 $X2=0 $Y2=0
cc_1022 N_A_1824_74#_c_1556_n N_A_2492_392#_c_1692_n 0.0089495f $X=12.385
+ $Y=1.885 $X2=0 $Y2=0
cc_1023 N_A_1824_74#_c_1542_n N_A_2492_392#_c_1684_n 0.00769864f $X=12.485
+ $Y=1.095 $X2=0 $Y2=0
cc_1024 N_A_1824_74#_c_1544_n N_A_2492_392#_c_1684_n 0.00167437f $X=12.295
+ $Y=1.095 $X2=0 $Y2=0
cc_1025 N_A_1824_74#_c_1541_n N_A_2492_392#_c_1686_n 0.00768781f $X=12.385
+ $Y=1.795 $X2=0 $Y2=0
cc_1026 N_A_1824_74#_c_1556_n N_A_2492_392#_c_1686_n 0.00189951f $X=12.385
+ $Y=1.885 $X2=0 $Y2=0
cc_1027 N_A_1824_74#_c_1544_n N_A_2492_392#_c_1687_n 0.00471821f $X=12.295
+ $Y=1.095 $X2=0 $Y2=0
cc_1028 N_A_1824_74#_c_1544_n N_A_2492_392#_c_1688_n 0.00503519f $X=12.295
+ $Y=1.095 $X2=0 $Y2=0
cc_1029 N_A_1824_74#_c_1553_n N_VPWR_c_1749_n 0.00975077f $X=11.8 $Y=2.375 $X2=0
+ $Y2=0
cc_1030 N_A_1824_74#_c_1554_n N_VPWR_c_1749_n 0.00807257f $X=11.8 $Y=2.465 $X2=0
+ $Y2=0
cc_1031 N_A_1824_74#_c_1539_n N_VPWR_c_1749_n 7.36409e-19 $X=12.295 $Y=1.26
+ $X2=0 $Y2=0
cc_1032 N_A_1824_74#_c_1556_n N_VPWR_c_1749_n 0.00991624f $X=12.385 $Y=1.885
+ $X2=0 $Y2=0
cc_1033 N_A_1824_74#_c_1556_n N_VPWR_c_1750_n 0.00456767f $X=12.385 $Y=1.885
+ $X2=0 $Y2=0
cc_1034 N_A_1824_74#_c_1554_n N_VPWR_c_1757_n 0.00445602f $X=11.8 $Y=2.465 $X2=0
+ $Y2=0
cc_1035 N_A_1824_74#_c_1557_n N_VPWR_c_1762_n 0.019583f $X=10.22 $Y=2.685 $X2=0
+ $Y2=0
cc_1036 N_A_1824_74#_c_1558_n N_VPWR_c_1762_n 0.00812764f $X=9.6 $Y=2.685 $X2=0
+ $Y2=0
cc_1037 N_A_1824_74#_c_1556_n N_VPWR_c_1763_n 0.00445602f $X=12.385 $Y=1.885
+ $X2=0 $Y2=0
cc_1038 N_A_1824_74#_c_1554_n N_VPWR_c_1744_n 0.00896763f $X=11.8 $Y=2.465 $X2=0
+ $Y2=0
cc_1039 N_A_1824_74#_c_1556_n N_VPWR_c_1744_n 0.00862869f $X=12.385 $Y=1.885
+ $X2=0 $Y2=0
cc_1040 N_A_1824_74#_c_1557_n N_VPWR_c_1744_n 0.025422f $X=10.22 $Y=2.685 $X2=0
+ $Y2=0
cc_1041 N_A_1824_74#_c_1558_n N_VPWR_c_1744_n 0.00936382f $X=9.6 $Y=2.685 $X2=0
+ $Y2=0
cc_1042 N_A_1824_74#_c_1557_n A_2037_508# 0.00191616f $X=10.22 $Y=2.685
+ $X2=-0.19 $Y2=-0.245
cc_1043 N_A_1824_74#_M1007_g N_VGND_c_2098_n 0.00182082f $X=11.495 $Y=0.58 $X2=0
+ $Y2=0
cc_1044 N_A_1824_74#_c_1545_n N_VGND_c_2098_n 0.014224f $X=10.22 $Y=0.645 $X2=0
+ $Y2=0
cc_1045 N_A_1824_74#_c_1550_n N_VGND_c_2098_n 0.0229174f $X=11.02 $Y=1.22 $X2=0
+ $Y2=0
cc_1046 N_A_1824_74#_M1007_g N_VGND_c_2099_n 0.00324482f $X=11.495 $Y=0.58 $X2=0
+ $Y2=0
cc_1047 N_A_1824_74#_c_1539_n N_VGND_c_2099_n 0.00356476f $X=12.295 $Y=1.26
+ $X2=0 $Y2=0
cc_1048 N_A_1824_74#_c_1542_n N_VGND_c_2099_n 0.00936719f $X=12.485 $Y=1.095
+ $X2=0 $Y2=0
cc_1049 N_A_1824_74#_c_1542_n N_VGND_c_2100_n 0.00296233f $X=12.485 $Y=1.095
+ $X2=0 $Y2=0
cc_1050 N_A_1824_74#_c_1545_n N_VGND_c_2109_n 0.0249458f $X=10.22 $Y=0.645 $X2=0
+ $Y2=0
cc_1051 N_A_1824_74#_M1007_g N_VGND_c_2110_n 0.00434272f $X=11.495 $Y=0.58 $X2=0
+ $Y2=0
cc_1052 N_A_1824_74#_c_1542_n N_VGND_c_2111_n 0.00383152f $X=12.485 $Y=1.095
+ $X2=0 $Y2=0
cc_1053 N_A_1824_74#_M1007_g N_VGND_c_2118_n 0.00825669f $X=11.495 $Y=0.58 $X2=0
+ $Y2=0
cc_1054 N_A_1824_74#_c_1542_n N_VGND_c_2118_n 0.00762539f $X=12.485 $Y=1.095
+ $X2=0 $Y2=0
cc_1055 N_A_1824_74#_c_1545_n N_VGND_c_2118_n 0.0310203f $X=10.22 $Y=0.645 $X2=0
+ $Y2=0
cc_1056 N_A_2492_392#_c_1691_n N_VPWR_c_1749_n 0.0405667f $X=12.61 $Y=2.105
+ $X2=0 $Y2=0
cc_1057 N_A_2492_392#_c_1689_n N_VPWR_c_1750_n 0.0180379f $X=13.395 $Y=1.765
+ $X2=0 $Y2=0
cc_1058 N_A_2492_392#_c_1690_n N_VPWR_c_1750_n 7.0907e-19 $X=13.845 $Y=1.765
+ $X2=0 $Y2=0
cc_1059 N_A_2492_392#_c_1685_n N_VPWR_c_1750_n 0.025458f $X=13.19 $Y=1.465 $X2=0
+ $Y2=0
cc_1060 N_A_2492_392#_c_1686_n N_VPWR_c_1750_n 0.0777543f $X=12.61 $Y=1.94 $X2=0
+ $Y2=0
cc_1061 N_A_2492_392#_c_1688_n N_VPWR_c_1750_n 0.00689404f $X=13.845 $Y=1.532
+ $X2=0 $Y2=0
cc_1062 N_A_2492_392#_c_1690_n N_VPWR_c_1752_n 0.0260843f $X=13.845 $Y=1.765
+ $X2=0 $Y2=0
cc_1063 N_A_2492_392#_c_1688_n N_VPWR_c_1752_n 9.39066e-19 $X=13.845 $Y=1.532
+ $X2=0 $Y2=0
cc_1064 N_A_2492_392#_c_1692_n N_VPWR_c_1763_n 0.0145938f $X=12.61 $Y=2.815
+ $X2=0 $Y2=0
cc_1065 N_A_2492_392#_c_1689_n N_VPWR_c_1764_n 0.00413917f $X=13.395 $Y=1.765
+ $X2=0 $Y2=0
cc_1066 N_A_2492_392#_c_1690_n N_VPWR_c_1764_n 0.00445602f $X=13.845 $Y=1.765
+ $X2=0 $Y2=0
cc_1067 N_A_2492_392#_c_1689_n N_VPWR_c_1744_n 0.00817726f $X=13.395 $Y=1.765
+ $X2=0 $Y2=0
cc_1068 N_A_2492_392#_c_1690_n N_VPWR_c_1744_n 0.00860566f $X=13.845 $Y=1.765
+ $X2=0 $Y2=0
cc_1069 N_A_2492_392#_c_1692_n N_VPWR_c_1744_n 0.0120466f $X=12.61 $Y=2.815
+ $X2=0 $Y2=0
cc_1070 N_A_2492_392#_c_1689_n N_Q_c_2074_n 0.00196498f $X=13.395 $Y=1.765 $X2=0
+ $Y2=0
cc_1071 N_A_2492_392#_c_1690_n N_Q_c_2074_n 0.0153501f $X=13.845 $Y=1.765 $X2=0
+ $Y2=0
cc_1072 N_A_2492_392#_c_1688_n N_Q_c_2074_n 0.0338785f $X=13.845 $Y=1.532 $X2=0
+ $Y2=0
cc_1073 N_A_2492_392#_M1023_g Q 0.0138248f $X=13.475 $Y=0.74 $X2=0 $Y2=0
cc_1074 N_A_2492_392#_M1041_g Q 0.0162403f $X=13.905 $Y=0.74 $X2=0 $Y2=0
cc_1075 N_A_2492_392#_c_1684_n Q 0.00465944f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1076 N_A_2492_392#_M1023_g Q 0.0018463f $X=13.475 $Y=0.74 $X2=0 $Y2=0
cc_1077 N_A_2492_392#_M1041_g Q 0.00299044f $X=13.905 $Y=0.74 $X2=0 $Y2=0
cc_1078 N_A_2492_392#_c_1685_n Q 0.02585f $X=13.19 $Y=1.465 $X2=0 $Y2=0
cc_1079 N_A_2492_392#_c_1688_n Q 0.015501f $X=13.845 $Y=1.532 $X2=0 $Y2=0
cc_1080 N_A_2492_392#_c_1684_n N_VGND_c_2099_n 0.0101431f $X=12.7 $Y=0.515 $X2=0
+ $Y2=0
cc_1081 N_A_2492_392#_M1023_g N_VGND_c_2100_n 0.00647412f $X=13.475 $Y=0.74
+ $X2=0 $Y2=0
cc_1082 N_A_2492_392#_c_1684_n N_VGND_c_2100_n 0.0505719f $X=12.7 $Y=0.515 $X2=0
+ $Y2=0
cc_1083 N_A_2492_392#_c_1685_n N_VGND_c_2100_n 0.0209147f $X=13.19 $Y=1.465
+ $X2=0 $Y2=0
cc_1084 N_A_2492_392#_c_1688_n N_VGND_c_2100_n 0.0058967f $X=13.845 $Y=1.532
+ $X2=0 $Y2=0
cc_1085 N_A_2492_392#_M1041_g N_VGND_c_2102_n 0.00647412f $X=13.905 $Y=0.74
+ $X2=0 $Y2=0
cc_1086 N_A_2492_392#_c_1684_n N_VGND_c_2111_n 0.0115122f $X=12.7 $Y=0.515 $X2=0
+ $Y2=0
cc_1087 N_A_2492_392#_M1023_g N_VGND_c_2112_n 0.00434272f $X=13.475 $Y=0.74
+ $X2=0 $Y2=0
cc_1088 N_A_2492_392#_M1041_g N_VGND_c_2112_n 0.00434272f $X=13.905 $Y=0.74
+ $X2=0 $Y2=0
cc_1089 N_A_2492_392#_M1023_g N_VGND_c_2118_n 0.00825283f $X=13.475 $Y=0.74
+ $X2=0 $Y2=0
cc_1090 N_A_2492_392#_M1041_g N_VGND_c_2118_n 0.00823942f $X=13.905 $Y=0.74
+ $X2=0 $Y2=0
cc_1091 N_A_2492_392#_c_1684_n N_VGND_c_2118_n 0.0095288f $X=12.7 $Y=0.515 $X2=0
+ $Y2=0
cc_1092 N_VPWR_M1027_d N_A_390_81#_c_1932_n 0.0103722f $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1093 N_VPWR_c_1745_n N_A_390_81#_c_1932_n 0.0214041f $X=3.26 $Y=2.815 $X2=0
+ $Y2=0
cc_1094 N_VPWR_c_1744_n N_A_390_81#_c_1932_n 0.0235488f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1095 N_VPWR_c_1753_n N_A_390_81#_c_1924_n 0.00543175f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1096 N_VPWR_c_1744_n N_A_390_81#_c_1924_n 0.0102994f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1097 N_VPWR_M1027_d N_A_390_81#_c_1925_n 8.43866e-19 $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1098 N_VPWR_c_1745_n N_A_390_81#_c_1925_n 0.0213647f $X=3.26 $Y=2.815 $X2=0
+ $Y2=0
cc_1099 N_VPWR_c_1753_n N_A_390_81#_c_1925_n 0.0207455f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1100 N_VPWR_c_1744_n N_A_390_81#_c_1925_n 0.0268061f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1101 N_VPWR_M1028_d N_A_390_81#_c_1926_n 0.00387164f $X=4.72 $Y=1.96 $X2=0
+ $Y2=0
cc_1102 N_VPWR_c_1746_n N_A_390_81#_c_1926_n 0.0167709f $X=4.87 $Y=2.835 $X2=0
+ $Y2=0
cc_1103 N_VPWR_c_1753_n N_A_390_81#_c_1926_n 7.54393e-19 $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1104 N_VPWR_c_1755_n N_A_390_81#_c_1926_n 0.0103722f $X=7.025 $Y=3.33 $X2=0
+ $Y2=0
cc_1105 N_VPWR_c_1744_n N_A_390_81#_c_1926_n 0.0213354f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1106 N_VPWR_c_1755_n N_A_390_81#_c_1927_n 0.00535093f $X=7.025 $Y=3.33 $X2=0
+ $Y2=0
cc_1107 N_VPWR_c_1744_n N_A_390_81#_c_1927_n 0.00675054f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1108 N_VPWR_c_1745_n N_A_390_81#_c_1931_n 0.00703114f $X=3.26 $Y=2.815 $X2=0
+ $Y2=0
cc_1109 N_VPWR_c_1760_n N_A_390_81#_c_1931_n 0.0144502f $X=3.095 $Y=3.33 $X2=0
+ $Y2=0
cc_1110 N_VPWR_c_1765_n N_A_390_81#_c_1931_n 0.0201674f $X=1.4 $Y=2.465 $X2=0
+ $Y2=0
cc_1111 N_VPWR_c_1744_n N_A_390_81#_c_1931_n 0.0119027f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1112 N_VPWR_c_1750_n N_Q_c_2074_n 0.0412253f $X=13.17 $Y=1.985 $X2=0 $Y2=0
cc_1113 N_VPWR_c_1752_n N_Q_c_2074_n 0.0435456f $X=14.12 $Y=1.985 $X2=0 $Y2=0
cc_1114 N_VPWR_c_1764_n N_Q_c_2074_n 0.0114703f $X=13.955 $Y=3.33 $X2=0 $Y2=0
cc_1115 N_VPWR_c_1744_n N_Q_c_2074_n 0.00946127f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1116 N_A_390_81#_c_1932_n A_512_464# 0.0136022f $X=3.445 $Y=2.43 $X2=-0.19
+ $Y2=-0.245
cc_1117 N_A_390_81#_M1006_d N_noxref_24_c_2234_n 0.00972395f $X=1.95 $Y=0.405
+ $X2=0 $Y2=0
cc_1118 N_A_390_81#_c_1916_n N_noxref_24_c_2234_n 0.0449825f $X=2.785 $Y=0.72
+ $X2=0 $Y2=0
cc_1119 N_A_390_81#_c_1916_n N_noxref_24_c_2248_n 0.0287162f $X=2.785 $Y=0.72
+ $X2=0 $Y2=0
cc_1120 N_A_390_81#_c_1916_n noxref_26 0.00127671f $X=2.785 $Y=0.72 $X2=-0.19
+ $Y2=-0.245
cc_1121 Q N_VGND_c_2100_n 0.0294122f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1122 Q N_VGND_c_2102_n 0.0294122f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1123 Q N_VGND_c_2112_n 0.0144922f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1124 Q N_VGND_c_2118_n 0.0118826f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1125 N_VGND_c_2096_n N_noxref_24_c_2234_n 0.0125993f $X=3.76 $Y=0.565 $X2=0
+ $Y2=0
cc_1126 N_VGND_c_2103_n N_noxref_24_c_2234_n 0.12976f $X=3.61 $Y=0 $X2=0 $Y2=0
cc_1127 N_VGND_c_2118_n N_noxref_24_c_2234_n 0.0752032f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1128 N_VGND_c_2095_n N_noxref_24_c_2235_n 0.0259561f $X=0.71 $Y=0.555 $X2=0
+ $Y2=0
cc_1129 N_VGND_c_2103_n N_noxref_24_c_2235_n 0.0225398f $X=3.61 $Y=0 $X2=0 $Y2=0
cc_1130 N_VGND_c_2118_n N_noxref_24_c_2235_n 0.0125704f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1131 N_noxref_24_c_2234_n noxref_25 0.0013394f $X=3.19 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1132 N_noxref_24_c_2234_n noxref_26 0.00130751f $X=3.19 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
