* File: sky130_fd_sc_ls__inv_8.pxi.spice
* Created: Fri Aug 28 13:28:49 2020
* 
x_PM_SKY130_FD_SC_LS__INV_8%A N_A_c_77_n N_A_M1000_g N_A_c_68_n N_A_M1001_g
+ N_A_c_69_n N_A_M1004_g N_A_c_78_n N_A_M1002_g N_A_M1005_g N_A_c_79_n
+ N_A_M1003_g N_A_M1009_g N_A_c_80_n N_A_M1006_g N_A_M1011_g N_A_c_81_n
+ N_A_M1007_g N_A_M1013_g N_A_c_82_n N_A_M1008_g N_A_M1014_g N_A_c_83_n
+ N_A_M1010_g N_A_c_75_n N_A_M1015_g N_A_c_85_n N_A_M1012_g A A A N_A_c_86_n
+ PM_SKY130_FD_SC_LS__INV_8%A
x_PM_SKY130_FD_SC_LS__INV_8%VPWR N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_M1006_d
+ N_VPWR_M1008_d N_VPWR_M1012_d N_VPWR_c_213_n N_VPWR_c_214_n N_VPWR_c_215_n
+ N_VPWR_c_216_n N_VPWR_c_217_n N_VPWR_c_218_n N_VPWR_c_219_n N_VPWR_c_220_n
+ N_VPWR_c_221_n VPWR N_VPWR_c_222_n N_VPWR_c_223_n N_VPWR_c_224_n
+ N_VPWR_c_225_n N_VPWR_c_226_n N_VPWR_c_212_n PM_SKY130_FD_SC_LS__INV_8%VPWR
x_PM_SKY130_FD_SC_LS__INV_8%Y N_Y_M1001_s N_Y_M1005_s N_Y_M1011_s N_Y_M1014_s
+ N_Y_M1000_s N_Y_M1003_s N_Y_M1007_s N_Y_M1010_s N_Y_c_281_n N_Y_c_300_n
+ N_Y_c_293_n N_Y_c_282_n N_Y_c_283_n N_Y_c_312_n N_Y_c_284_n N_Y_c_294_n
+ N_Y_c_285_n N_Y_c_326_n N_Y_c_286_n N_Y_c_295_n N_Y_c_296_n N_Y_c_287_n
+ N_Y_c_288_n N_Y_c_297_n N_Y_c_289_n N_Y_c_352_n N_Y_c_290_n N_Y_c_389_n
+ N_Y_c_291_n Y PM_SKY130_FD_SC_LS__INV_8%Y
x_PM_SKY130_FD_SC_LS__INV_8%VGND N_VGND_M1001_d N_VGND_M1004_d N_VGND_M1009_d
+ N_VGND_M1013_d N_VGND_M1015_d N_VGND_c_414_n N_VGND_c_415_n N_VGND_c_416_n
+ N_VGND_c_417_n N_VGND_c_418_n N_VGND_c_419_n N_VGND_c_420_n N_VGND_c_421_n
+ N_VGND_c_422_n N_VGND_c_423_n N_VGND_c_424_n VGND N_VGND_c_425_n
+ N_VGND_c_426_n N_VGND_c_427_n N_VGND_c_428_n PM_SKY130_FD_SC_LS__INV_8%VGND
cc_1 VNB N_A_c_68_n 0.0184811f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.2
cc_2 VNB N_A_c_69_n 0.0148647f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.2
cc_3 VNB N_A_M1005_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=0.74
cc_4 VNB N_A_M1009_g 0.0234581f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=0.74
cc_5 VNB N_A_M1011_g 0.0239956f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=0.74
cc_6 VNB N_A_M1013_g 0.0235862f $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=0.74
cc_7 VNB N_A_M1014_g 0.02357f $X=-0.19 $Y=-0.245 $X2=3.3 $Y2=0.74
cc_8 VNB N_A_c_75_n 0.18624f $X=-0.19 $Y=-0.245 $X2=3.73 $Y2=1.35
cc_9 VNB N_A_M1015_g 0.0274509f $X=-0.19 $Y=-0.245 $X2=3.73 $Y2=0.74
cc_10 VNB N_VPWR_c_212_n 0.183584f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=1.482
cc_11 VNB N_Y_c_281_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.35
cc_12 VNB N_Y_c_282_n 0.00324651f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=2.4
cc_13 VNB N_Y_c_283_n 0.00176308f $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=1.35
cc_14 VNB N_Y_c_284_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=2.4
cc_15 VNB N_Y_c_285_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=3.305 $Y2=1.765
cc_16 VNB N_Y_c_286_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_287_n 0.00671548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_288_n 0.00241914f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.482
cc_19 VNB N_Y_c_289_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=1.515
cc_20 VNB N_Y_c_290_n 0.00458554f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=1.482
cc_21 VNB N_Y_c_291_n 0.00183274f $X=-0.19 $Y=-0.245 $X2=3.305 $Y2=1.482
cc_22 VNB Y 0.0327695f $X=-0.19 $Y=-0.245 $X2=3.73 $Y2=1.482
cc_23 VNB N_VGND_c_414_n 0.0111565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_415_n 0.0498215f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_25 VNB N_VGND_c_416_n 0.0026136f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=0.74
cc_26 VNB N_VGND_c_417_n 0.00498656f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=2.4
cc_27 VNB N_VGND_c_418_n 0.00817312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_419_n 0.0150576f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=2.4
cc_29 VNB N_VGND_c_420_n 0.0321594f $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=1.35
cc_30 VNB N_VGND_c_421_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_422_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=1.765
cc_32 VNB N_VGND_c_423_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=2.4
cc_33 VNB N_VGND_c_424_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=3.3 $Y2=1.35
cc_34 VNB N_VGND_c_425_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_426_n 0.0168561f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_36 VNB N_VGND_c_427_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.515
cc_37 VNB N_VGND_c_428_n 0.256334f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=1.482
cc_38 VPB N_A_c_77_n 0.0177026f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_39 VPB N_A_c_78_n 0.0153817f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_40 VPB N_A_c_79_n 0.0158901f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_41 VPB N_A_c_80_n 0.0155091f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.765
cc_42 VPB N_A_c_81_n 0.0150742f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=1.765
cc_43 VPB N_A_c_82_n 0.0153553f $X=-0.19 $Y=1.66 $X2=2.805 $Y2=1.765
cc_44 VPB N_A_c_83_n 0.0156611f $X=-0.19 $Y=1.66 $X2=3.305 $Y2=1.765
cc_45 VPB N_A_c_75_n 0.113901f $X=-0.19 $Y=1.66 $X2=3.73 $Y2=1.35
cc_46 VPB N_A_c_85_n 0.0174155f $X=-0.19 $Y=1.66 $X2=3.755 $Y2=1.765
cc_47 VPB N_A_c_86_n 0.0120353f $X=-0.19 $Y=1.66 $X2=2.085 $Y2=1.515
cc_48 VPB N_VPWR_c_213_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_214_n 0.0639451f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_50 VPB N_VPWR_c_215_n 0.00594454f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.765
cc_51 VPB N_VPWR_c_216_n 0.00504372f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=0.74
cc_52 VPB N_VPWR_c_217_n 0.00734988f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=2.4
cc_53 VPB N_VPWR_c_218_n 0.0125099f $X=-0.19 $Y=1.66 $X2=2.73 $Y2=0.74
cc_54 VPB N_VPWR_c_219_n 0.0594616f $X=-0.19 $Y=1.66 $X2=2.805 $Y2=1.765
cc_55 VPB N_VPWR_c_220_n 0.0164465f $X=-0.19 $Y=1.66 $X2=3.3 $Y2=0.74
cc_56 VPB N_VPWR_c_221_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_222_n 0.0185253f $X=-0.19 $Y=1.66 $X2=3.305 $Y2=2.4
cc_58 VPB N_VPWR_c_223_n 0.0196495f $X=-0.19 $Y=1.66 $X2=3.755 $Y2=1.765
cc_59 VPB N_VPWR_c_224_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.482
cc_60 VPB N_VPWR_c_225_n 0.00614127f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.482
cc_61 VPB N_VPWR_c_226_n 0.00460249f $X=-0.19 $Y=1.66 $X2=2.085 $Y2=1.482
cc_62 VPB N_VPWR_c_212_n 0.0704964f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=1.482
cc_63 VPB N_Y_c_293_n 0.00216998f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=1.765
cc_64 VPB N_Y_c_294_n 0.00257348f $X=-0.19 $Y=1.66 $X2=3.3 $Y2=0.74
cc_65 VPB N_Y_c_295_n 0.00259215f $X=-0.19 $Y=1.66 $X2=3.755 $Y2=2.4
cc_66 VPB N_Y_c_296_n 0.00180921f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_67 VPB N_Y_c_297_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.482
cc_68 N_A_c_77_n N_VPWR_c_214_n 0.0110944f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_69 N_A_c_77_n N_VPWR_c_215_n 5.55114e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_70 N_A_c_78_n N_VPWR_c_215_n 0.0110935f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_71 N_A_c_79_n N_VPWR_c_215_n 0.0068696f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_72 N_A_c_80_n N_VPWR_c_216_n 0.00526215f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A_c_81_n N_VPWR_c_216_n 0.0106464f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_74 N_A_c_82_n N_VPWR_c_216_n 5.37805e-19 $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_75 N_A_c_81_n N_VPWR_c_217_n 5.87963e-19 $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A_c_82_n N_VPWR_c_217_n 0.0165883f $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_77 N_A_c_83_n N_VPWR_c_217_n 0.00804662f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_78 N_A_c_75_n N_VPWR_c_217_n 0.00809737f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_79 N_A_c_85_n N_VPWR_c_219_n 0.0261486f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A_c_81_n N_VPWR_c_220_n 0.00413917f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A_c_82_n N_VPWR_c_220_n 0.00413917f $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_c_77_n N_VPWR_c_222_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_83 N_A_c_78_n N_VPWR_c_222_n 0.00413917f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_84 N_A_c_79_n N_VPWR_c_223_n 0.00445602f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A_c_80_n N_VPWR_c_223_n 0.00445602f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A_c_83_n N_VPWR_c_224_n 0.00445602f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_87 N_A_c_85_n N_VPWR_c_224_n 0.00445602f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A_c_77_n N_VPWR_c_212_n 0.00861084f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A_c_78_n N_VPWR_c_212_n 0.00817726f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A_c_79_n N_VPWR_c_212_n 0.00857378f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A_c_80_n N_VPWR_c_212_n 0.00857589f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A_c_81_n N_VPWR_c_212_n 0.00817726f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A_c_82_n N_VPWR_c_212_n 0.00817726f $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A_c_83_n N_VPWR_c_212_n 0.00857378f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A_c_85_n N_VPWR_c_212_n 0.00860594f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A_c_68_n N_Y_c_281_n 0.00814975f $X=0.51 $Y=1.2 $X2=0 $Y2=0
cc_97 N_A_c_69_n N_Y_c_281_n 3.97481e-19 $X=0.94 $Y=1.2 $X2=0 $Y2=0
cc_98 N_A_c_77_n N_Y_c_300_n 0.00203651f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_c_75_n N_Y_c_300_n 0.00123888f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_100 N_A_c_86_n N_Y_c_300_n 0.0193936f $X=2.085 $Y=1.515 $X2=0 $Y2=0
cc_101 N_A_c_77_n N_Y_c_293_n 0.00955225f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_c_78_n N_Y_c_293_n 0.00605728f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A_c_69_n N_Y_c_282_n 0.0130918f $X=0.94 $Y=1.2 $X2=0 $Y2=0
cc_104 N_A_M1005_g N_Y_c_282_n 0.0130918f $X=1.37 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_c_75_n N_Y_c_282_n 0.00224206f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_106 N_A_c_86_n N_Y_c_282_n 0.0517342f $X=2.085 $Y=1.515 $X2=0 $Y2=0
cc_107 N_A_c_68_n N_Y_c_283_n 0.00486135f $X=0.51 $Y=1.2 $X2=0 $Y2=0
cc_108 N_A_c_75_n N_Y_c_283_n 0.00301484f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_109 N_A_c_86_n N_Y_c_283_n 0.0213612f $X=2.085 $Y=1.515 $X2=0 $Y2=0
cc_110 N_A_c_78_n N_Y_c_312_n 0.0129585f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A_c_79_n N_Y_c_312_n 0.0122806f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_112 N_A_c_75_n N_Y_c_312_n 0.00176917f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_113 N_A_c_86_n N_Y_c_312_n 0.0475354f $X=2.085 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A_M1005_g N_Y_c_284_n 3.92313e-19 $X=1.37 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A_M1009_g N_Y_c_284_n 3.92313e-19 $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A_c_78_n N_Y_c_294_n 8.85795e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A_c_79_n N_Y_c_294_n 0.0100941f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_118 N_A_c_80_n N_Y_c_294_n 0.0105452f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A_c_81_n N_Y_c_294_n 6.69308e-19 $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A_M1009_g N_Y_c_285_n 0.0134851f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A_M1011_g N_Y_c_285_n 0.0145021f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A_c_75_n N_Y_c_285_n 0.00388688f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_123 N_A_c_86_n N_Y_c_285_n 0.0438012f $X=2.085 $Y=1.515 $X2=0 $Y2=0
cc_124 N_A_c_80_n N_Y_c_326_n 0.0119563f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A_c_81_n N_Y_c_326_n 0.0170871f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A_c_75_n N_Y_c_326_n 0.00227731f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_127 N_A_c_86_n N_Y_c_326_n 0.0282713f $X=2.085 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A_M1009_g N_Y_c_286_n 9.06576e-19 $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A_M1011_g N_Y_c_286_n 0.00945641f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_M1013_g N_Y_c_286_n 0.00837625f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A_M1014_g N_Y_c_286_n 2.47834e-19 $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A_c_81_n N_Y_c_295_n 0.00368201f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A_c_82_n N_Y_c_295_n 0.00180034f $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A_c_75_n N_Y_c_295_n 0.0114492f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_135 N_A_c_86_n N_Y_c_295_n 0.00984427f $X=2.085 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A_c_81_n N_Y_c_296_n 0.0039133f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A_c_82_n N_Y_c_296_n 0.00301623f $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A_M1013_g N_Y_c_287_n 0.011986f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_M1014_g N_Y_c_287_n 0.011986f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A_c_75_n N_Y_c_287_n 0.0402923f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_141 N_A_M1013_g N_Y_c_288_n 6.56051e-19 $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A_M1014_g N_Y_c_288_n 0.0110703f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A_M1015_g N_Y_c_288_n 0.00114583f $X=3.73 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A_c_82_n N_Y_c_297_n 5.5832e-19 $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A_c_83_n N_Y_c_297_n 0.0140077f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A_c_75_n N_Y_c_297_n 0.022394f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_147 N_A_c_85_n N_Y_c_297_n 0.015803f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A_c_75_n N_Y_c_289_n 0.00234043f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_149 N_A_c_86_n N_Y_c_289_n 0.0146029f $X=2.085 $Y=1.515 $X2=0 $Y2=0
cc_150 N_A_c_79_n N_Y_c_352_n 4.27055e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A_c_80_n N_Y_c_352_n 4.27055e-19 $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A_c_75_n N_Y_c_352_n 0.00144091f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_153 N_A_c_86_n N_Y_c_352_n 0.0237598f $X=2.085 $Y=1.515 $X2=0 $Y2=0
cc_154 N_A_M1011_g N_Y_c_290_n 0.0078432f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_M1013_g N_Y_c_290_n 0.00547674f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_M1014_g N_Y_c_290_n 4.05789e-19 $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A_c_75_n N_Y_c_290_n 0.0128858f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_158 N_A_c_86_n N_Y_c_290_n 0.0169547f $X=2.085 $Y=1.515 $X2=0 $Y2=0
cc_159 N_A_M1014_g N_Y_c_291_n 0.00298831f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_c_75_n N_Y_c_291_n 0.0120112f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_161 N_A_M1015_g N_Y_c_291_n 0.00536013f $X=3.73 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A_c_75_n Y 0.0174567f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_163 N_A_M1015_g Y 0.0111608f $X=3.73 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A_c_68_n N_VGND_c_415_n 0.00511131f $X=0.51 $Y=1.2 $X2=0 $Y2=0
cc_165 N_A_c_68_n N_VGND_c_416_n 5.19194e-19 $X=0.51 $Y=1.2 $X2=0 $Y2=0
cc_166 N_A_c_69_n N_VGND_c_416_n 0.0108127f $X=0.94 $Y=1.2 $X2=0 $Y2=0
cc_167 N_A_M1005_g N_VGND_c_416_n 0.0106755f $X=1.37 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A_M1009_g N_VGND_c_416_n 4.71636e-19 $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A_M1005_g N_VGND_c_417_n 4.71636e-19 $X=1.37 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A_M1009_g N_VGND_c_417_n 0.0106899f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A_M1011_g N_VGND_c_417_n 0.00432843f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A_M1013_g N_VGND_c_418_n 0.00563364f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A_M1014_g N_VGND_c_418_n 0.0055442f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A_c_75_n N_VGND_c_418_n 0.00117726f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_175 N_A_M1014_g N_VGND_c_420_n 5.47e-19 $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_M1015_g N_VGND_c_420_n 0.0117247f $X=3.73 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A_M1005_g N_VGND_c_421_n 0.00383152f $X=1.37 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A_M1009_g N_VGND_c_421_n 0.00383152f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A_M1011_g N_VGND_c_423_n 0.00434272f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A_M1013_g N_VGND_c_423_n 0.00434272f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A_c_68_n N_VGND_c_425_n 0.00434272f $X=0.51 $Y=1.2 $X2=0 $Y2=0
cc_182 N_A_c_69_n N_VGND_c_425_n 0.00383152f $X=0.94 $Y=1.2 $X2=0 $Y2=0
cc_183 N_A_M1014_g N_VGND_c_426_n 0.00434272f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A_M1015_g N_VGND_c_426_n 0.00383152f $X=3.73 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A_c_68_n N_VGND_c_428_n 0.00823992f $X=0.51 $Y=1.2 $X2=0 $Y2=0
cc_186 N_A_c_69_n N_VGND_c_428_n 0.0075754f $X=0.94 $Y=1.2 $X2=0 $Y2=0
cc_187 N_A_M1005_g N_VGND_c_428_n 0.0075754f $X=1.37 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A_M1009_g N_VGND_c_428_n 0.0075754f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A_M1011_g N_VGND_c_428_n 0.00820718f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A_M1013_g N_VGND_c_428_n 0.00821294f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A_M1014_g N_VGND_c_428_n 0.00821294f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A_M1015_g N_VGND_c_428_n 0.0075754f $X=3.73 $Y=0.74 $X2=0 $Y2=0
cc_193 N_VPWR_c_214_n N_Y_c_300_n 0.0121024f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_194 N_VPWR_c_214_n N_Y_c_293_n 0.0564818f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_195 N_VPWR_c_215_n N_Y_c_293_n 0.0462948f $X=1.18 $Y=2.455 $X2=0 $Y2=0
cc_196 N_VPWR_c_222_n N_Y_c_293_n 0.0110241f $X=1.015 $Y=3.33 $X2=0 $Y2=0
cc_197 N_VPWR_c_212_n N_Y_c_293_n 0.00909194f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_198 N_VPWR_M1002_d N_Y_c_312_n 0.00455969f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_199 N_VPWR_c_215_n N_Y_c_312_n 0.0202249f $X=1.18 $Y=2.455 $X2=0 $Y2=0
cc_200 N_VPWR_c_215_n N_Y_c_294_n 0.0266809f $X=1.18 $Y=2.455 $X2=0 $Y2=0
cc_201 N_VPWR_c_216_n N_Y_c_294_n 0.0462948f $X=2.13 $Y=2.455 $X2=0 $Y2=0
cc_202 N_VPWR_c_223_n N_Y_c_294_n 0.014552f $X=2.045 $Y=3.33 $X2=0 $Y2=0
cc_203 N_VPWR_c_212_n N_Y_c_294_n 0.0119791f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_204 N_VPWR_M1006_d N_Y_c_326_n 0.00384138f $X=1.98 $Y=1.84 $X2=0 $Y2=0
cc_205 N_VPWR_c_216_n N_Y_c_326_n 0.0154248f $X=2.13 $Y=2.455 $X2=0 $Y2=0
cc_206 N_VPWR_c_217_n N_Y_c_295_n 0.00846293f $X=3.03 $Y=1.985 $X2=0 $Y2=0
cc_207 N_VPWR_c_216_n N_Y_c_296_n 0.0440249f $X=2.13 $Y=2.455 $X2=0 $Y2=0
cc_208 N_VPWR_c_217_n N_Y_c_296_n 0.0560128f $X=3.03 $Y=1.985 $X2=0 $Y2=0
cc_209 N_VPWR_c_220_n N_Y_c_296_n 0.00749631f $X=2.865 $Y=3.33 $X2=0 $Y2=0
cc_210 N_VPWR_c_212_n N_Y_c_296_n 0.0062048f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_211 N_VPWR_c_217_n N_Y_c_287_n 0.0250577f $X=3.03 $Y=1.985 $X2=0 $Y2=0
cc_212 N_VPWR_c_217_n N_Y_c_297_n 0.0451069f $X=3.03 $Y=1.985 $X2=0 $Y2=0
cc_213 N_VPWR_c_219_n N_Y_c_297_n 0.0451069f $X=4.03 $Y=1.985 $X2=0 $Y2=0
cc_214 N_VPWR_c_224_n N_Y_c_297_n 0.014552f $X=3.865 $Y=3.33 $X2=0 $Y2=0
cc_215 N_VPWR_c_212_n N_Y_c_297_n 0.0119791f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_216 N_VPWR_c_217_n N_Y_c_389_n 0.0123817f $X=3.03 $Y=1.985 $X2=0 $Y2=0
cc_217 N_VPWR_c_219_n Y 0.0265821f $X=4.03 $Y=1.985 $X2=0 $Y2=0
cc_218 N_Y_c_282_n N_VGND_M1004_d 0.00176461f $X=1.5 $Y=1.095 $X2=0 $Y2=0
cc_219 N_Y_c_285_n N_VGND_M1009_d 0.00250873f $X=2.35 $Y=1.095 $X2=0 $Y2=0
cc_220 N_Y_c_281_n N_VGND_c_415_n 0.0233636f $X=0.725 $Y=0.515 $X2=0 $Y2=0
cc_221 N_Y_c_283_n N_VGND_c_415_n 0.00555794f $X=0.81 $Y=1.095 $X2=0 $Y2=0
cc_222 N_Y_c_281_n N_VGND_c_416_n 0.0182902f $X=0.725 $Y=0.515 $X2=0 $Y2=0
cc_223 N_Y_c_282_n N_VGND_c_416_n 0.0170777f $X=1.5 $Y=1.095 $X2=0 $Y2=0
cc_224 N_Y_c_284_n N_VGND_c_416_n 0.0182488f $X=1.585 $Y=0.515 $X2=0 $Y2=0
cc_225 N_Y_c_284_n N_VGND_c_417_n 0.0182488f $X=1.585 $Y=0.515 $X2=0 $Y2=0
cc_226 N_Y_c_285_n N_VGND_c_417_n 0.0209867f $X=2.35 $Y=1.095 $X2=0 $Y2=0
cc_227 N_Y_c_286_n N_VGND_c_417_n 0.0191765f $X=2.515 $Y=0.515 $X2=0 $Y2=0
cc_228 N_Y_c_286_n N_VGND_c_418_n 0.0240544f $X=2.515 $Y=0.515 $X2=0 $Y2=0
cc_229 N_Y_c_287_n N_VGND_c_418_n 0.028246f $X=3.35 $Y=1.38 $X2=0 $Y2=0
cc_230 N_Y_c_288_n N_VGND_c_418_n 0.0232199f $X=3.515 $Y=0.515 $X2=0 $Y2=0
cc_231 N_Y_c_288_n N_VGND_c_420_n 0.0240263f $X=3.515 $Y=0.515 $X2=0 $Y2=0
cc_232 Y N_VGND_c_420_n 0.026488f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_233 N_Y_c_284_n N_VGND_c_421_n 0.00749631f $X=1.585 $Y=0.515 $X2=0 $Y2=0
cc_234 N_Y_c_286_n N_VGND_c_423_n 0.0144922f $X=2.515 $Y=0.515 $X2=0 $Y2=0
cc_235 N_Y_c_281_n N_VGND_c_425_n 0.0109942f $X=0.725 $Y=0.515 $X2=0 $Y2=0
cc_236 N_Y_c_288_n N_VGND_c_426_n 0.0114405f $X=3.515 $Y=0.515 $X2=0 $Y2=0
cc_237 N_Y_c_281_n N_VGND_c_428_n 0.00904371f $X=0.725 $Y=0.515 $X2=0 $Y2=0
cc_238 N_Y_c_284_n N_VGND_c_428_n 0.0062048f $X=1.585 $Y=0.515 $X2=0 $Y2=0
cc_239 N_Y_c_286_n N_VGND_c_428_n 0.0118826f $X=2.515 $Y=0.515 $X2=0 $Y2=0
cc_240 N_Y_c_288_n N_VGND_c_428_n 0.00941304f $X=3.515 $Y=0.515 $X2=0 $Y2=0
