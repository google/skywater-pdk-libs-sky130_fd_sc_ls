* File: sky130_fd_sc_ls__a21o_1.pex.spice
* Created: Wed Sep  2 10:48:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__A21O_1%A_81_264# 1 2 7 9 10 12 14 15 24 26 30 32 34
+ 35
c61 35 0 1.84796e-19 $X=1.425 $Y=1.95
c62 10 0 8.11701e-20 $X=1.13 $Y=1.47
r63 34 35 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=2.115
+ $X2=1.425 $Y2=1.95
r64 28 30 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.97 $Y=1.11
+ $X2=1.97 $Y2=0.805
r65 27 32 3.70735 $w=2.5e-07 $l=2.23495e-07 $layer=LI1_cond $X=1.415 $Y=1.195
+ $X2=1.33 $Y2=1.38
r66 26 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.805 $Y=1.195
+ $X2=1.97 $Y2=1.11
r67 26 27 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.805 $Y=1.195
+ $X2=1.415 $Y2=1.195
r68 22 34 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=1.425 $Y=2.13
+ $X2=1.425 $Y2=2.115
r69 22 24 21.9284 $w=3.58e-07 $l=6.85e-07 $layer=LI1_cond $X=1.425 $Y=2.13
+ $X2=1.425 $Y2=2.815
r70 20 32 2.76166 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=1.33 $Y=1.65 $X2=1.33
+ $Y2=1.38
r71 20 35 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.33 $Y=1.65 $X2=1.33
+ $Y2=1.95
r72 18 36 2.36275 $w=3.06e-07 $l=1.5e-08 $layer=POLY_cond $X=0.58 $Y=1.485
+ $X2=0.58 $Y2=1.47
r73 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.485 $X2=0.59 $Y2=1.485
r74 15 32 3.70735 $w=2.5e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.245 $Y=1.485
+ $X2=1.33 $Y2=1.38
r75 15 17 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=1.245 $Y=1.485
+ $X2=0.59 $Y2=1.485
r76 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.205 $Y=1.395
+ $X2=1.205 $Y2=0.95
r77 11 36 19.4347 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.755 $Y=1.47
+ $X2=0.58 $Y2=1.47
r78 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.13 $Y=1.47
+ $X2=1.205 $Y2=1.395
r79 10 11 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.13 $Y=1.47
+ $X2=0.755 $Y2=1.47
r80 7 18 56.6494 $w=3.06e-07 $l=3.19687e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.58 $Y2=1.485
r81 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
r82 2 34 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=1.96 $X2=1.52 $Y2=2.115
r83 2 24 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=1.96 $X2=1.52 $Y2=2.815
r84 1 30 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.83
+ $Y=0.68 $X2=1.97 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LS__A21O_1%B1 1 3 6 8
c31 8 0 8.11701e-20 $X=1.68 $Y=1.665
r32 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.615 $X2=1.67 $Y2=1.615
r33 4 11 38.5916 $w=2.93e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.755 $Y=1.45
+ $X2=1.67 $Y2=1.615
r34 4 6 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.755 $Y=1.45
+ $X2=1.755 $Y2=1
r35 1 11 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=1.745 $Y=1.885
+ $X2=1.67 $Y2=1.615
r36 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.745 $Y=1.885
+ $X2=1.745 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__A21O_1%A1 3 5 7 8
c34 5 0 4.69421e-20 $X=2.195 $Y=1.885
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.615 $X2=2.21 $Y2=1.615
r36 5 11 55.8646 $w=2.93e-07 $l=2.77399e-07 $layer=POLY_cond $X=2.195 $Y=1.885
+ $X2=2.21 $Y2=1.615
r37 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.195 $Y=1.885
+ $X2=2.195 $Y2=2.46
r38 1 11 38.5916 $w=2.93e-07 $l=1.77059e-07 $layer=POLY_cond $X=2.185 $Y=1.45
+ $X2=2.21 $Y2=1.615
r39 1 3 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.185 $Y=1.45
+ $X2=2.185 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_LS__A21O_1%A2 4 5 6 7 9 14 16 23
r36 16 23 3.89033 $w=4.13e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=0.462
+ $X2=3.005 $Y2=0.462
r37 14 18 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.81 $Y=0.405
+ $X2=2.66 $Y2=0.405
r38 13 23 7.13417 $w=3.13e-07 $l=1.95e-07 $layer=LI1_cond $X=2.81 $Y=0.412
+ $X2=3.005 $Y2=0.412
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.81
+ $Y=0.405 $X2=2.81 $Y2=0.405
r40 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.675 $Y=1.885
+ $X2=2.675 $Y2=2.46
r41 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.675 $Y=1.795 $X2=2.675
+ $Y2=1.885
r42 5 10 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.675 $Y=1.485
+ $X2=2.675 $Y2=1.395
r43 5 6 120.5 $w=1.8e-07 $l=3.1e-07 $layer=POLY_cond $X=2.675 $Y=1.485 $X2=2.675
+ $Y2=1.795
r44 4 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.66 $Y=1 $X2=2.66
+ $Y2=1.395
r45 1 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.66 $Y=0.57
+ $X2=2.66 $Y2=0.405
r46 1 4 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.66 $Y=0.57 $X2=2.66
+ $Y2=1
.ends

.subckt PM_SKY130_FD_SC_LS__A21O_1%X 1 2 9 10 13 15 16 17 24 33
r20 22 24 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=0.26 $Y=1.995 $X2=0.26
+ $Y2=2.035
r21 16 17 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.405
+ $X2=0.26 $Y2=2.775
r22 15 22 0.75732 $w=3.48e-07 $l=2.3e-08 $layer=LI1_cond $X=0.26 $Y=1.972
+ $X2=0.26 $Y2=1.995
r23 15 33 8.06043 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=0.26 $Y=1.972
+ $X2=0.26 $Y2=1.82
r24 15 16 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=0.26 $Y=2.057
+ $X2=0.26 $Y2=2.405
r25 15 24 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=0.26 $Y=2.057
+ $X2=0.26 $Y2=2.035
r26 11 13 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=0.95 $Y=0.98
+ $X2=0.95 $Y2=0.885
r27 9 11 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.825 $Y=1.065
+ $X2=0.95 $Y2=0.98
r28 9 10 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=0.825 $Y=1.065
+ $X2=0.255 $Y2=1.065
r29 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.15
+ $X2=0.255 $Y2=1.065
r30 7 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=1.15 $X2=0.17
+ $Y2=1.82
r31 2 15 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=1.985
r32 2 17 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.815
r33 1 13 182 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_NDIFF $count=1 $X=0.865
+ $Y=0.58 $X2=0.99 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_LS__A21O_1%VPWR 1 2 9 15 18 19 20 22 35 36 39
r36 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r42 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r43 27 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.76 $Y2=3.33
r44 27 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 22 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.76 $Y2=3.33
r48 22 24 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 20 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 20 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 18 32 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 18 19 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.335 $Y=3.33 $X2=2.435
+ $Y2=3.33
r53 17 35 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.535 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 17 19 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.535 $Y=3.33 $X2=2.435
+ $Y2=3.33
r55 13 19 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=3.245
+ $X2=2.435 $Y2=3.33
r56 13 15 43.8091 $w=1.98e-07 $l=7.9e-07 $layer=LI1_cond $X=2.435 $Y=3.245
+ $X2=2.435 $Y2=2.455
r57 9 12 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.76 $Y=1.985
+ $X2=0.76 $Y2=2.815
r58 7 39 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=3.33
r59 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.76 $Y=3.245 $X2=0.76
+ $Y2=2.815
r60 2 15 300 $w=1.7e-07 $l=5.71577e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=1.96 $X2=2.435 $Y2=2.455
r61 1 12 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.815
r62 1 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__A21O_1%A_364_392# 1 2 7 9 11 13 15
c31 13 0 4.69421e-20 $X=2.9 $Y=2.12
r32 13 20 2.68829 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.9 $Y=2.12 $X2=2.9
+ $Y2=2.03
r33 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.9 $Y=2.12 $X2=2.9
+ $Y2=2.815
r34 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=2.035
+ $X2=1.97 $Y2=2.035
r35 11 20 5.07788 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=2.735 $Y=2.035
+ $X2=2.9 $Y2=2.03
r36 11 12 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.735 $Y=2.035
+ $X2=2.135 $Y2=2.035
r37 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.97 $Y=2.12 $X2=1.97
+ $Y2=2.035
r38 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.97 $Y=2.12 $X2=1.97
+ $Y2=2.815
r39 2 20 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.75
+ $Y=1.96 $X2=2.9 $Y2=2.105
r40 2 15 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.75
+ $Y=1.96 $X2=2.9 $Y2=2.815
r41 1 18 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=1.82
+ $Y=1.96 $X2=1.97 $Y2=2.115
r42 1 9 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.82
+ $Y=1.96 $X2=1.97 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__A21O_1%VGND 1 2 9 12 13 14 16 17 19 20 21 26 39 40
r52 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r53 37 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r54 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r55 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r56 30 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r57 29 33 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r58 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r59 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r60 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r61 21 24 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=0.925
+ $X2=2.875 $Y2=1.09
r62 19 36 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.16
+ $Y2=0
r63 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.39
+ $Y2=0
r64 18 39 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=3.12
+ $Y2=0
r65 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.39
+ $Y2=0
r66 16 33 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.2
+ $Y2=0
r67 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.42
+ $Y2=0
r68 15 36 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1.585 $Y=0 $X2=2.16
+ $Y2=0
r69 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.585 $Y=0 $X2=1.42
+ $Y2=0
r70 13 21 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0.925
+ $X2=2.875 $Y2=0.925
r71 13 14 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.71 $Y=0.925
+ $X2=2.475 $Y2=0.925
r72 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.39 $Y=0.84
+ $X2=2.475 $Y2=0.925
r73 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=0.085
+ $X2=2.39 $Y2=0
r74 11 12 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.39 $Y=0.085
+ $X2=2.39 $Y2=0.84
r75 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.42 $Y=0.085 $X2=1.42
+ $Y2=0
r76 7 9 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=1.42 $Y=0.085 $X2=1.42
+ $Y2=0.775
r77 2 24 182 $w=1.7e-07 $l=4.74868e-07 $layer=licon1_NDIFF $count=1 $X=2.735
+ $Y=0.68 $X2=2.875 $Y2=1.09
r78 1 9 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.28
+ $Y=0.58 $X2=1.42 $Y2=0.775
.ends

