* File: sky130_fd_sc_ls__dfxtp_4.spice
* Created: Fri Aug 28 13:16:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__dfxtp_4.pex.spice"
.subckt sky130_fd_sc_ls__dfxtp_4  VNB VPB CLK D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1025 N_VGND_M1025_d N_CLK_M1025_g N_A_27_74#_M1025_s VNB NSHORT L=0.15 W=0.74
+ AD=0.17575 AS=0.2109 PD=1.215 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1022 N_A_206_368#_M1022_d N_A_27_74#_M1022_g N_VGND_M1025_d VNB NSHORT L=0.15
+ W=0.74 AD=0.2516 AS=0.17575 PD=2.16 PS=1.215 NRD=8.916 NRS=31.62 M=1 R=4.93333
+ SA=75000.8 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1019 N_A_437_503#_M1019_d N_D_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.355025 PD=0.7 PS=2.6 NRD=0 NRS=225.792 M=1 R=2.8 SA=75000.5
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1020 N_A_544_485#_M1020_d N_A_27_74#_M1020_g N_A_437_503#_M1019_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0756875 AS=0.0588 PD=0.83 PS=0.7 NRD=4.284 NRS=0 M=1 R=2.8
+ SA=75001 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1017 A_735_102# N_A_206_368#_M1017_g N_A_544_485#_M1020_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0756875 PD=0.63 PS=0.83 NRD=14.28 NRS=8.568 M=1 R=2.8
+ SA=75001.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_696_458#_M1011_g A_735_102# VNB NSHORT L=0.15 W=0.42
+ AD=0.170728 AS=0.0441 PD=1.18206 PS=0.63 NRD=100.416 NRS=14.28 M=1 R=2.8
+ SA=75001.5 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_696_458#_M1005_d N_A_544_485#_M1005_g N_VGND_M1011_d VNB NSHORT
+ L=0.15 W=0.55 AD=0.099 AS=0.223572 PD=0.985 PS=1.54794 NRD=0 NRS=76.68 M=1
+ R=3.66667 SA=75001.9 SB=75001.2 A=0.0825 P=1.4 MULT=1
MM1021 N_A_1034_424#_M1021_d N_A_206_368#_M1021_g N_A_696_458#_M1005_d VNB
+ NSHORT L=0.15 W=0.55 AD=0.122021 AS=0.099 PD=1.11701 PS=0.985 NRD=24 NRS=0 M=1
+ R=3.66667 SA=75002.2 SB=75001 A=0.0825 P=1.4 MULT=1
MM1028 A_1178_124# N_A_27_74#_M1028_g N_A_1034_424#_M1021_d VNB NSHORT L=0.15
+ W=0.42 AD=0.06615 AS=0.0931794 PD=0.735 PS=0.85299 NRD=29.28 NRS=12.852 M=1
+ R=2.8 SA=75002.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_1226_296#_M1014_g A_1178_124# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.06615 PD=1.41 PS=0.735 NRD=0 NRS=29.28 M=1 R=2.8 SA=75003.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_1034_424#_M1024_g N_A_1226_296#_M1024_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.1147 AS=0.2109 PD=1.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1000 N_Q_M1000_d N_A_1226_296#_M1000_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1184 AS=0.1147 PD=1.06 PS=1.05 NRD=6.48 NRS=4.86 M=1 R=4.93333 SA=75000.7
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1004 N_Q_M1000_d N_A_1226_296#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1184 AS=0.111 PD=1.06 PS=1.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1012 N_Q_M1012_d N_A_1226_296#_M1012_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.111 PD=1.02 PS=1.04 NRD=0 NRS=3.24 M=1 R=4.93333 SA=75001.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1030 N_Q_M1012_d N_A_1226_296#_M1030_g N_VGND_M1030_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VPWR_M1015_d N_CLK_M1015_g N_A_27_74#_M1015_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1016 N_A_206_368#_M1016_d N_A_27_74#_M1016_g N_VPWR_M1015_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1008 N_A_437_503#_M1008_d N_D_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.088725 AS=0.2544 PD=0.895 PS=2.2 NRD=46.886 NRS=258.306 M=1 R=2.8
+ SA=75000.4 SB=75005.5 A=0.063 P=1.14 MULT=1
MM1010 N_A_544_485#_M1010_d N_A_206_368#_M1010_g N_A_437_503#_M1008_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.088725 AS=0.088725 PD=0.895 PS=0.895 NRD=4.6886
+ NRS=4.6886 M=1 R=2.8 SA=75000.8 SB=75005 A=0.063 P=1.14 MULT=1
MM1006 A_651_503# N_A_27_74#_M1006_g N_A_544_485#_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.088725 PD=0.66 PS=0.895 NRD=30.4759 NRS=44.5417 M=1
+ R=2.8 SA=75001.2 SB=75005.9 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_696_458#_M1009_g A_651_503# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1599 AS=0.0504 PD=1.15667 PS=0.66 NRD=152.773 NRS=30.4759 M=1 R=2.8
+ SA=75001.6 SB=75005.5 A=0.063 P=1.14 MULT=1
MM1027 N_A_696_458#_M1027_d N_A_544_485#_M1027_g N_VPWR_M1009_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.3198 PD=1.37 PS=2.31333 NRD=0 NRS=76.3769 M=1
+ R=5.6 SA=75001.3 SB=75002.9 A=0.126 P=1.98 MULT=1
MM1018 N_A_1034_424#_M1018_d N_A_27_74#_M1018_g N_A_696_458#_M1027_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1904 AS=0.2226 PD=1.63333 PS=1.37 NRD=2.3443 NRS=56.2829
+ M=1 R=5.6 SA=75002 SB=75002.2 A=0.126 P=1.98 MULT=1
MM1001 A_1141_508# N_A_206_368#_M1001_g N_A_1034_424#_M1018_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.09975 AS=0.0952 PD=0.895 PS=0.816667 NRD=85.5965 NRS=80.5139 M=1
+ R=2.8 SA=75003.5 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1023 N_VPWR_M1023_d N_A_1226_296#_M1023_g A_1141_508# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0868 AS=0.09975 PD=0.796667 PS=0.895 NRD=7.0329 NRS=85.5965 M=1
+ R=2.8 SA=75004.1 SB=75003.1 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1023_d N_A_1034_424#_M1003_g N_A_1226_296#_M1003_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1736 AS=0.126 PD=1.59333 PS=1.14 NRD=14.0658 NRS=2.3443 M=1
+ R=5.6 SA=75002.4 SB=75002.6 A=0.126 P=1.98 MULT=1
MM1029 N_VPWR_M1029_d N_A_1034_424#_M1029_g N_A_1226_296#_M1003_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.174 AS=0.126 PD=1.29 PS=1.14 NRD=22.261 NRS=2.3443 M=1
+ R=5.6 SA=75002.9 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1002 N_Q_M1002_d N_A_1226_296#_M1002_g N_VPWR_M1029_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.232 PD=1.42 PS=1.72 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.6 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1007 N_Q_M1002_d N_A_1226_296#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1013 N_Q_M1013_d N_A_1226_296#_M1013_g N_VPWR_M1007_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1026 N_Q_M1013_d N_A_1226_296#_M1026_g N_VPWR_M1026_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.9 SB=75000.2 A=0.168 P=2.54 MULT=1
DX31_noxref VNB VPB NWDIODE A=18.5628 P=23.68
c_212 VPB 0 1.17955e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__dfxtp_4.pxi.spice"
*
.ends
*
*
