* NGSPICE file created from sky130_fd_sc_ls__o221ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 Y C1 a_27_84# VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=1.4578e+12p ps=1.43e+07u
M1001 a_508_368# B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=1.4e+12p pd=1.146e+07u as=2.716e+12p ps=2.053e+07u
M1002 Y C1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=2.1e+12p pd=1.719e+07u as=0p ps=0u
M1003 a_483_74# B2 a_27_84# VNB nshort w=740000u l=150000u
+  ad=1.9758e+12p pd=1.866e+07u as=0p ps=0u
M1004 VGND A2 a_483_74# VNB nshort w=740000u l=150000u
+  ad=9.916e+11p pd=8.6e+06u as=0p ps=0u
M1005 a_483_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B2 a_508_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A2 a_1288_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=1.4056e+12p ps=1.147e+07u
M1008 a_27_84# B1 a_483_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_84# B1 a_483_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_508_368# B2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_483_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR B1 a_508_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1288_368# A2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR B1 a_508_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_483_74# B2 a_27_84# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_508_368# B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_84# B2 a_483_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_483_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1288_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A1 a_1288_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y C1 a_27_84# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A2 a_483_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y C1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR C1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR A1 a_1288_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y B2 a_508_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y A2 a_1288_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_27_84# B2 a_483_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND A1 a_483_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_483_74# B1 a_27_84# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND A1 a_483_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR C1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1288_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_483_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_483_74# B1 a_27_84# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_508_368# B2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1288_368# A2 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_27_84# C1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_27_84# C1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

