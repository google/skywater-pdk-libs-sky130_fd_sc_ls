# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__fa_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__fa_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.044000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.245000 0.835000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.044000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345000 1.260000 1.835000 1.575000 ;
        RECT 1.665000 1.575000 1.835000 1.950000 ;
        RECT 1.665000 1.950000 2.650000 2.120000 ;
        RECT 2.480000 1.245000 2.810000 1.745000 ;
        RECT 2.480000 1.745000 6.595000 1.780000 ;
        RECT 2.480000 1.780000 6.085000 1.890000 ;
        RECT 2.480000 1.890000 4.620000 1.915000 ;
        RECT 2.480000 1.915000 2.650000 1.950000 ;
        RECT 3.950000 1.260000 4.280000 1.745000 ;
        RECT 4.450000 1.720000 6.595000 1.745000 ;
        RECT 5.915000 1.260000 6.340000 1.550000 ;
        RECT 5.915000 1.550000 6.595000 1.720000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.783000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005000 1.180000 2.275000 1.780000 ;
        RECT 3.005000 1.180000 3.215000 1.260000 ;
        RECT 3.005000 1.260000 3.740000 1.575000 ;
        RECT 5.430000 1.180000 5.745000 1.550000 ;
      LAYER mcon ;
        RECT 2.075000 1.210000 2.245000 1.380000 ;
        RECT 3.035000 1.210000 3.205000 1.380000 ;
        RECT 5.435000 1.210000 5.605000 1.380000 ;
      LAYER met1 ;
        RECT 2.015000 1.180000 2.305000 1.225000 ;
        RECT 2.015000 1.225000 5.665000 1.365000 ;
        RECT 2.015000 1.365000 2.305000 1.410000 ;
        RECT 2.975000 1.180000 3.265000 1.225000 ;
        RECT 2.975000 1.365000 3.265000 1.410000 ;
        RECT 5.375000 1.180000 5.665000 1.225000 ;
        RECT 5.375000 1.365000 5.665000 1.410000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.145000 1.820000 10.435000 1.990000 ;
        RECT  9.145000 1.990000  9.475000 2.980000 ;
        RECT  9.305000 0.390000  9.555000 0.980000 ;
        RECT  9.305000 0.980000 10.425000 1.150000 ;
        RECT 10.095000 1.990000 10.435000 2.980000 ;
        RECT 10.165000 0.390000 10.425000 0.980000 ;
        RECT 10.165000 1.150000 10.425000 1.550000 ;
        RECT 10.165000 1.550000 10.435000 1.820000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.245000 1.840000 8.525000 2.010000 ;
        RECT 7.245000 2.010000 7.575000 2.980000 ;
        RECT 7.265000 0.920000 8.615000 1.170000 ;
        RECT 8.195000 2.010000 8.525000 2.980000 ;
        RECT 8.285000 1.170000 8.525000 1.840000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.040000 0.085000 ;
        RECT  0.625000  0.085000  1.155000 0.410000 ;
        RECT  3.175000  0.085000  3.505000 0.670000 ;
        RECT  4.155000  0.085000  4.485000 0.410000 ;
        RECT  6.755000  0.085000  7.085000 0.410000 ;
        RECT  7.775000  0.085000  8.105000 0.410000 ;
        RECT  8.795000  0.085000  9.125000 0.410000 ;
        RECT  9.735000  0.085000  9.985000 0.810000 ;
        RECT 10.595000  0.085000 10.925000 1.170000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 11.040000 3.415000 ;
        RECT  0.645000 2.425000  0.815000 3.245000 ;
        RECT  3.170000 2.085000  3.500000 3.245000 ;
        RECT  4.170000 2.425000  4.570000 3.245000 ;
        RECT  6.795000 2.290000  7.045000 3.245000 ;
        RECT  7.775000 2.180000  8.025000 3.245000 ;
        RECT  8.725000 1.820000  8.975000 3.245000 ;
        RECT  9.675000 2.160000  9.925000 3.245000 ;
        RECT 10.625000 1.820000 10.875000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.350000 0.445000 0.580000 ;
      RECT 0.115000 0.580000 1.965000 0.670000 ;
      RECT 0.115000 0.670000 1.495000 0.750000 ;
      RECT 0.115000 0.750000 0.445000 1.075000 ;
      RECT 0.115000 1.950000 0.445000 2.085000 ;
      RECT 0.115000 2.085000 1.155000 2.255000 ;
      RECT 0.115000 2.255000 0.445000 2.980000 ;
      RECT 0.985000 2.255000 1.155000 2.630000 ;
      RECT 0.985000 2.630000 2.005000 2.960000 ;
      RECT 1.005000 0.920000 5.255000 1.010000 ;
      RECT 1.005000 1.010000 1.835000 1.090000 ;
      RECT 1.005000 1.090000 1.175000 1.745000 ;
      RECT 1.005000 1.745000 1.495000 1.915000 ;
      RECT 1.325000 0.350000 1.965000 0.580000 ;
      RECT 1.325000 1.915000 1.495000 2.290000 ;
      RECT 1.325000 2.290000 2.540000 2.460000 ;
      RECT 1.665000 0.840000 3.555000 0.920000 ;
      RECT 2.135000 0.350000 2.465000 0.840000 ;
      RECT 2.210000 2.460000 2.540000 2.755000 ;
      RECT 3.385000 1.010000 5.255000 1.090000 ;
      RECT 3.670000 2.085000 5.070000 2.255000 ;
      RECT 3.670000 2.255000 4.000000 2.755000 ;
      RECT 3.725000 0.350000 3.975000 0.580000 ;
      RECT 3.725000 0.580000 4.915000 0.750000 ;
      RECT 4.665000 0.350000 4.915000 0.580000 ;
      RECT 4.740000 2.255000 5.070000 2.755000 ;
      RECT 4.930000 1.090000 5.255000 1.220000 ;
      RECT 4.930000 1.220000 5.260000 1.550000 ;
      RECT 5.085000 0.255000 6.425000 0.425000 ;
      RECT 5.085000 0.425000 5.255000 0.920000 ;
      RECT 5.240000 2.060000 7.075000 2.120000 ;
      RECT 5.240000 2.120000 6.425000 2.230000 ;
      RECT 5.240000 2.230000 5.570000 2.755000 ;
      RECT 5.425000 0.595000 5.675000 0.840000 ;
      RECT 5.425000 0.840000 6.085000 0.920000 ;
      RECT 5.425000 0.920000 7.075000 1.010000 ;
      RECT 5.915000 1.010000 7.075000 1.090000 ;
      RECT 6.255000 0.425000 6.425000 0.580000 ;
      RECT 6.255000 0.580000 9.135000 0.750000 ;
      RECT 6.255000 1.950000 7.075000 2.060000 ;
      RECT 6.905000 1.090000 7.075000 1.340000 ;
      RECT 6.905000 1.340000 8.105000 1.670000 ;
      RECT 6.905000 1.670000 7.075000 1.950000 ;
      RECT 8.965000 0.750000 9.135000 1.320000 ;
      RECT 8.965000 1.320000 9.955000 1.650000 ;
  END
END sky130_fd_sc_ls__fa_4
