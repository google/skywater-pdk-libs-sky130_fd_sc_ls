* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_69_392# C1 a_154_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_154_392# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 X a_154_392# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 a_334_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_1081_39# A2 a_888_105# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_1081_39# A1 a_154_392# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 VPWR A1 a_334_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_154_392# C1 a_69_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_154_392# A1 a_1081_39# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 VPWR a_154_392# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X10 VGND C1 a_154_392# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 VPWR A2 a_334_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_154_392# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 VPWR a_154_392# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 VGND a_154_392# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 VGND A3 a_888_105# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 X a_154_392# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 VGND a_154_392# X VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X18 VPWR A3 a_334_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_154_392# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 a_334_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_888_105# A2 a_1081_39# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 a_334_392# B1 a_69_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 VGND B1 a_154_392# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 a_888_105# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 a_69_392# B1 a_334_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_334_392# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 X a_154_392# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
.ends
