* File: sky130_fd_sc_ls__or3_4.pxi.spice
* Created: Wed Sep  2 11:24:59 2020
* 
x_PM_SKY130_FD_SC_LS__OR3_4%A N_A_c_93_n N_A_c_105_n N_A_M1002_g N_A_c_94_n
+ N_A_c_107_n N_A_M1006_g N_A_M1004_g N_A_c_95_n N_A_c_96_n N_A_c_97_n
+ N_A_c_98_n N_A_c_99_n A N_A_c_101_n N_A_c_102_n A PM_SKY130_FD_SC_LS__OR3_4%A
x_PM_SKY130_FD_SC_LS__OR3_4%B N_B_c_187_n N_B_M1000_g N_B_c_188_n N_B_M1003_g
+ N_B_M1012_g B B B B N_B_c_190_n PM_SKY130_FD_SC_LS__OR3_4%B
x_PM_SKY130_FD_SC_LS__OR3_4%C N_C_c_246_n N_C_c_253_n N_C_M1013_g N_C_c_247_n
+ N_C_c_255_n N_C_M1016_g N_C_c_248_n N_C_M1008_g N_C_c_249_n C N_C_c_250_n
+ N_C_c_251_n PM_SKY130_FD_SC_LS__OR3_4%C
x_PM_SKY130_FD_SC_LS__OR3_4%A_302_388# N_A_302_388#_M1008_s N_A_302_388#_M1012_d
+ N_A_302_388#_M1013_d N_A_302_388#_c_314_n N_A_302_388#_M1005_g
+ N_A_302_388#_M1001_g N_A_302_388#_M1007_g N_A_302_388#_c_315_n
+ N_A_302_388#_M1010_g N_A_302_388#_c_316_n N_A_302_388#_M1011_g
+ N_A_302_388#_M1009_g N_A_302_388#_c_317_n N_A_302_388#_M1014_g
+ N_A_302_388#_M1015_g N_A_302_388#_c_307_n N_A_302_388#_c_326_n
+ N_A_302_388#_c_330_n N_A_302_388#_c_308_n N_A_302_388#_c_309_n
+ N_A_302_388#_c_333_n N_A_302_388#_c_310_n N_A_302_388#_c_311_n
+ N_A_302_388#_c_404_p N_A_302_388#_c_355_n N_A_302_388#_c_341_n
+ N_A_302_388#_c_312_n N_A_302_388#_c_313_n PM_SKY130_FD_SC_LS__OR3_4%A_302_388#
x_PM_SKY130_FD_SC_LS__OR3_4%VPWR N_VPWR_M1002_s N_VPWR_M1006_s N_VPWR_M1010_s
+ N_VPWR_M1014_s N_VPWR_c_470_n N_VPWR_c_471_n N_VPWR_c_472_n N_VPWR_c_473_n
+ N_VPWR_c_474_n N_VPWR_c_475_n VPWR N_VPWR_c_476_n N_VPWR_c_477_n
+ N_VPWR_c_478_n N_VPWR_c_479_n N_VPWR_c_480_n N_VPWR_c_469_n
+ PM_SKY130_FD_SC_LS__OR3_4%VPWR
x_PM_SKY130_FD_SC_LS__OR3_4%A_116_388# N_A_116_388#_M1002_d N_A_116_388#_M1003_d
+ N_A_116_388#_c_541_n N_A_116_388#_c_539_n N_A_116_388#_c_550_n
+ N_A_116_388#_c_544_n N_A_116_388#_c_540_n N_A_116_388#_c_546_n
+ PM_SKY130_FD_SC_LS__OR3_4%A_116_388#
x_PM_SKY130_FD_SC_LS__OR3_4%A_206_388# N_A_206_388#_M1000_s N_A_206_388#_M1016_s
+ N_A_206_388#_c_576_n PM_SKY130_FD_SC_LS__OR3_4%A_206_388#
x_PM_SKY130_FD_SC_LS__OR3_4%X N_X_M1001_d N_X_M1009_d N_X_M1005_d N_X_M1011_d
+ N_X_c_590_n N_X_c_597_n N_X_c_591_n N_X_c_592_n N_X_c_598_n N_X_c_599_n
+ N_X_c_600_n N_X_c_593_n N_X_c_594_n N_X_c_601_n N_X_c_602_n N_X_c_595_n X X
+ PM_SKY130_FD_SC_LS__OR3_4%X
x_PM_SKY130_FD_SC_LS__OR3_4%VGND N_VGND_M1008_d N_VGND_M1004_d N_VGND_M1007_s
+ N_VGND_M1015_s N_VGND_c_673_n N_VGND_c_674_n N_VGND_c_675_n N_VGND_c_676_n
+ N_VGND_c_677_n N_VGND_c_678_n VGND N_VGND_c_679_n N_VGND_c_680_n
+ N_VGND_c_681_n N_VGND_c_682_n N_VGND_c_683_n N_VGND_c_684_n N_VGND_c_685_n
+ PM_SKY130_FD_SC_LS__OR3_4%VGND
cc_1 VNB N_A_c_93_n 0.00241604f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.775
cc_2 VNB N_A_c_94_n 0.00642334f $X=-0.19 $Y=-0.245 $X2=2.89 $Y2=1.775
cc_3 VNB N_A_c_95_n 0.00249471f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.445
cc_4 VNB N_A_c_96_n 0.156212f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.445
cc_5 VNB N_A_c_97_n 0.0390478f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=1.195
cc_6 VNB N_A_c_98_n 0.00249596f $X=-0.19 $Y=-0.245 $X2=2.905 $Y2=1.195
cc_7 VNB N_A_c_99_n 0.032308f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=1.385
cc_8 VNB A 0.00692367f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_9 VNB N_A_c_101_n 0.0410223f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_10 VNB N_A_c_102_n 0.0176807f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=1.22
cc_11 VNB A 0.00534102f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.295
cc_12 VNB N_B_c_187_n 0.0192391f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.63
cc_13 VNB N_B_c_188_n 0.0165947f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.44
cc_14 VNB N_B_M1012_g 0.0292678f $X=-0.19 $Y=-0.245 $X2=2.89 $Y2=2.44
cc_15 VNB N_B_c_190_n 0.00863455f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=1.385
cc_16 VNB N_C_c_246_n 0.00649245f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.775
cc_17 VNB N_C_c_247_n 0.00671204f $X=-0.19 $Y=-0.245 $X2=2.89 $Y2=1.775
cc_18 VNB N_C_c_248_n 0.0167983f $X=-0.19 $Y=-0.245 $X2=2.93 $Y2=1.22
cc_19 VNB N_C_c_249_n 0.0571927f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.445
cc_20 VNB N_C_c_250_n 0.0972169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_C_c_251_n 0.00245092f $X=-0.19 $Y=-0.245 $X2=2.905 $Y2=1.385
cc_22 VNB N_A_302_388#_M1001_g 0.0204334f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.445
cc_23 VNB N_A_302_388#_M1007_g 0.0211635f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=1.195
cc_24 VNB N_A_302_388#_M1009_g 0.02167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_302_388#_M1015_g 0.0232609f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.465
cc_26 VNB N_A_302_388#_c_307_n 0.00530233f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=1.385
cc_27 VNB N_A_302_388#_c_308_n 0.00124938f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.295
cc_28 VNB N_A_302_388#_c_309_n 0.00279725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_302_388#_c_310_n 0.00113959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_302_388#_c_311_n 2.94743e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_302_388#_c_312_n 0.00237265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_302_388#_c_313_n 0.104036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_469_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_590_n 0.0017961f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.445
cc_35 VNB N_X_c_591_n 0.00311091f $X=-0.19 $Y=-0.245 $X2=2.905 $Y2=1.385
cc_36 VNB N_X_c_592_n 0.00138775f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=1.385
cc_37 VNB N_X_c_593_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_38 VNB N_X_c_594_n 0.00874592f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_39 VNB N_X_c_595_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=1.55
cc_40 VNB X 0.0264317f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.295
cc_41 VNB N_VGND_c_673_n 0.00595424f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.445
cc_42 VNB N_VGND_c_674_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.445
cc_43 VNB N_VGND_c_675_n 0.00499383f $X=-0.19 $Y=-0.245 $X2=2.905 $Y2=1.195
cc_44 VNB N_VGND_c_676_n 0.00425095f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=1.385
cc_45 VNB N_VGND_c_677_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_46 VNB N_VGND_c_678_n 0.0258474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_679_n 0.0588809f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.125
cc_48 VNB N_VGND_c_680_n 0.0153327f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=1.22
cc_49 VNB N_VGND_c_681_n 0.0191617f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.33
cc_50 VNB N_VGND_c_682_n 0.00614151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_683_n 0.00613227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_684_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_685_n 0.320708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VPB N_A_c_93_n 0.00949753f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.775
cc_55 VPB N_A_c_105_n 0.0256936f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.865
cc_56 VPB N_A_c_94_n 0.00672248f $X=-0.19 $Y=1.66 $X2=2.89 $Y2=1.775
cc_57 VPB N_A_c_107_n 0.0222666f $X=-0.19 $Y=1.66 $X2=2.89 $Y2=1.865
cc_58 VPB N_B_c_187_n 0.0326652f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.63
cc_59 VPB N_B_c_188_n 0.0325849f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.44
cc_60 VPB N_B_c_190_n 0.012713f $X=-0.19 $Y=1.66 $X2=2.92 $Y2=1.385
cc_61 VPB N_C_c_246_n 0.0048061f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.775
cc_62 VPB N_C_c_253_n 0.020717f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.865
cc_63 VPB N_C_c_247_n 0.00496865f $X=-0.19 $Y=1.66 $X2=2.89 $Y2=1.775
cc_64 VPB N_C_c_255_n 0.020853f $X=-0.19 $Y=1.66 $X2=2.89 $Y2=1.865
cc_65 VPB N_A_302_388#_c_314_n 0.0155697f $X=-0.19 $Y=1.66 $X2=2.89 $Y2=2.44
cc_66 VPB N_A_302_388#_c_315_n 0.0147322f $X=-0.19 $Y=1.66 $X2=2.905 $Y2=1.195
cc_67 VPB N_A_302_388#_c_316_n 0.0152457f $X=-0.19 $Y=1.66 $X2=2.92 $Y2=1.385
cc_68 VPB N_A_302_388#_c_317_n 0.0164089f $X=-0.19 $Y=1.66 $X2=0.35 $Y2=0.445
cc_69 VPB N_A_302_388#_c_311_n 0.00182944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_302_388#_c_313_n 0.0262207f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_470_n 0.0106521f $X=-0.19 $Y=1.66 $X2=2.93 $Y2=0.74
cc_72 VPB N_VPWR_c_471_n 0.0535635f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.445
cc_73 VPB N_VPWR_c_472_n 0.00654918f $X=-0.19 $Y=1.66 $X2=2.905 $Y2=1.195
cc_74 VPB N_VPWR_c_473_n 0.00504372f $X=-0.19 $Y=1.66 $X2=2.92 $Y2=1.385
cc_75 VPB N_VPWR_c_474_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_76 VPB N_VPWR_c_475_n 0.0428822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_476_n 0.0707163f $X=-0.19 $Y=1.66 $X2=0.35 $Y2=1.125
cc_78 VPB N_VPWR_c_477_n 0.0164465f $X=-0.19 $Y=1.66 $X2=2.92 $Y2=1.22
cc_79 VPB N_VPWR_c_478_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.33
cc_80 VPB N_VPWR_c_479_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_480_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_469_n 0.091515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_116_388#_c_539_n 0.00223287f $X=-0.19 $Y=1.66 $X2=2.93 $Y2=0.74
cc_84 VPB N_A_116_388#_c_540_n 0.00298259f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=1.195
cc_85 VPB N_A_206_388#_c_576_n 0.00859266f $X=-0.19 $Y=1.66 $X2=2.93 $Y2=1.22
cc_86 VPB N_X_c_597_n 0.00180921f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=1.195
cc_87 VPB N_X_c_598_n 0.00217622f $X=-0.19 $Y=1.66 $X2=2.92 $Y2=1.385
cc_88 VPB N_X_c_599_n 0.00133248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_X_c_600_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_X_c_601_n 0.00826668f $X=-0.19 $Y=1.66 $X2=0.35 $Y2=1.63
cc_91 VPB N_X_c_602_n 0.00187476f $X=-0.19 $Y=1.66 $X2=2.92 $Y2=1.22
cc_92 VPB X 0.00690691f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.295
cc_93 N_A_c_105_n N_B_c_187_n 0.0135232f $X=0.505 $Y=1.865 $X2=-0.19 $Y2=-0.245
cc_94 N_A_c_97_n N_B_c_187_n 0.00656481f $X=2.755 $Y=1.195 $X2=-0.19 $Y2=-0.245
cc_95 N_A_c_101_n N_B_c_187_n 0.0202515f $X=0.27 $Y=1.465 $X2=-0.19 $Y2=-0.245
cc_96 N_A_c_94_n N_B_c_188_n 0.0108762f $X=2.89 $Y=1.775 $X2=0 $Y2=0
cc_97 N_A_c_107_n N_B_c_188_n 0.0331104f $X=2.89 $Y=1.865 $X2=0 $Y2=0
cc_98 N_A_c_97_n N_B_c_188_n 0.00424898f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_99 N_A_c_99_n N_B_c_188_n 0.0063017f $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_100 N_A_c_97_n N_B_M1012_g 0.010633f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_101 N_A_c_98_n N_B_M1012_g 0.00124415f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_102 N_A_c_99_n N_B_M1012_g 0.0127642f $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_103 N_A_c_102_n N_B_M1012_g 0.0212043f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_104 N_A_c_94_n N_B_c_190_n 0.00128931f $X=2.89 $Y=1.775 $X2=0 $Y2=0
cc_105 N_A_c_97_n N_B_c_190_n 0.145451f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_106 N_A_c_98_n N_B_c_190_n 0.00662177f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_107 N_A_c_99_n N_B_c_190_n 3.44095e-19 $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_108 N_A_c_101_n N_B_c_190_n 0.00644662f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_109 A N_B_c_190_n 0.0150931f $X=0.24 $Y=1.295 $X2=0 $Y2=0
cc_110 N_A_c_97_n N_C_c_248_n 0.00518557f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_111 N_A_c_97_n N_C_c_249_n 0.0255921f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_112 N_A_c_95_n N_C_c_250_n 0.00317605f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_113 N_A_c_96_n N_C_c_250_n 0.0259948f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_114 N_A_c_97_n N_C_c_250_n 0.0149653f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_115 N_A_c_95_n N_C_c_251_n 0.0170535f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_116 N_A_c_96_n N_C_c_251_n 0.00315685f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_117 N_A_c_97_n N_C_c_251_n 0.0249544f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_118 N_A_c_98_n N_A_302_388#_M1012_d 0.00108111f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_119 N_A_c_94_n N_A_302_388#_c_314_n 0.00281018f $X=2.89 $Y=1.775 $X2=0 $Y2=0
cc_120 N_A_c_107_n N_A_302_388#_c_314_n 0.0224878f $X=2.89 $Y=1.865 $X2=0 $Y2=0
cc_121 N_A_c_98_n N_A_302_388#_M1001_g 3.74191e-19 $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_122 N_A_c_99_n N_A_302_388#_M1001_g 0.0035568f $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_123 N_A_c_102_n N_A_302_388#_M1001_g 0.0249349f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_124 N_A_c_107_n N_A_302_388#_c_326_n 0.0166706f $X=2.89 $Y=1.865 $X2=0 $Y2=0
cc_125 N_A_c_97_n N_A_302_388#_c_326_n 0.00574781f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_126 N_A_c_98_n N_A_302_388#_c_326_n 0.00909601f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_127 N_A_c_99_n N_A_302_388#_c_326_n 0.00134002f $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_128 N_A_c_97_n N_A_302_388#_c_330_n 0.0424115f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_129 N_A_c_97_n N_A_302_388#_c_308_n 0.0243069f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_130 N_A_c_102_n N_A_302_388#_c_309_n 0.00627897f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_131 N_A_c_98_n N_A_302_388#_c_333_n 0.0112121f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_132 N_A_c_99_n N_A_302_388#_c_333_n 9.11899e-19 $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_133 N_A_c_102_n N_A_302_388#_c_333_n 0.00865712f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_134 N_A_c_98_n N_A_302_388#_c_310_n 0.014585f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_135 N_A_c_99_n N_A_302_388#_c_310_n 5.12525e-19 $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_136 N_A_c_102_n N_A_302_388#_c_310_n 0.00373084f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_137 N_A_c_94_n N_A_302_388#_c_311_n 0.00462819f $X=2.89 $Y=1.775 $X2=0 $Y2=0
cc_138 N_A_c_107_n N_A_302_388#_c_311_n 0.00163564f $X=2.89 $Y=1.865 $X2=0 $Y2=0
cc_139 N_A_c_97_n N_A_302_388#_c_341_n 0.0157928f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_140 N_A_c_98_n N_A_302_388#_c_341_n 0.0080232f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_141 N_A_c_99_n N_A_302_388#_c_341_n 4.47709e-19 $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_142 N_A_c_102_n N_A_302_388#_c_341_n 7.14557e-19 $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_143 N_A_c_94_n N_A_302_388#_c_312_n 9.95864e-19 $X=2.89 $Y=1.775 $X2=0 $Y2=0
cc_144 N_A_c_98_n N_A_302_388#_c_312_n 0.0209458f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_145 N_A_c_99_n N_A_302_388#_c_312_n 0.00176886f $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_146 N_A_c_94_n N_A_302_388#_c_313_n 0.00649469f $X=2.89 $Y=1.775 $X2=0 $Y2=0
cc_147 N_A_c_98_n N_A_302_388#_c_313_n 2.43886e-19 $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_148 N_A_c_99_n N_A_302_388#_c_313_n 0.0124829f $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_149 N_A_c_105_n N_VPWR_c_471_n 0.00929585f $X=0.505 $Y=1.865 $X2=0 $Y2=0
cc_150 N_A_c_101_n N_VPWR_c_471_n 0.00182202f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_151 A N_VPWR_c_471_n 0.0148078f $X=0.24 $Y=1.295 $X2=0 $Y2=0
cc_152 N_A_c_107_n N_VPWR_c_472_n 0.00915455f $X=2.89 $Y=1.865 $X2=0 $Y2=0
cc_153 N_A_c_105_n N_VPWR_c_476_n 0.00548284f $X=0.505 $Y=1.865 $X2=0 $Y2=0
cc_154 N_A_c_107_n N_VPWR_c_476_n 0.00548284f $X=2.89 $Y=1.865 $X2=0 $Y2=0
cc_155 N_A_c_105_n N_VPWR_c_469_n 0.00539454f $X=0.505 $Y=1.865 $X2=0 $Y2=0
cc_156 N_A_c_107_n N_VPWR_c_469_n 0.00539454f $X=2.89 $Y=1.865 $X2=0 $Y2=0
cc_157 N_A_c_105_n N_A_116_388#_c_541_n 0.00490148f $X=0.505 $Y=1.865 $X2=0
+ $Y2=0
cc_158 N_A_c_97_n N_A_116_388#_c_541_n 6.30791e-19 $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_159 N_A_c_105_n N_A_116_388#_c_539_n 0.00482252f $X=0.505 $Y=1.865 $X2=0
+ $Y2=0
cc_160 N_A_c_107_n N_A_116_388#_c_544_n 0.00280333f $X=2.89 $Y=1.865 $X2=0 $Y2=0
cc_161 N_A_c_107_n N_A_116_388#_c_540_n 0.00472936f $X=2.89 $Y=1.865 $X2=0 $Y2=0
cc_162 N_A_c_105_n N_A_116_388#_c_546_n 0.00183357f $X=0.505 $Y=1.865 $X2=0
+ $Y2=0
cc_163 N_A_c_98_n N_VGND_M1004_d 5.36408e-19 $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_164 N_A_c_102_n N_VGND_c_673_n 4.07914e-19 $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_165 N_A_c_102_n N_VGND_c_674_n 0.00434272f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_166 N_A_c_102_n N_VGND_c_675_n 0.0030773f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_167 N_A_c_95_n N_VGND_c_679_n 0.0191905f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_168 N_A_c_96_n N_VGND_c_679_n 0.00793088f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A_c_95_n N_VGND_c_685_n 0.012382f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_170 N_A_c_96_n N_VGND_c_685_n 0.00575727f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_171 N_A_c_102_n N_VGND_c_685_n 0.00431597f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_172 N_B_c_190_n N_C_c_246_n 0.0100513f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_173 N_B_c_187_n N_C_c_253_n 0.0371776f $X=0.955 $Y=1.865 $X2=0 $Y2=0
cc_174 N_B_c_190_n N_C_c_253_n 0.00442044f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_175 N_B_c_190_n N_C_c_247_n 0.0103797f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_176 N_B_c_188_n N_C_c_255_n 0.0353468f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_177 N_B_c_190_n N_C_c_255_n 0.00240362f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_178 N_B_M1012_g N_C_c_248_n 0.0303957f $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_179 N_B_c_187_n N_C_c_249_n 0.0266597f $X=0.955 $Y=1.865 $X2=0 $Y2=0
cc_180 N_B_c_188_n N_C_c_249_n 0.0180818f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_181 N_B_M1012_g N_C_c_249_n 0.00483407f $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B_c_190_n N_C_c_249_n 0.0172417f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_183 N_B_M1012_g N_A_302_388#_c_307_n 3.40036e-19 $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_184 N_B_c_188_n N_A_302_388#_c_326_n 0.0149684f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_185 N_B_M1012_g N_A_302_388#_c_330_n 0.0122153f $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_186 N_B_M1012_g N_A_302_388#_c_309_n 0.0022446f $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_187 N_B_c_187_n N_A_302_388#_c_355_n 0.00115622f $X=0.955 $Y=1.865 $X2=0
+ $Y2=0
cc_188 N_B_c_188_n N_A_302_388#_c_355_n 3.66649e-19 $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_189 N_B_c_190_n N_A_302_388#_c_355_n 0.0688717f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_190 N_B_c_190_n N_A_302_388#_c_312_n 0.00244434f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_191 N_B_c_187_n N_VPWR_c_476_n 0.00547215f $X=0.955 $Y=1.865 $X2=0 $Y2=0
cc_192 N_B_c_188_n N_VPWR_c_476_n 0.00547215f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_193 N_B_c_187_n N_VPWR_c_469_n 0.00539454f $X=0.955 $Y=1.865 $X2=0 $Y2=0
cc_194 N_B_c_188_n N_VPWR_c_469_n 0.00539454f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_195 N_B_c_187_n N_A_116_388#_c_541_n 2.09661e-19 $X=0.955 $Y=1.865 $X2=0
+ $Y2=0
cc_196 N_B_c_190_n N_A_116_388#_c_541_n 0.0166452f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_197 N_B_c_187_n N_A_116_388#_c_539_n 0.00457212f $X=0.955 $Y=1.865 $X2=0
+ $Y2=0
cc_198 N_B_c_187_n N_A_116_388#_c_550_n 0.0137656f $X=0.955 $Y=1.865 $X2=0 $Y2=0
cc_199 N_B_c_188_n N_A_116_388#_c_550_n 0.0127563f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_200 N_B_c_190_n N_A_116_388#_c_550_n 0.0166363f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_201 N_B_c_188_n N_A_116_388#_c_540_n 0.00231881f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_202 N_B_c_187_n N_A_206_388#_c_576_n 0.00312019f $X=0.955 $Y=1.865 $X2=0
+ $Y2=0
cc_203 N_B_c_188_n N_A_206_388#_c_576_n 0.0029807f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_204 N_B_M1012_g N_VGND_c_673_n 0.0065526f $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_205 N_B_M1012_g N_VGND_c_674_n 0.00413917f $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_206 N_B_M1012_g N_VGND_c_685_n 0.00399073f $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_207 N_C_c_248_n N_A_302_388#_c_307_n 0.0064141f $X=1.93 $Y=1.185 $X2=0 $Y2=0
cc_208 N_C_c_250_n N_A_302_388#_c_307_n 0.004172f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_209 N_C_c_251_n N_A_302_388#_c_307_n 0.0331922f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_210 N_C_c_255_n N_A_302_388#_c_326_n 0.00857129f $X=1.885 $Y=1.865 $X2=0
+ $Y2=0
cc_211 N_C_c_248_n N_A_302_388#_c_330_n 0.00871095f $X=1.93 $Y=1.185 $X2=0 $Y2=0
cc_212 N_C_c_248_n N_A_302_388#_c_308_n 7.15561e-19 $X=1.93 $Y=1.185 $X2=0 $Y2=0
cc_213 N_C_c_249_n N_A_302_388#_c_308_n 0.00114784f $X=1.885 $Y=1.345 $X2=0
+ $Y2=0
cc_214 N_C_c_250_n N_A_302_388#_c_308_n 0.00179824f $X=1.215 $Y=0.435 $X2=0
+ $Y2=0
cc_215 N_C_c_251_n N_A_302_388#_c_308_n 0.0143345f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_216 N_C_c_253_n N_A_302_388#_c_355_n 0.00519335f $X=1.435 $Y=1.865 $X2=0
+ $Y2=0
cc_217 N_C_c_255_n N_A_302_388#_c_355_n 0.00209181f $X=1.885 $Y=1.865 $X2=0
+ $Y2=0
cc_218 N_C_c_249_n N_A_302_388#_c_355_n 3.55714e-19 $X=1.885 $Y=1.345 $X2=0
+ $Y2=0
cc_219 N_C_c_253_n N_VPWR_c_476_n 0.00401361f $X=1.435 $Y=1.865 $X2=0 $Y2=0
cc_220 N_C_c_255_n N_VPWR_c_476_n 0.00401361f $X=1.885 $Y=1.865 $X2=0 $Y2=0
cc_221 N_C_c_253_n N_VPWR_c_469_n 0.00539454f $X=1.435 $Y=1.865 $X2=0 $Y2=0
cc_222 N_C_c_255_n N_VPWR_c_469_n 0.00539454f $X=1.885 $Y=1.865 $X2=0 $Y2=0
cc_223 N_C_c_253_n N_A_116_388#_c_550_n 0.0126399f $X=1.435 $Y=1.865 $X2=0 $Y2=0
cc_224 N_C_c_255_n N_A_116_388#_c_550_n 0.0113838f $X=1.885 $Y=1.865 $X2=0 $Y2=0
cc_225 N_C_c_253_n N_A_206_388#_c_576_n 0.010492f $X=1.435 $Y=1.865 $X2=0 $Y2=0
cc_226 N_C_c_255_n N_A_206_388#_c_576_n 0.0105055f $X=1.885 $Y=1.865 $X2=0 $Y2=0
cc_227 N_C_c_248_n N_VGND_c_673_n 0.00349022f $X=1.93 $Y=1.185 $X2=0 $Y2=0
cc_228 N_C_c_251_n N_VGND_c_673_n 0.00220313f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_229 N_C_c_248_n N_VGND_c_679_n 0.00434272f $X=1.93 $Y=1.185 $X2=0 $Y2=0
cc_230 N_C_c_250_n N_VGND_c_679_n 0.00637453f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_231 N_C_c_251_n N_VGND_c_679_n 0.0203268f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_232 N_C_c_248_n N_VGND_c_685_n 0.00436049f $X=1.93 $Y=1.185 $X2=0 $Y2=0
cc_233 N_C_c_250_n N_VGND_c_685_n 0.00418281f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_234 N_C_c_251_n N_VGND_c_685_n 0.0124484f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_235 N_A_302_388#_c_326_n N_VPWR_M1006_s 0.00966885f $X=3.225 $Y=2.035 $X2=0
+ $Y2=0
cc_236 N_A_302_388#_c_311_n N_VPWR_M1006_s 0.00135024f $X=3.31 $Y=1.95 $X2=0
+ $Y2=0
cc_237 N_A_302_388#_c_314_n N_VPWR_c_472_n 0.0111999f $X=3.425 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_A_302_388#_c_315_n N_VPWR_c_472_n 5.35985e-19 $X=3.875 $Y=1.765 $X2=0
+ $Y2=0
cc_239 N_A_302_388#_c_326_n N_VPWR_c_472_n 0.022569f $X=3.225 $Y=2.035 $X2=0
+ $Y2=0
cc_240 N_A_302_388#_c_314_n N_VPWR_c_473_n 5.83721e-19 $X=3.425 $Y=1.765 $X2=0
+ $Y2=0
cc_241 N_A_302_388#_c_315_n N_VPWR_c_473_n 0.0133451f $X=3.875 $Y=1.765 $X2=0
+ $Y2=0
cc_242 N_A_302_388#_c_316_n N_VPWR_c_473_n 0.00630489f $X=4.325 $Y=1.765 $X2=0
+ $Y2=0
cc_243 N_A_302_388#_c_317_n N_VPWR_c_475_n 0.00993564f $X=4.775 $Y=1.765 $X2=0
+ $Y2=0
cc_244 N_A_302_388#_c_314_n N_VPWR_c_477_n 0.00413917f $X=3.425 $Y=1.765 $X2=0
+ $Y2=0
cc_245 N_A_302_388#_c_315_n N_VPWR_c_477_n 0.00413917f $X=3.875 $Y=1.765 $X2=0
+ $Y2=0
cc_246 N_A_302_388#_c_316_n N_VPWR_c_478_n 0.00445602f $X=4.325 $Y=1.765 $X2=0
+ $Y2=0
cc_247 N_A_302_388#_c_317_n N_VPWR_c_478_n 0.00445602f $X=4.775 $Y=1.765 $X2=0
+ $Y2=0
cc_248 N_A_302_388#_c_314_n N_VPWR_c_469_n 0.00817726f $X=3.425 $Y=1.765 $X2=0
+ $Y2=0
cc_249 N_A_302_388#_c_315_n N_VPWR_c_469_n 0.00817726f $X=3.875 $Y=1.765 $X2=0
+ $Y2=0
cc_250 N_A_302_388#_c_316_n N_VPWR_c_469_n 0.00857589f $X=4.325 $Y=1.765 $X2=0
+ $Y2=0
cc_251 N_A_302_388#_c_317_n N_VPWR_c_469_n 0.00861084f $X=4.775 $Y=1.765 $X2=0
+ $Y2=0
cc_252 N_A_302_388#_c_326_n N_A_116_388#_M1003_d 0.00713316f $X=3.225 $Y=2.035
+ $X2=0 $Y2=0
cc_253 N_A_302_388#_M1013_d N_A_116_388#_c_550_n 0.00392879f $X=1.51 $Y=1.94
+ $X2=0 $Y2=0
cc_254 N_A_302_388#_c_326_n N_A_116_388#_c_550_n 0.0273439f $X=3.225 $Y=2.035
+ $X2=0 $Y2=0
cc_255 N_A_302_388#_c_355_n N_A_116_388#_c_550_n 0.015935f $X=1.825 $Y=2.075
+ $X2=0 $Y2=0
cc_256 N_A_302_388#_c_326_n N_A_116_388#_c_544_n 0.0202766f $X=3.225 $Y=2.035
+ $X2=0 $Y2=0
cc_257 N_A_302_388#_c_326_n N_A_206_388#_M1016_s 0.00551997f $X=3.225 $Y=2.035
+ $X2=0 $Y2=0
cc_258 N_A_302_388#_M1013_d N_A_206_388#_c_576_n 0.00200574f $X=1.51 $Y=1.94
+ $X2=0 $Y2=0
cc_259 N_A_302_388#_M1001_g N_X_c_590_n 0.00492137f $X=3.43 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A_302_388#_M1007_g N_X_c_590_n 3.97599e-19 $X=3.865 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_302_388#_c_333_n N_X_c_590_n 0.0133617f $X=3.225 $Y=0.855 $X2=0 $Y2=0
cc_262 N_A_302_388#_c_310_n N_X_c_590_n 0.00133388f $X=3.31 $Y=1.3 $X2=0 $Y2=0
cc_263 N_A_302_388#_c_314_n N_X_c_597_n 0.0061914f $X=3.425 $Y=1.765 $X2=0 $Y2=0
cc_264 N_A_302_388#_c_315_n N_X_c_597_n 0.00438646f $X=3.875 $Y=1.765 $X2=0
+ $Y2=0
cc_265 N_A_302_388#_c_326_n N_X_c_597_n 0.0117532f $X=3.225 $Y=2.035 $X2=0 $Y2=0
cc_266 N_A_302_388#_M1007_g N_X_c_591_n 0.0127819f $X=3.865 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A_302_388#_M1009_g N_X_c_591_n 0.0113778f $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A_302_388#_c_404_p N_X_c_591_n 0.0492576f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_269 N_A_302_388#_c_313_n N_X_c_591_n 0.00358729f $X=4.775 $Y=1.532 $X2=0
+ $Y2=0
cc_270 N_A_302_388#_M1001_g N_X_c_592_n 7.34064e-19 $X=3.43 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A_302_388#_c_310_n N_X_c_592_n 0.0134529f $X=3.31 $Y=1.3 $X2=0 $Y2=0
cc_272 N_A_302_388#_c_404_p N_X_c_592_n 0.014338f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_273 N_A_302_388#_c_313_n N_X_c_592_n 0.00244604f $X=4.775 $Y=1.532 $X2=0
+ $Y2=0
cc_274 N_A_302_388#_c_315_n N_X_c_598_n 0.0130724f $X=3.875 $Y=1.765 $X2=0 $Y2=0
cc_275 N_A_302_388#_c_316_n N_X_c_598_n 0.0119563f $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_276 N_A_302_388#_c_404_p N_X_c_598_n 0.0477127f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_277 N_A_302_388#_c_313_n N_X_c_598_n 0.00919355f $X=4.775 $Y=1.532 $X2=0
+ $Y2=0
cc_278 N_A_302_388#_c_314_n N_X_c_599_n 8.17608e-19 $X=3.425 $Y=1.765 $X2=0
+ $Y2=0
cc_279 N_A_302_388#_c_326_n N_X_c_599_n 0.00174806f $X=3.225 $Y=2.035 $X2=0
+ $Y2=0
cc_280 N_A_302_388#_c_311_n N_X_c_599_n 0.0118751f $X=3.31 $Y=1.95 $X2=0 $Y2=0
cc_281 N_A_302_388#_c_404_p N_X_c_599_n 0.0143367f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_282 N_A_302_388#_c_313_n N_X_c_599_n 0.00421663f $X=4.775 $Y=1.532 $X2=0
+ $Y2=0
cc_283 N_A_302_388#_c_315_n N_X_c_600_n 7.68526e-19 $X=3.875 $Y=1.765 $X2=0
+ $Y2=0
cc_284 N_A_302_388#_c_316_n N_X_c_600_n 0.012705f $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_285 N_A_302_388#_c_317_n N_X_c_600_n 0.017229f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_286 N_A_302_388#_M1007_g N_X_c_593_n 7.04495e-19 $X=3.865 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A_302_388#_M1009_g N_X_c_593_n 0.00953543f $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_288 N_A_302_388#_M1015_g N_X_c_593_n 3.97481e-19 $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_289 N_A_302_388#_M1015_g N_X_c_594_n 0.0160474f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_290 N_A_302_388#_c_404_p N_X_c_594_n 0.00221753f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_291 N_A_302_388#_c_317_n N_X_c_601_n 0.0152503f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_292 N_A_302_388#_c_313_n N_X_c_601_n 5.4426e-19 $X=4.775 $Y=1.532 $X2=0 $Y2=0
cc_293 N_A_302_388#_c_316_n N_X_c_602_n 9.3899e-19 $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_294 N_A_302_388#_c_317_n N_X_c_602_n 0.00114764f $X=4.775 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A_302_388#_c_404_p N_X_c_602_n 0.0252322f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_296 N_A_302_388#_c_313_n N_X_c_602_n 0.00805362f $X=4.775 $Y=1.532 $X2=0
+ $Y2=0
cc_297 N_A_302_388#_M1009_g N_X_c_595_n 9.7541e-19 $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_298 N_A_302_388#_c_404_p N_X_c_595_n 0.0209731f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_299 N_A_302_388#_c_313_n N_X_c_595_n 0.00232957f $X=4.775 $Y=1.532 $X2=0
+ $Y2=0
cc_300 N_A_302_388#_c_317_n X 0.00133808f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_301 N_A_302_388#_M1015_g X 0.0067245f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_302 N_A_302_388#_c_404_p X 0.0206535f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_303 N_A_302_388#_c_313_n X 0.0158588f $X=4.775 $Y=1.532 $X2=0 $Y2=0
cc_304 N_A_302_388#_c_330_n N_VGND_M1008_d 0.00507735f $X=2.55 $Y=0.855
+ $X2=-0.19 $Y2=-0.245
cc_305 N_A_302_388#_c_333_n N_VGND_M1004_d 0.00807426f $X=3.225 $Y=0.855 $X2=0
+ $Y2=0
cc_306 N_A_302_388#_c_310_n N_VGND_M1004_d 0.00203236f $X=3.31 $Y=1.3 $X2=0
+ $Y2=0
cc_307 N_A_302_388#_c_307_n N_VGND_c_673_n 0.0101711f $X=1.715 $Y=0.515 $X2=0
+ $Y2=0
cc_308 N_A_302_388#_c_330_n N_VGND_c_673_n 0.0204503f $X=2.55 $Y=0.855 $X2=0
+ $Y2=0
cc_309 N_A_302_388#_c_309_n N_VGND_c_673_n 0.0101711f $X=2.715 $Y=0.515 $X2=0
+ $Y2=0
cc_310 N_A_302_388#_c_309_n N_VGND_c_674_n 0.014415f $X=2.715 $Y=0.515 $X2=0
+ $Y2=0
cc_311 N_A_302_388#_M1001_g N_VGND_c_675_n 0.00690871f $X=3.43 $Y=0.74 $X2=0
+ $Y2=0
cc_312 N_A_302_388#_M1007_g N_VGND_c_675_n 4.02157e-19 $X=3.865 $Y=0.74 $X2=0
+ $Y2=0
cc_313 N_A_302_388#_c_309_n N_VGND_c_675_n 0.0101711f $X=2.715 $Y=0.515 $X2=0
+ $Y2=0
cc_314 N_A_302_388#_c_333_n N_VGND_c_675_n 0.0211625f $X=3.225 $Y=0.855 $X2=0
+ $Y2=0
cc_315 N_A_302_388#_M1001_g N_VGND_c_676_n 4.57455e-19 $X=3.43 $Y=0.74 $X2=0
+ $Y2=0
cc_316 N_A_302_388#_M1007_g N_VGND_c_676_n 0.00897549f $X=3.865 $Y=0.74 $X2=0
+ $Y2=0
cc_317 N_A_302_388#_M1009_g N_VGND_c_676_n 0.00497505f $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_318 N_A_302_388#_M1009_g N_VGND_c_678_n 5.12327e-19 $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_319 N_A_302_388#_M1015_g N_VGND_c_678_n 0.0110492f $X=4.785 $Y=0.74 $X2=0
+ $Y2=0
cc_320 N_A_302_388#_c_307_n N_VGND_c_679_n 0.014415f $X=1.715 $Y=0.515 $X2=0
+ $Y2=0
cc_321 N_A_302_388#_M1001_g N_VGND_c_680_n 0.00383152f $X=3.43 $Y=0.74 $X2=0
+ $Y2=0
cc_322 N_A_302_388#_M1007_g N_VGND_c_680_n 0.00383152f $X=3.865 $Y=0.74 $X2=0
+ $Y2=0
cc_323 N_A_302_388#_M1009_g N_VGND_c_681_n 0.00434272f $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_324 N_A_302_388#_M1015_g N_VGND_c_681_n 0.00383152f $X=4.785 $Y=0.74 $X2=0
+ $Y2=0
cc_325 N_A_302_388#_M1001_g N_VGND_c_685_n 0.00708259f $X=3.43 $Y=0.74 $X2=0
+ $Y2=0
cc_326 N_A_302_388#_M1007_g N_VGND_c_685_n 0.0075759f $X=3.865 $Y=0.74 $X2=0
+ $Y2=0
cc_327 N_A_302_388#_M1009_g N_VGND_c_685_n 0.00821839f $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_328 N_A_302_388#_M1015_g N_VGND_c_685_n 0.0075754f $X=4.785 $Y=0.74 $X2=0
+ $Y2=0
cc_329 N_A_302_388#_c_307_n N_VGND_c_685_n 0.0119404f $X=1.715 $Y=0.515 $X2=0
+ $Y2=0
cc_330 N_A_302_388#_c_330_n N_VGND_c_685_n 0.0118074f $X=2.55 $Y=0.855 $X2=0
+ $Y2=0
cc_331 N_A_302_388#_c_309_n N_VGND_c_685_n 0.0119404f $X=2.715 $Y=0.515 $X2=0
+ $Y2=0
cc_332 N_A_302_388#_c_333_n N_VGND_c_685_n 0.00714277f $X=3.225 $Y=0.855 $X2=0
+ $Y2=0
cc_333 N_VPWR_c_471_n N_A_116_388#_c_541_n 0.0275535f $X=0.28 $Y=2.085 $X2=0
+ $Y2=0
cc_334 N_VPWR_c_471_n N_A_116_388#_c_539_n 0.0275831f $X=0.28 $Y=2.085 $X2=0
+ $Y2=0
cc_335 N_VPWR_c_476_n N_A_116_388#_c_539_n 0.0102021f $X=3.035 $Y=3.33 $X2=0
+ $Y2=0
cc_336 N_VPWR_c_469_n N_A_116_388#_c_539_n 0.00903636f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_337 N_VPWR_c_469_n N_A_116_388#_c_550_n 0.0142759f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_472_n N_A_116_388#_c_544_n 0.017515f $X=3.2 $Y=2.455 $X2=0 $Y2=0
cc_339 N_VPWR_c_472_n N_A_116_388#_c_540_n 0.0282274f $X=3.2 $Y=2.455 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_476_n N_A_116_388#_c_540_n 0.0134917f $X=3.035 $Y=3.33 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_469_n N_A_116_388#_c_540_n 0.0119489f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_471_n N_A_116_388#_c_546_n 0.0121024f $X=0.28 $Y=2.085 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_476_n N_A_206_388#_c_576_n 0.049596f $X=3.035 $Y=3.33 $X2=0
+ $Y2=0
cc_344 N_VPWR_c_469_n N_A_206_388#_c_576_n 0.0461161f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_472_n N_X_c_597_n 0.0449718f $X=3.2 $Y=2.455 $X2=0 $Y2=0
cc_346 N_VPWR_c_473_n N_X_c_597_n 0.0535896f $X=4.1 $Y=2.305 $X2=0 $Y2=0
cc_347 N_VPWR_c_477_n N_X_c_597_n 0.00749631f $X=3.935 $Y=3.33 $X2=0 $Y2=0
cc_348 N_VPWR_c_469_n N_X_c_597_n 0.0062048f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_349 N_VPWR_M1010_s N_X_c_598_n 0.00222494f $X=3.95 $Y=1.84 $X2=0 $Y2=0
cc_350 N_VPWR_c_473_n N_X_c_598_n 0.0154248f $X=4.1 $Y=2.305 $X2=0 $Y2=0
cc_351 N_VPWR_c_473_n N_X_c_600_n 0.0563525f $X=4.1 $Y=2.305 $X2=0 $Y2=0
cc_352 N_VPWR_c_475_n N_X_c_600_n 0.0563525f $X=5 $Y=2.305 $X2=0 $Y2=0
cc_353 N_VPWR_c_478_n N_X_c_600_n 0.014552f $X=4.915 $Y=3.33 $X2=0 $Y2=0
cc_354 N_VPWR_c_469_n N_X_c_600_n 0.0119791f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_355 N_VPWR_M1014_s N_X_c_601_n 0.0036905f $X=4.85 $Y=1.84 $X2=0 $Y2=0
cc_356 N_VPWR_c_475_n N_X_c_601_n 0.0214215f $X=5 $Y=2.305 $X2=0 $Y2=0
cc_357 N_A_116_388#_c_550_n N_A_206_388#_M1000_s 0.00639049f $X=2.5 $Y=2.455
+ $X2=-0.19 $Y2=1.66
cc_358 N_A_116_388#_c_550_n N_A_206_388#_M1016_s 0.0055195f $X=2.5 $Y=2.455
+ $X2=0 $Y2=0
cc_359 N_A_116_388#_c_539_n N_A_206_388#_c_576_n 0.0176833f $X=0.73 $Y=2.795
+ $X2=0 $Y2=0
cc_360 N_A_116_388#_c_550_n N_A_206_388#_c_576_n 0.0689258f $X=2.5 $Y=2.455
+ $X2=0 $Y2=0
cc_361 N_A_116_388#_c_540_n N_A_206_388#_c_576_n 0.0111988f $X=2.665 $Y=2.795
+ $X2=0 $Y2=0
cc_362 N_X_c_591_n N_VGND_M1007_s 0.00402642f $X=4.405 $Y=1.045 $X2=0 $Y2=0
cc_363 N_X_c_594_n N_VGND_M1015_s 0.00338075f $X=4.925 $Y=1.045 $X2=0 $Y2=0
cc_364 N_X_c_590_n N_VGND_c_675_n 0.0173183f $X=3.65 $Y=0.515 $X2=0 $Y2=0
cc_365 N_X_c_590_n N_VGND_c_676_n 0.0157999f $X=3.65 $Y=0.515 $X2=0 $Y2=0
cc_366 N_X_c_591_n N_VGND_c_676_n 0.0154151f $X=4.405 $Y=1.045 $X2=0 $Y2=0
cc_367 N_X_c_593_n N_VGND_c_676_n 0.0251662f $X=4.57 $Y=0.515 $X2=0 $Y2=0
cc_368 N_X_c_593_n N_VGND_c_678_n 0.0164981f $X=4.57 $Y=0.515 $X2=0 $Y2=0
cc_369 N_X_c_594_n N_VGND_c_678_n 0.023173f $X=4.925 $Y=1.045 $X2=0 $Y2=0
cc_370 N_X_c_590_n N_VGND_c_680_n 0.00749631f $X=3.65 $Y=0.515 $X2=0 $Y2=0
cc_371 N_X_c_593_n N_VGND_c_681_n 0.0109942f $X=4.57 $Y=0.515 $X2=0 $Y2=0
cc_372 N_X_c_590_n N_VGND_c_685_n 0.0062048f $X=3.65 $Y=0.515 $X2=0 $Y2=0
cc_373 N_X_c_593_n N_VGND_c_685_n 0.00904371f $X=4.57 $Y=0.515 $X2=0 $Y2=0
