* File: sky130_fd_sc_ls__o2111a_2.spice
* Created: Wed Sep  2 11:16:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o2111a_2.pex.spice"
.subckt sky130_fd_sc_ls__o2111a_2  VNB VPB A1 A2 B1 C1 D1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D1	D1
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A1_M1008_g N_A_54_74#_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.2627 PD=1.16 PS=2.19 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1000 N_A_54_74#_M1000_d N_A2_M1000_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1554 PD=1.09 PS=1.16 NRD=11.34 NRS=11.34 M=1 R=4.93333
+ SA=75000.8 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1012 A_369_74# N_B1_M1012_g N_A_54_74#_M1000_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1147 AS=0.1295 PD=1.05 PS=1.09 NRD=16.212 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1005 A_461_74# N_C1_M1005_g A_369_74# VNB NSHORT L=0.15 W=0.74 AD=0.1554
+ AS=0.1147 PD=1.16 PS=1.05 NRD=25.128 NRS=16.212 M=1 R=4.93333 SA=75001.8
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1010 N_A_236_368#_M1010_d N_D1_M1010_g A_461_74# VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75002.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A_236_368#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A_236_368#_M1011_g N_X_M1001_s VNB NSHORT L=0.15 W=0.74
+ AD=0.222 AS=0.1036 PD=2.08 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 A_152_368# N_A1_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75003.8 A=0.15 P=2.3 MULT=1
MM1013 N_A_236_368#_M1013_d N_A2_M1013_g A_152_368# VPB PHIGHVT L=0.15 W=1
+ AD=0.21 AS=0.135 PD=1.42 PS=1.27 NRD=25.5903 NRS=15.7403 M=1 R=6.66667
+ SA=75000.6 SB=75003.4 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_B1_M1009_g N_A_236_368#_M1013_d VPB PHIGHVT L=0.15 W=1
+ AD=0.245 AS=0.21 PD=1.49 PS=1.42 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75001.2 SB=75002.8 A=0.15 P=2.3 MULT=1
MM1004 N_A_236_368#_M1004_d N_C1_M1004_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.245 PD=1.35 PS=1.49 NRD=1.9503 NRS=29.55 M=1 R=6.66667
+ SA=75001.8 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_D1_M1007_g N_A_236_368#_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.406509 AS=0.175 PD=1.83962 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75002.3 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1003 N_X_M1003_d N_A_236_368#_M1003_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.455291 PD=1.42 PS=2.06038 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1006 N_X_M1003_d N_A_236_368#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.4 SB=75000.3 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ls__o2111a_2.pxi.spice"
*
.ends
*
*
