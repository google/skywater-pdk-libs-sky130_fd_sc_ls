* File: sky130_fd_sc_ls__ha_2.spice
* Created: Fri Aug 28 13:27:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__ha_2.pex.spice"
.subckt sky130_fd_sc_ls__ha_2  VNB VPB B A VPWR SUM COUT VGND
* 
* VGND	VGND
* COUT	COUT
* SUM	SUM
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1013 A_114_74# N_B_M1013_g N_A_27_74#_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_M1010_g A_114_74# VNB NSHORT L=0.15 W=0.74 AD=0.1036
+ AS=0.0888 PD=1.02 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6 SB=75001
+ A=0.111 P=1.78 MULT=1
MM1000 N_A_278_74#_M1000_d N_A_M1000_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_B_M1009_g N_A_278_74#_M1000_d VNB NSHORT L=0.15 W=0.74
+ AD=0.19515 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_A_278_74#_M1015_d N_A_27_74#_M1015_g N_A_391_388#_M1015_s VNB NSHORT
+ L=0.15 W=0.74 AD=0.2011 AS=0.201625 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_SUM_M1003_d N_A_391_388#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1221 AS=0.1962 PD=1.07 PS=2.05 NRD=4.044 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1012 N_SUM_M1003_d N_A_391_388#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1221 AS=0.1036 PD=1.07 PS=1.02 NRD=4.044 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1012_s N_A_27_74#_M1008_g N_COUT_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A_27_74#_M1017_g N_COUT_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_27_74#_M1005_d N_B_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75004.9 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_27_74#_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.17925 AS=0.15 PD=1.375 PS=1.3 NRD=6.8753 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75004.4 A=0.15 P=2.3 MULT=1
MM1002 A_307_388# N_A_M1002_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.17925 PD=1.27 PS=1.375 NRD=15.7403 NRS=7.8603 M=1 R=6.66667 SA=75001.2
+ SB=75004 A=0.15 P=2.3 MULT=1
MM1016 N_A_391_388#_M1016_d N_B_M1016_g A_307_388# VPB PHIGHVT L=0.15 W=1
+ AD=0.495 AS=0.135 PD=1.99 PS=1.27 NRD=137.88 NRS=15.7403 M=1 R=6.66667
+ SA=75001.6 SB=75003.6 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_A_27_74#_M1011_g N_A_391_388#_M1016_d VPB PHIGHVT L=0.15
+ W=1 AD=0.364953 AS=0.495 PD=1.75 PS=1.99 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75002.7 SB=75002.5 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1011_d N_A_391_388#_M1001_g N_SUM_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.408747 AS=0.168 PD=1.96 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75003.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1014_d N_A_391_388#_M1014_g N_SUM_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1004 N_COUT_M1004_d N_A_27_74#_M1004_g N_VPWR_M1014_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1007 N_COUT_M1004_d N_A_27_74#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ls__ha_2.pxi.spice"
*
.ends
*
*
