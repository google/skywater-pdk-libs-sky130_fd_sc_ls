* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__ha_1 A B VGND VNB VPB VPWR COUT SUM
X0 VPWR B a_239_294# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 a_83_260# a_239_294# a_305_130# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 a_239_294# B a_695_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 VPWR a_239_294# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X4 a_386_392# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_305_130# B VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 SUM a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 VGND a_239_294# COUT VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 a_239_294# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X9 VPWR a_239_294# a_83_260# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 VGND A a_305_130# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 SUM a_83_260# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 a_83_260# B a_386_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_695_119# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
