* File: sky130_fd_sc_ls__and4_4.spice
* Created: Fri Aug 28 13:05:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__and4_4.pex.spice"
.subckt sky130_fd_sc_ls__and4_4  VNB VPB A B D C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* D	D
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_A_119_119#_M1002_d N_B_M1002_g N_A_32_119#_M1002_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75003.4 A=0.096 P=1.58 MULT=1
MM1001 N_A_116_392#_M1001_d N_A_M1001_g N_A_119_119#_M1002_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1003 N_A_116_392#_M1001_d N_A_M1003_g N_A_119_119#_M1003_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1016 N_A_119_119#_M1003_s N_B_M1016_g N_A_32_119#_M1016_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1019 N_A_463_119#_M1019_d N_C_M1019_g N_A_32_119#_M1016_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.9 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1012 N_VGND_M1012_d N_D_M1012_g N_A_463_119#_M1019_d VNB NSHORT L=0.15 W=0.64
+ AD=0.170525 AS=0.0896 PD=1.285 PS=0.92 NRD=39.636 NRS=0 M=1 R=4.26667
+ SA=75002.4 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1018 N_VGND_M1012_d N_D_M1018_g N_A_463_119#_M1018_s VNB NSHORT L=0.15 W=0.64
+ AD=0.170525 AS=0.0896 PD=1.285 PS=0.92 NRD=39.636 NRS=0 M=1 R=4.26667
+ SA=75002.9 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1020 N_A_463_119#_M1018_s N_C_M1020_g N_A_32_119#_M1020_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1705 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75003.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1007_d N_A_116_392#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2405 AS=0.1147 PD=2.13 PS=1.05 NRD=6.48 NRS=4.86 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_116_392#_M1013_g N_X_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1147 PD=1.09 PS=1.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1013_d N_A_116_392#_M1021_g N_X_M1021_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1022_d N_A_116_392#_M1022_g N_X_M1021_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2146 AS=0.1036 PD=2.06 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_A_116_392#_M1017_d N_B_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75005.9 A=0.15 P=2.3 MULT=1
MM1000 N_A_116_392#_M1017_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.7
+ SB=75005.5 A=0.15 P=2.3 MULT=1
MM1015 N_A_116_392#_M1015_d N_A_M1015_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1575 AS=0.15 PD=1.315 PS=1.3 NRD=4.9053 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75005 A=0.15 P=2.3 MULT=1
MM1023 N_A_116_392#_M1015_d N_B_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1
+ AD=0.1575 AS=0.175 PD=1.315 PS=1.35 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.6 SB=75004.6 A=0.15 P=2.3 MULT=1
MM1006 N_A_116_392#_M1006_d N_C_M1006_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75002.1 SB=75004.1 A=0.15 P=2.3 MULT=1
MM1004 N_A_116_392#_M1006_d N_D_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.3675 PD=1.3 PS=1.735 NRD=1.9503 NRS=2.9353 M=1 R=6.66667
+ SA=75002.5 SB=75003.6 A=0.15 P=2.3 MULT=1
MM1010 N_A_116_392#_M1010_d N_D_M1010_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.3675 PD=1.35 PS=1.735 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75003.4 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1009 N_A_116_392#_M1010_d N_C_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.208396 PD=1.35 PS=1.4434 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75003.9 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1005_d N_A_116_392#_M1005_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.233404 PD=1.47 PS=1.6166 NRD=10.5395 NRS=12.2928 M=1 R=7.46667
+ SA=75004 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1008 N_X_M1005_d N_A_116_392#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.5 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1011 N_X_M1011_d N_A_116_392#_M1011_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75005
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1014 N_X_M1011_d N_A_116_392#_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75005.4 SB=75000.3 A=0.168 P=2.54 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.206 P=17.92
c_70 VNB 0 4.03451e-19 $X=0 $Y=0
c_131 VPB 0 8.82342e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__and4_4.pxi.spice"
*
.ends
*
*
