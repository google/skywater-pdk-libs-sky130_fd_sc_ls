* File: sky130_fd_sc_ls__sedfxbp_1.pxi.spice
* Created: Fri Aug 28 14:06:51 2020
* 
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%D N_D_c_337_n N_D_c_342_n N_D_c_343_n
+ N_D_M1023_g N_D_M1013_g N_D_c_339_n D D N_D_c_340_n N_D_c_341_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_1%D
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%A_161_394# N_A_161_394#_M1012_s
+ N_A_161_394#_M1019_s N_A_161_394#_c_387_n N_A_161_394#_M1029_g
+ N_A_161_394#_M1009_g N_A_161_394#_c_388_n N_A_161_394#_c_380_n
+ N_A_161_394#_c_381_n N_A_161_394#_c_382_n N_A_161_394#_c_383_n
+ N_A_161_394#_c_390_n N_A_161_394#_c_391_n N_A_161_394#_c_384_n
+ N_A_161_394#_c_392_n N_A_161_394#_c_393_n N_A_161_394#_c_385_n
+ N_A_161_394#_c_386_n N_A_161_394#_c_396_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_1%A_161_394#
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%DE N_DE_M1014_g N_DE_c_492_n N_DE_c_493_n
+ N_DE_c_499_n N_DE_c_500_n N_DE_M1019_g N_DE_c_494_n N_DE_M1012_g N_DE_c_501_n
+ N_DE_c_502_n N_DE_M1020_g N_DE_c_495_n N_DE_c_503_n DE N_DE_c_496_n
+ N_DE_c_497_n N_DE_c_498_n PM_SKY130_FD_SC_LS__SEDFXBP_1%DE
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%A_575_305# N_A_575_305#_M1028_d
+ N_A_575_305#_M1002_d N_A_575_305#_M1001_g N_A_575_305#_c_594_n
+ N_A_575_305#_c_595_n N_A_575_305#_M1011_g N_A_575_305#_c_578_n
+ N_A_575_305#_M1032_g N_A_575_305#_c_579_n N_A_575_305#_c_580_n
+ N_A_575_305#_c_596_n N_A_575_305#_M1039_g N_A_575_305#_c_581_n
+ N_A_575_305#_c_582_n N_A_575_305#_M1040_g N_A_575_305#_M1000_g
+ N_A_575_305#_c_584_n N_A_575_305#_c_585_n N_A_575_305#_c_600_n
+ N_A_575_305#_c_586_n N_A_575_305#_c_587_n N_A_575_305#_c_588_n
+ N_A_575_305#_c_589_n N_A_575_305#_c_590_n N_A_575_305#_c_591_n
+ N_A_575_305#_c_601_n N_A_575_305#_c_602_n N_A_575_305#_c_603_n
+ N_A_575_305#_c_592_n N_A_575_305#_c_593_n N_A_575_305#_c_606_n
+ N_A_575_305#_c_607_n PM_SKY130_FD_SC_LS__SEDFXBP_1%A_575_305#
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%A_667_87# N_A_667_87#_M1037_s
+ N_A_667_87#_M1003_s N_A_667_87#_c_836_n N_A_667_87#_M1026_g
+ N_A_667_87#_c_837_n N_A_667_87#_c_838_n N_A_667_87#_c_843_n
+ N_A_667_87#_M1007_g N_A_667_87#_c_839_n N_A_667_87#_c_867_p
+ N_A_667_87#_c_840_n N_A_667_87#_c_845_n N_A_667_87#_c_846_n
+ N_A_667_87#_c_841_n N_A_667_87#_c_842_n N_A_667_87#_c_847_n
+ N_A_667_87#_c_848_n N_A_667_87#_c_849_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_1%A_667_87#
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%SCD N_SCD_c_927_n N_SCD_c_932_n N_SCD_M1033_g
+ N_SCD_M1024_g SCD N_SCD_c_930_n PM_SKY130_FD_SC_LS__SEDFXBP_1%SCD
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%SCE N_SCE_c_978_n N_SCE_M1021_g N_SCE_c_979_n
+ N_SCE_c_980_n N_SCE_c_981_n N_SCE_c_982_n N_SCE_M1003_g N_SCE_M1037_g
+ N_SCE_c_973_n N_SCE_c_974_n N_SCE_M1010_g SCE N_SCE_c_976_n N_SCE_c_977_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_1%SCE
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%CLK N_CLK_c_1052_n N_CLK_M1034_g N_CLK_c_1053_n
+ N_CLK_M1015_g CLK PM_SKY130_FD_SC_LS__SEDFXBP_1%CLK
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%A_1549_74# N_A_1549_74#_M1004_d
+ N_A_1549_74#_M1008_d N_A_1549_74#_c_1111_n N_A_1549_74#_M1017_g
+ N_A_1549_74#_M1043_g N_A_1549_74#_M1018_g N_A_1549_74#_c_1112_n
+ N_A_1549_74#_c_1113_n N_A_1549_74#_c_1114_n N_A_1549_74#_M1006_g
+ N_A_1549_74#_c_1088_n N_A_1549_74#_c_1089_n N_A_1549_74#_c_1090_n
+ N_A_1549_74#_c_1091_n N_A_1549_74#_c_1116_n N_A_1549_74#_c_1092_n
+ N_A_1549_74#_c_1093_n N_A_1549_74#_c_1094_n N_A_1549_74#_c_1184_p
+ N_A_1549_74#_c_1095_n N_A_1549_74#_c_1096_n N_A_1549_74#_c_1097_n
+ N_A_1549_74#_c_1098_n N_A_1549_74#_c_1099_n N_A_1549_74#_c_1100_n
+ N_A_1549_74#_c_1101_n N_A_1549_74#_c_1102_n N_A_1549_74#_c_1103_n
+ N_A_1549_74#_c_1119_n N_A_1549_74#_c_1104_n N_A_1549_74#_c_1105_n
+ N_A_1549_74#_c_1106_n N_A_1549_74#_c_1107_n N_A_1549_74#_c_1108_n
+ N_A_1549_74#_c_1109_n N_A_1549_74#_c_1110_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_1%A_1549_74#
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%A_1348_368# N_A_1348_368#_M1015_d
+ N_A_1348_368#_M1034_d N_A_1348_368#_M1004_g N_A_1348_368#_c_1319_n
+ N_A_1348_368#_c_1333_n N_A_1348_368#_M1008_g N_A_1348_368#_c_1320_n
+ N_A_1348_368#_M1042_g N_A_1348_368#_c_1335_n N_A_1348_368#_c_1336_n
+ N_A_1348_368#_M1025_g N_A_1348_368#_c_1322_n N_A_1348_368#_M1030_g
+ N_A_1348_368#_M1031_g N_A_1348_368#_c_1324_n N_A_1348_368#_c_1325_n
+ N_A_1348_368#_c_1326_n N_A_1348_368#_c_1327_n N_A_1348_368#_c_1328_n
+ N_A_1348_368#_c_1329_n N_A_1348_368#_c_1330_n N_A_1348_368#_c_1341_n
+ N_A_1348_368#_c_1342_n N_A_1348_368#_c_1343_n N_A_1348_368#_c_1344_n
+ N_A_1348_368#_c_1345_n N_A_1348_368#_c_1346_n N_A_1348_368#_c_1347_n
+ N_A_1348_368#_c_1348_n N_A_1348_368#_c_1331_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_1%A_1348_368#
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%A_1972_92# N_A_1972_92#_M1035_d
+ N_A_1972_92#_M1005_d N_A_1972_92#_M1022_g N_A_1972_92#_c_1517_n
+ N_A_1972_92#_c_1530_n N_A_1972_92#_M1041_g N_A_1972_92#_c_1518_n
+ N_A_1972_92#_c_1519_n N_A_1972_92#_c_1532_n N_A_1972_92#_M1038_g
+ N_A_1972_92#_c_1520_n N_A_1972_92#_M1016_g N_A_1972_92#_c_1521_n
+ N_A_1972_92#_c_1533_n N_A_1972_92#_c_1522_n N_A_1972_92#_c_1523_n
+ N_A_1972_92#_c_1524_n N_A_1972_92#_c_1525_n N_A_1972_92#_c_1526_n
+ N_A_1972_92#_c_1527_n N_A_1972_92#_c_1528_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_1%A_1972_92#
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%A_1747_118# N_A_1747_118#_M1042_d
+ N_A_1747_118#_M1017_d N_A_1747_118#_c_1623_n N_A_1747_118#_M1005_g
+ N_A_1747_118#_M1035_g N_A_1747_118#_c_1625_n N_A_1747_118#_c_1630_n
+ N_A_1747_118#_c_1650_n N_A_1747_118#_c_1626_n N_A_1747_118#_c_1631_n
+ N_A_1747_118#_c_1632_n N_A_1747_118#_c_1627_n N_A_1747_118#_c_1628_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_1%A_1747_118#
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%A_2463_74# N_A_2463_74#_M1018_d
+ N_A_2463_74#_M1030_d N_A_2463_74#_M1028_g N_A_2463_74#_c_1715_n
+ N_A_2463_74#_c_1727_n N_A_2463_74#_M1002_g N_A_2463_74#_c_1716_n
+ N_A_2463_74#_c_1717_n N_A_2463_74#_c_1718_n N_A_2463_74#_M1036_g
+ N_A_2463_74#_c_1719_n N_A_2463_74#_c_1720_n N_A_2463_74#_c_1729_n
+ N_A_2463_74#_M1027_g N_A_2463_74#_c_1800_n N_A_2463_74#_c_1721_n
+ N_A_2463_74#_c_1722_n N_A_2463_74#_c_1730_n N_A_2463_74#_c_1731_n
+ N_A_2463_74#_c_1732_n N_A_2463_74#_c_1723_n N_A_2463_74#_c_1724_n
+ N_A_2463_74#_c_1734_n N_A_2463_74#_c_1725_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_1%A_2463_74#
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%A_27_90# N_A_27_90#_M1013_s N_A_27_90#_M1001_d
+ N_A_27_90#_M1023_s N_A_27_90#_M1011_d N_A_27_90#_c_1869_n N_A_27_90#_c_1875_n
+ N_A_27_90#_c_1876_n N_A_27_90#_c_1877_n N_A_27_90#_c_1878_n
+ N_A_27_90#_c_1879_n N_A_27_90#_c_1908_n N_A_27_90#_c_1880_n
+ N_A_27_90#_c_1881_n N_A_27_90#_c_1870_n N_A_27_90#_c_1871_n
+ N_A_27_90#_c_1872_n N_A_27_90#_c_1883_n N_A_27_90#_c_1873_n
+ N_A_27_90#_c_1884_n PM_SKY130_FD_SC_LS__SEDFXBP_1%A_27_90#
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%VPWR N_VPWR_M1029_d N_VPWR_M1019_d
+ N_VPWR_M1003_d N_VPWR_M1034_s N_VPWR_M1008_s N_VPWR_M1041_d N_VPWR_M1038_s
+ N_VPWR_M1039_d N_VPWR_M1027_d N_VPWR_c_1992_n N_VPWR_c_1993_n N_VPWR_c_1994_n
+ N_VPWR_c_1995_n N_VPWR_c_1996_n N_VPWR_c_1997_n N_VPWR_c_1998_n
+ N_VPWR_c_1999_n N_VPWR_c_2000_n VPWR N_VPWR_c_2001_n N_VPWR_c_2002_n
+ N_VPWR_c_2003_n N_VPWR_c_2004_n N_VPWR_c_2005_n N_VPWR_c_2006_n
+ N_VPWR_c_2007_n N_VPWR_c_2008_n N_VPWR_c_2009_n N_VPWR_c_2010_n
+ N_VPWR_c_1991_n N_VPWR_c_2012_n N_VPWR_c_2013_n N_VPWR_c_2014_n
+ N_VPWR_c_2015_n N_VPWR_c_2016_n N_VPWR_c_2017_n N_VPWR_c_2018_n
+ N_VPWR_c_2019_n N_VPWR_c_2020_n PM_SKY130_FD_SC_LS__SEDFXBP_1%VPWR
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%A_697_113# N_A_697_113#_M1026_d
+ N_A_697_113#_M1010_d N_A_697_113#_M1042_s N_A_697_113#_M1021_d
+ N_A_697_113#_M1007_d N_A_697_113#_M1017_s N_A_697_113#_c_2180_n
+ N_A_697_113#_c_2181_n N_A_697_113#_c_2182_n N_A_697_113#_c_2183_n
+ N_A_697_113#_c_2208_n N_A_697_113#_c_2184_n N_A_697_113#_c_2173_n
+ N_A_697_113#_c_2186_n N_A_697_113#_c_2187_n N_A_697_113#_c_2174_n
+ N_A_697_113#_c_2175_n N_A_697_113#_c_2200_n N_A_697_113#_c_2265_n
+ N_A_697_113#_c_2176_n N_A_697_113#_c_2188_n N_A_697_113#_c_2189_n
+ N_A_697_113#_c_2177_n N_A_697_113#_c_2178_n N_A_697_113#_c_2191_n
+ N_A_697_113#_c_2192_n N_A_697_113#_c_2193_n N_A_697_113#_c_2179_n
+ N_A_697_113#_c_2333_n PM_SKY130_FD_SC_LS__SEDFXBP_1%A_697_113#
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%Q N_Q_M1036_s N_Q_M1027_s N_Q_c_2349_n Q Q Q Q
+ PM_SKY130_FD_SC_LS__SEDFXBP_1%Q
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%Q_N N_Q_N_M1000_d N_Q_N_M1040_d N_Q_N_c_2375_n
+ N_Q_N_c_2376_n Q_N Q_N Q_N Q_N N_Q_N_c_2377_n
+ PM_SKY130_FD_SC_LS__SEDFXBP_1%Q_N
x_PM_SKY130_FD_SC_LS__SEDFXBP_1%VGND N_VGND_M1014_d N_VGND_M1012_d
+ N_VGND_M1037_d N_VGND_M1015_s N_VGND_M1004_s N_VGND_M1022_d N_VGND_M1016_s
+ N_VGND_M1032_d N_VGND_M1036_d N_VGND_c_2397_n N_VGND_c_2398_n N_VGND_c_2399_n
+ N_VGND_c_2400_n N_VGND_c_2401_n N_VGND_c_2402_n N_VGND_c_2403_n
+ N_VGND_c_2404_n N_VGND_c_2405_n N_VGND_c_2406_n N_VGND_c_2407_n
+ N_VGND_c_2408_n VGND N_VGND_c_2409_n N_VGND_c_2410_n N_VGND_c_2411_n
+ N_VGND_c_2412_n N_VGND_c_2413_n N_VGND_c_2414_n N_VGND_c_2415_n
+ N_VGND_c_2416_n N_VGND_c_2417_n N_VGND_c_2418_n N_VGND_c_2419_n
+ N_VGND_c_2420_n N_VGND_c_2421_n N_VGND_c_2422_n N_VGND_c_2423_n
+ N_VGND_c_2424_n PM_SKY130_FD_SC_LS__SEDFXBP_1%VGND
cc_1 VNB N_D_c_337_n 0.0257586f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.545
cc_2 VNB N_D_M1013_g 0.0256701f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.66
cc_3 VNB N_D_c_339_n 0.00860311f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.73
cc_4 VNB N_D_c_340_n 0.0206728f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.225
cc_5 VNB N_D_c_341_n 0.00878149f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.225
cc_6 VNB N_A_161_394#_M1009_g 0.0423657f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.73
cc_7 VNB N_A_161_394#_c_380_n 0.00324511f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.06
cc_8 VNB N_A_161_394#_c_381_n 0.0197974f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.225
cc_9 VNB N_A_161_394#_c_382_n 0.00679172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_161_394#_c_383_n 0.00111842f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.295
cc_11 VNB N_A_161_394#_c_384_n 0.00912528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_161_394#_c_385_n 0.00271375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_161_394#_c_386_n 0.0145505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_DE_M1014_g 0.0239075f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.73
cc_15 VNB N_DE_c_492_n 0.0395716f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_16 VNB N_DE_c_493_n 0.00619153f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_17 VNB N_DE_c_494_n 0.0178603f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_18 VNB N_DE_c_495_n 0.0214729f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.295
cc_19 VNB N_DE_c_496_n 0.0168283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_DE_c_497_n 0.00465944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_DE_c_498_n 0.0167209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_575_305#_M1001_g 0.0404596f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.66
cc_23 VNB N_A_575_305#_c_578_n 0.0170882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_575_305#_c_579_n 0.0388921f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.225
cc_25 VNB N_A_575_305#_c_580_n 0.00716124f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.06
cc_26 VNB N_A_575_305#_c_581_n 0.0339623f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.665
cc_27 VNB N_A_575_305#_c_582_n 0.0335406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_575_305#_M1000_g 0.028168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_575_305#_c_584_n 0.00491486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_575_305#_c_585_n 0.0084524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_575_305#_c_586_n 0.0143213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_575_305#_c_587_n 0.00367455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_575_305#_c_588_n 7.76083e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_575_305#_c_589_n 0.00299714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_575_305#_c_590_n 0.00913009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_575_305#_c_591_n 0.00436426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_575_305#_c_592_n 0.0156253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_575_305#_c_593_n 0.00259103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_667_87#_c_836_n 0.0161363f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_40 VNB N_A_667_87#_c_837_n 0.0369865f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.66
cc_41 VNB N_A_667_87#_c_838_n 0.00865069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_667_87#_c_839_n 0.00887253f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.225
cc_43 VNB N_A_667_87#_c_840_n 0.0354104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_667_87#_c_841_n 0.0614006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_667_87#_c_842_n 0.0158654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_SCD_c_927_n 0.0106811f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.545
cc_47 VNB N_SCD_M1024_g 0.0164747f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.06
cc_48 VNB SCD 0.0189074f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.66
cc_49 VNB N_SCD_c_930_n 0.0339713f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_50 VNB N_SCE_M1037_g 0.0487723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_SCE_c_973_n 0.0654138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_SCE_c_974_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.225
cc_53 VNB N_SCE_M1010_g 0.0375422f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.06
cc_54 VNB N_SCE_c_976_n 0.0177212f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.665
cc_55 VNB N_SCE_c_977_n 0.0042092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_CLK_c_1052_n 0.0458321f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.245
cc_57 VNB N_CLK_c_1053_n 0.0216597f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.155
cc_58 VNB CLK 0.0136832f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_59 VNB N_A_1549_74#_M1018_g 0.0355212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1549_74#_c_1088_n 0.00575788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1549_74#_c_1089_n 0.00955967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1549_74#_c_1090_n 0.0208222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1549_74#_c_1091_n 0.00361019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1549_74#_c_1092_n 0.023079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1549_74#_c_1093_n 0.00421456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1549_74#_c_1094_n 0.00772673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1549_74#_c_1095_n 0.00921403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1549_74#_c_1096_n 0.00195347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1549_74#_c_1097_n 0.00956756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1549_74#_c_1098_n 0.00506047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1549_74#_c_1099_n 0.00321401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1549_74#_c_1100_n 0.00319118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1549_74#_c_1101_n 0.00111521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1549_74#_c_1102_n 0.018076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1549_74#_c_1103_n 0.00733234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1549_74#_c_1104_n 0.00139474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1549_74#_c_1105_n 0.00653741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1549_74#_c_1106_n 0.0345165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1549_74#_c_1107_n 0.00292381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1549_74#_c_1108_n 0.0300273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1549_74#_c_1109_n 0.0195571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1549_74#_c_1110_n 0.0196812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1348_368#_M1004_g 0.048522f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.66
cc_84 VNB N_A_1348_368#_c_1319_n 0.00519935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1348_368#_c_1320_n 0.0125595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1348_368#_M1042_g 0.0493193f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.06
cc_87 VNB N_A_1348_368#_c_1322_n 0.015283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1348_368#_M1031_g 0.05116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1348_368#_c_1324_n 0.0179649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1348_368#_c_1325_n 0.00499721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1348_368#_c_1326_n 0.00200062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1348_368#_c_1327_n 0.00806055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1348_368#_c_1328_n 0.0115444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1348_368#_c_1329_n 3.04083e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1348_368#_c_1330_n 0.0112028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1348_368#_c_1331_n 0.00385141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1972_92#_M1022_g 0.0228279f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.66
cc_98 VNB N_A_1972_92#_c_1517_n 0.0142601f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.73
cc_99 VNB N_A_1972_92#_c_1518_n 0.0341591f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.225
cc_100 VNB N_A_1972_92#_c_1519_n 0.00889414f $X=-0.19 $Y=-0.245 $X2=0.62
+ $Y2=1.225
cc_101 VNB N_A_1972_92#_c_1520_n 0.0198235f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.295
cc_102 VNB N_A_1972_92#_c_1521_n 0.0125353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1972_92#_c_1522_n 0.00549523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1972_92#_c_1523_n 0.00260597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1972_92#_c_1524_n 0.00191104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1972_92#_c_1525_n 0.0590469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1972_92#_c_1526_n 0.031165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1972_92#_c_1527_n 0.00283223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1972_92#_c_1528_n 0.00172958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_1747_118#_c_1623_n 0.0204185f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.64
cc_111 VNB N_A_1747_118#_M1035_g 0.0427559f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.73
cc_112 VNB N_A_1747_118#_c_1625_n 0.0146697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1747_118#_c_1626_n 2.63561e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1747_118#_c_1627_n 0.00102942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_1747_118#_c_1628_n 0.0100709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_2463_74#_M1028_g 0.0251625f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.66
cc_117 VNB N_A_2463_74#_c_1715_n 0.0084305f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.73
cc_118 VNB N_A_2463_74#_c_1716_n 0.0576991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_2463_74#_c_1717_n 0.0377417f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.225
cc_120 VNB N_A_2463_74#_c_1718_n 0.0168831f $X=-0.19 $Y=-0.245 $X2=0.62
+ $Y2=1.225
cc_121 VNB N_A_2463_74#_c_1719_n 0.0155027f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.225
cc_122 VNB N_A_2463_74#_c_1720_n 0.0176486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_2463_74#_c_1721_n 0.00286498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_2463_74#_c_1722_n 0.0026364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_2463_74#_c_1723_n 0.00208726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_2463_74#_c_1724_n 0.00164929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_2463_74#_c_1725_n 0.00329462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_27_90#_c_1869_n 0.03964f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_129 VNB N_A_27_90#_c_1870_n 0.00395727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_27_90#_c_1871_n 0.00687596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_27_90#_c_1872_n 0.0135101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_27_90#_c_1873_n 0.00780487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VPWR_c_1991_n 0.681144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_697_113#_c_2173_n 0.0180421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_697_113#_c_2174_n 0.00995796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_697_113#_c_2175_n 0.00376624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_697_113#_c_2176_n 0.0161278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_A_697_113#_c_2177_n 0.0104448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_A_697_113#_c_2178_n 0.00835877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_697_113#_c_2179_n 0.0112976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_Q_c_2349_n 0.00610717f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.66
cc_142 VNB N_Q_N_c_2375_n 0.0266902f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.66
cc_143 VNB N_Q_N_c_2376_n 0.00950103f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_144 VNB N_Q_N_c_2377_n 0.0239414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2397_n 0.0229784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2398_n 0.0301741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2399_n 0.00778394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2400_n 0.00867342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2401_n 0.0098347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2402_n 0.0124808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2403_n 0.00590394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2404_n 0.0103909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2405_n 0.0214209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2406_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2407_n 0.0329502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2408_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2409_n 0.0354476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2410_n 0.0668922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2411_n 0.0209223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2412_n 0.0598226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2413_n 0.0296513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2414_n 0.0363431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2415_n 0.0193429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2416_n 0.89f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2417_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2418_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2419_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2420_n 0.0062513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2421_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2422_n 0.0403351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2423_n 0.0275281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2424_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VPB N_D_c_342_n 0.026035f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.155
cc_174 VPB N_D_c_343_n 0.0251075f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_175 VPB N_D_c_339_n 0.0106593f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.73
cc_176 VPB N_D_c_341_n 0.00420103f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.225
cc_177 VPB N_A_161_394#_c_387_n 0.0181954f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_178 VPB N_A_161_394#_c_388_n 0.0468826f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_179 VPB N_A_161_394#_c_381_n 0.026082f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.225
cc_180 VPB N_A_161_394#_c_390_n 0.0131197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_161_394#_c_391_n 0.00336961f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.665
cc_182 VPB N_A_161_394#_c_392_n 0.00823568f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_161_394#_c_393_n 0.011445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_161_394#_c_385_n 0.00169193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_161_394#_c_386_n 0.0174379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_161_394#_c_396_n 0.00141199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_DE_c_499_n 0.0205675f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=0.66
cc_188 VPB N_DE_c_500_n 0.0184461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_DE_c_501_n 0.0391066f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.225
cc_190 VPB N_DE_c_502_n 0.0165101f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.225
cc_191 VPB N_DE_c_503_n 0.00724793f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.665
cc_192 VPB N_DE_c_496_n 0.0123746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_DE_c_497_n 0.00346054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_575_305#_c_594_n 0.0224025f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.73
cc_195 VPB N_A_575_305#_c_595_n 0.0217529f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_196 VPB N_A_575_305#_c_596_n 0.0551894f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.225
cc_197 VPB N_A_575_305#_c_581_n 0.0211417f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.665
cc_198 VPB N_A_575_305#_c_582_n 0.0289703f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_575_305#_c_585_n 0.00585284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_575_305#_c_600_n 0.00185536f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_575_305#_c_601_n 0.0662214f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_575_305#_c_602_n 0.00214501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_575_305#_c_603_n 0.0024988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_575_305#_c_592_n 0.0195159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_575_305#_c_593_n 0.00388881f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_575_305#_c_606_n 0.00489778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_575_305#_c_607_n 0.00461807f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_667_87#_c_843_n 0.0623088f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.73
cc_209 VPB N_A_667_87#_c_840_n 0.0436189f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_667_87#_c_845_n 0.0038203f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_667_87#_c_846_n 0.0288765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_667_87#_c_847_n 0.00341614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_667_87#_c_848_n 0.00621254f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_667_87#_c_849_n 0.00775817f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_SCD_c_927_n 0.0285682f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.545
cc_216 VPB N_SCD_c_932_n 0.0210132f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.73
cc_217 VPB N_SCE_c_978_n 0.0160619f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.245
cc_218 VPB N_SCE_c_979_n 0.0872209f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.155
cc_219 VPB N_SCE_c_980_n 0.0128697f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_220 VPB N_SCE_c_981_n 0.0206854f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_221 VPB N_SCE_c_982_n 0.00702891f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.06
cc_222 VPB N_SCE_M1003_g 0.00927731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_SCE_c_976_n 0.0110457f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.665
cc_224 VPB N_SCE_c_977_n 0.00259215f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_CLK_c_1052_n 0.0300141f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.245
cc_226 VPB N_A_1549_74#_c_1111_n 0.0202965f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_227 VPB N_A_1549_74#_c_1112_n 0.00498378f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.225
cc_228 VPB N_A_1549_74#_c_1113_n 0.0126529f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.225
cc_229 VPB N_A_1549_74#_c_1114_n 0.0219728f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.225
cc_230 VPB N_A_1549_74#_c_1088_n 0.0190642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_1549_74#_c_1116_n 0.0108227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_1549_74#_c_1101_n 0.00362877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_1549_74#_c_1103_n 2.75058e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_1549_74#_c_1119_n 0.0560771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_1549_74#_c_1110_n 0.0208843f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_1348_368#_c_1319_n 0.00684676f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_1348_368#_c_1333_n 0.0207807f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_238 VPB N_A_1348_368#_c_1320_n 0.0150145f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_1348_368#_c_1335_n 0.0440712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_1348_368#_c_1336_n 0.0723303f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_1348_368#_c_1322_n 0.0417731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_1348_368#_c_1324_n 0.0132907f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_1348_368#_c_1325_n 0.00167153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_1348_368#_c_1326_n 0.00693389f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_1348_368#_c_1341_n 0.0056838f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_1348_368#_c_1342_n 0.00264345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_1348_368#_c_1343_n 0.0107744f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_1348_368#_c_1344_n 0.00103733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_1348_368#_c_1345_n 0.00413334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_1348_368#_c_1346_n 0.0362079f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_1348_368#_c_1347_n 0.00311017f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_A_1348_368#_c_1348_n 0.00829487f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_A_1348_368#_c_1331_n 0.00222147f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_A_1972_92#_c_1517_n 0.040329f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.73
cc_255 VPB N_A_1972_92#_c_1530_n 0.0219277f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_256 VPB N_A_1972_92#_c_1519_n 0.00857421f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.225
cc_257 VPB N_A_1972_92#_c_1532_n 0.0308626f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.06
cc_258 VPB N_A_1972_92#_c_1533_n 0.00461792f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_A_1972_92#_c_1523_n 0.00968251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_A_1747_118#_c_1623_n 0.0453428f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_261 VPB N_A_1747_118#_c_1630_n 0.00288391f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.06
cc_262 VPB N_A_1747_118#_c_1631_n 0.00639558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_A_1747_118#_c_1632_n 0.00199044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_1747_118#_c_1627_n 4.51094e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_A_1747_118#_c_1628_n 0.00634007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_A_2463_74#_c_1715_n 0.00875712f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.73
cc_267 VPB N_A_2463_74#_c_1727_n 0.0265917f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_268 VPB N_A_2463_74#_c_1720_n 8.80765e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_A_2463_74#_c_1729_n 0.0268658f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.295
cc_270 VPB N_A_2463_74#_c_1730_n 0.00565678f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_2463_74#_c_1731_n 0.0134523f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_A_2463_74#_c_1732_n 0.00205362f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_A_2463_74#_c_1724_n 5.43958e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_2463_74#_c_1734_n 0.00367038f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_A_27_90#_c_1869_n 0.0306822f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_276 VPB N_A_27_90#_c_1875_n 0.0224775f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.225
cc_277 VPB N_A_27_90#_c_1876_n 0.0136f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.225
cc_278 VPB N_A_27_90#_c_1877_n 0.00998336f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_27_90#_c_1878_n 0.00949465f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.295
cc_280 VPB N_A_27_90#_c_1879_n 0.00349119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_27_90#_c_1880_n 0.00660395f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_A_27_90#_c_1881_n 0.00109302f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_27_90#_c_1871_n 0.0094187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_A_27_90#_c_1883_n 0.0126424f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_27_90#_c_1884_n 0.00468081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_VPWR_c_1992_n 0.00600898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_VPWR_c_1993_n 0.00543965f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_288 VPB N_VPWR_c_1994_n 0.00573048f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_289 VPB N_VPWR_c_1995_n 0.0102206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_VPWR_c_1996_n 0.0220341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_1997_n 0.0115779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_VPWR_c_1998_n 0.0162479f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_VPWR_c_1999_n 0.00608393f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_VPWR_c_2000_n 0.0112275f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_VPWR_c_2001_n 0.029813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_2002_n 0.0296515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_VPWR_c_2003_n 0.0599825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_VPWR_c_2004_n 0.0313657f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_2005_n 0.0335097f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_300 VPB N_VPWR_c_2006_n 0.0567382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_301 VPB N_VPWR_c_2007_n 0.0242802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_302 VPB N_VPWR_c_2008_n 0.0643658f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_303 VPB N_VPWR_c_2009_n 0.0339005f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_2010_n 0.0192773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_305 VPB N_VPWR_c_1991_n 0.194333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_2012_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_2013_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_2014_n 0.00467461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_309 VPB N_VPWR_c_2015_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_310 VPB N_VPWR_c_2016_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_2017_n 0.00615076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_312 VPB N_VPWR_c_2018_n 0.00632182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_313 VPB N_VPWR_c_2019_n 0.010962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_314 VPB N_VPWR_c_2020_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_315 VPB N_A_697_113#_c_2180_n 0.00236938f $X=-0.19 $Y=1.66 $X2=0.645
+ $Y2=1.225
cc_316 VPB N_A_697_113#_c_2181_n 0.00457103f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_317 VPB N_A_697_113#_c_2182_n 0.0077302f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.665
cc_318 VPB N_A_697_113#_c_2183_n 7.12198e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_319 VPB N_A_697_113#_c_2184_n 3.43064e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_320 VPB N_A_697_113#_c_2173_n 0.0160595f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_321 VPB N_A_697_113#_c_2186_n 0.0219398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_322 VPB N_A_697_113#_c_2187_n 0.00112537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_323 VPB N_A_697_113#_c_2188_n 0.00168863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_324 VPB N_A_697_113#_c_2189_n 0.011749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_325 VPB N_A_697_113#_c_2178_n 0.0114561f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_326 VPB N_A_697_113#_c_2191_n 0.00824945f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_327 VPB N_A_697_113#_c_2192_n 0.0046419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_328 VPB N_A_697_113#_c_2193_n 0.00735455f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_329 VPB N_Q_c_2349_n 0.00381055f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=0.66
cc_330 VPB Q 0.00674277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_331 VPB Q 0.0140623f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.06
cc_332 VPB Q_N 0.0100754f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_333 VPB Q_N 0.042262f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.295
cc_334 VPB N_Q_N_c_2377_n 0.00776947f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_335 N_D_c_343_n N_A_161_394#_c_387_n 0.0437552f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_336 N_D_c_342_n N_A_161_394#_c_388_n 0.018058f $X=0.505 $Y=2.155 $X2=0 $Y2=0
cc_337 N_D_c_341_n N_A_161_394#_c_388_n 8.40458e-19 $X=0.62 $Y=1.225 $X2=0 $Y2=0
cc_338 N_D_c_337_n N_A_161_394#_c_380_n 0.00140836f $X=0.6 $Y=1.545 $X2=0 $Y2=0
cc_339 N_D_c_342_n N_A_161_394#_c_380_n 0.00102045f $X=0.505 $Y=2.155 $X2=0
+ $Y2=0
cc_340 N_D_c_341_n N_A_161_394#_c_380_n 0.0374911f $X=0.62 $Y=1.225 $X2=0 $Y2=0
cc_341 N_D_c_337_n N_A_161_394#_c_381_n 0.0147863f $X=0.6 $Y=1.545 $X2=0 $Y2=0
cc_342 N_D_c_342_n N_A_161_394#_c_381_n 0.00688788f $X=0.505 $Y=2.155 $X2=0
+ $Y2=0
cc_343 N_D_c_341_n N_A_161_394#_c_381_n 0.00214371f $X=0.62 $Y=1.225 $X2=0 $Y2=0
cc_344 N_D_c_340_n N_A_161_394#_c_383_n 5.92811e-19 $X=0.62 $Y=1.225 $X2=0 $Y2=0
cc_345 N_D_c_341_n N_A_161_394#_c_383_n 0.0135781f $X=0.62 $Y=1.225 $X2=0 $Y2=0
cc_346 N_D_c_342_n N_A_161_394#_c_391_n 7.41315e-19 $X=0.505 $Y=2.155 $X2=0
+ $Y2=0
cc_347 N_D_M1013_g N_DE_M1014_g 0.0235118f $X=0.71 $Y=0.66 $X2=0 $Y2=0
cc_348 N_D_c_340_n N_DE_c_493_n 0.0235118f $X=0.62 $Y=1.225 $X2=0 $Y2=0
cc_349 N_D_c_341_n N_DE_c_493_n 0.001576f $X=0.62 $Y=1.225 $X2=0 $Y2=0
cc_350 N_D_c_343_n N_A_27_90#_c_1869_n 0.00154775f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_351 N_D_M1013_g N_A_27_90#_c_1869_n 0.0066353f $X=0.71 $Y=0.66 $X2=0 $Y2=0
cc_352 N_D_c_340_n N_A_27_90#_c_1869_n 0.0340525f $X=0.62 $Y=1.225 $X2=0 $Y2=0
cc_353 N_D_c_341_n N_A_27_90#_c_1869_n 0.0545845f $X=0.62 $Y=1.225 $X2=0 $Y2=0
cc_354 N_D_c_343_n N_A_27_90#_c_1875_n 0.00907263f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_355 N_D_c_343_n N_A_27_90#_c_1876_n 0.0136133f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_356 N_D_c_339_n N_A_27_90#_c_1876_n 9.37516e-19 $X=0.6 $Y=1.73 $X2=0 $Y2=0
cc_357 N_D_c_341_n N_A_27_90#_c_1876_n 0.0137727f $X=0.62 $Y=1.225 $X2=0 $Y2=0
cc_358 N_D_M1013_g N_A_27_90#_c_1872_n 0.00620944f $X=0.71 $Y=0.66 $X2=0 $Y2=0
cc_359 N_D_c_340_n N_A_27_90#_c_1872_n 0.00272163f $X=0.62 $Y=1.225 $X2=0 $Y2=0
cc_360 N_D_c_341_n N_A_27_90#_c_1872_n 0.0107166f $X=0.62 $Y=1.225 $X2=0 $Y2=0
cc_361 N_D_c_343_n N_A_27_90#_c_1883_n 0.00237313f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_362 N_D_c_343_n N_VPWR_c_1992_n 0.0015335f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_363 N_D_c_343_n N_VPWR_c_2001_n 0.00445602f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_364 N_D_c_343_n N_VPWR_c_1991_n 0.00861358f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_365 N_D_M1013_g N_VGND_c_2397_n 0.00212753f $X=0.71 $Y=0.66 $X2=0 $Y2=0
cc_366 N_D_M1013_g N_VGND_c_2409_n 0.00497885f $X=0.71 $Y=0.66 $X2=0 $Y2=0
cc_367 N_D_M1013_g N_VGND_c_2416_n 0.00520574f $X=0.71 $Y=0.66 $X2=0 $Y2=0
cc_368 N_A_161_394#_c_384_n N_DE_M1014_g 0.00497053f $X=1.875 $Y=0.775 $X2=0
+ $Y2=0
cc_369 N_A_161_394#_c_382_n N_DE_c_492_n 0.0193426f $X=1.71 $Y=1.195 $X2=0 $Y2=0
cc_370 N_A_161_394#_c_383_n N_DE_c_492_n 0.00569077f $X=1.355 $Y=1.195 $X2=0
+ $Y2=0
cc_371 N_A_161_394#_c_384_n N_DE_c_492_n 0.0035123f $X=1.875 $Y=0.775 $X2=0
+ $Y2=0
cc_372 N_A_161_394#_c_381_n N_DE_c_493_n 0.0182409f $X=1.19 $Y=1.615 $X2=0 $Y2=0
cc_373 N_A_161_394#_c_383_n N_DE_c_493_n 0.00994624f $X=1.355 $Y=1.195 $X2=0
+ $Y2=0
cc_374 N_A_161_394#_c_380_n N_DE_c_499_n 8.54735e-19 $X=1.19 $Y=1.615 $X2=0
+ $Y2=0
cc_375 N_A_161_394#_c_381_n N_DE_c_499_n 0.0031603f $X=1.19 $Y=1.615 $X2=0 $Y2=0
cc_376 N_A_161_394#_c_393_n N_DE_c_499_n 0.0100993f $X=2.335 $Y=2.035 $X2=0
+ $Y2=0
cc_377 N_A_161_394#_c_385_n N_DE_c_499_n 0.00321563f $X=2.5 $Y=1.69 $X2=0 $Y2=0
cc_378 N_A_161_394#_c_392_n N_DE_c_500_n 0.00429303f $X=1.8 $Y=2.515 $X2=0 $Y2=0
cc_379 N_A_161_394#_M1009_g N_DE_c_494_n 0.0184318f $X=2.59 $Y=0.775 $X2=0 $Y2=0
cc_380 N_A_161_394#_c_384_n N_DE_c_494_n 0.00860606f $X=1.875 $Y=0.775 $X2=0
+ $Y2=0
cc_381 N_A_161_394#_c_393_n N_DE_c_501_n 0.0152013f $X=2.335 $Y=2.035 $X2=0
+ $Y2=0
cc_382 N_A_161_394#_c_386_n N_DE_c_501_n 0.0181536f $X=2.5 $Y=1.69 $X2=0 $Y2=0
cc_383 N_A_161_394#_c_382_n N_DE_c_495_n 0.00511954f $X=1.71 $Y=1.195 $X2=0
+ $Y2=0
cc_384 N_A_161_394#_c_384_n N_DE_c_495_n 0.0060005f $X=1.875 $Y=0.775 $X2=0
+ $Y2=0
cc_385 N_A_161_394#_c_388_n N_DE_c_503_n 0.0031603f $X=0.895 $Y=2.107 $X2=0
+ $Y2=0
cc_386 N_A_161_394#_c_392_n N_DE_c_503_n 0.00589429f $X=1.8 $Y=2.515 $X2=0 $Y2=0
cc_387 N_A_161_394#_c_393_n N_DE_c_503_n 0.00696573f $X=2.335 $Y=2.035 $X2=0
+ $Y2=0
cc_388 N_A_161_394#_M1009_g N_DE_c_496_n 0.00178228f $X=2.59 $Y=0.775 $X2=0
+ $Y2=0
cc_389 N_A_161_394#_c_380_n N_DE_c_496_n 3.17712e-19 $X=1.19 $Y=1.615 $X2=0
+ $Y2=0
cc_390 N_A_161_394#_c_381_n N_DE_c_496_n 0.00868804f $X=1.19 $Y=1.615 $X2=0
+ $Y2=0
cc_391 N_A_161_394#_c_382_n N_DE_c_496_n 9.53276e-19 $X=1.71 $Y=1.195 $X2=0
+ $Y2=0
cc_392 N_A_161_394#_c_393_n N_DE_c_496_n 0.00119763f $X=2.335 $Y=2.035 $X2=0
+ $Y2=0
cc_393 N_A_161_394#_c_385_n N_DE_c_496_n 8.11706e-19 $X=2.5 $Y=1.69 $X2=0 $Y2=0
cc_394 N_A_161_394#_c_386_n N_DE_c_496_n 0.0169432f $X=2.5 $Y=1.69 $X2=0 $Y2=0
cc_395 N_A_161_394#_c_396_n N_DE_c_496_n 0.00354118f $X=1.8 $Y=2.035 $X2=0 $Y2=0
cc_396 N_A_161_394#_M1009_g N_DE_c_497_n 4.1165e-19 $X=2.59 $Y=0.775 $X2=0 $Y2=0
cc_397 N_A_161_394#_c_380_n N_DE_c_497_n 0.0230897f $X=1.19 $Y=1.615 $X2=0 $Y2=0
cc_398 N_A_161_394#_c_381_n N_DE_c_497_n 0.00270561f $X=1.19 $Y=1.615 $X2=0
+ $Y2=0
cc_399 N_A_161_394#_c_382_n N_DE_c_497_n 0.0387962f $X=1.71 $Y=1.195 $X2=0 $Y2=0
cc_400 N_A_161_394#_c_390_n N_DE_c_497_n 0.0118552f $X=1.715 $Y=2.035 $X2=0
+ $Y2=0
cc_401 N_A_161_394#_c_393_n N_DE_c_497_n 0.0144321f $X=2.335 $Y=2.035 $X2=0
+ $Y2=0
cc_402 N_A_161_394#_c_385_n N_DE_c_497_n 0.0145619f $X=2.5 $Y=1.69 $X2=0 $Y2=0
cc_403 N_A_161_394#_c_386_n N_DE_c_497_n 9.49267e-19 $X=2.5 $Y=1.69 $X2=0 $Y2=0
cc_404 N_A_161_394#_c_396_n N_DE_c_497_n 0.0145018f $X=1.8 $Y=2.035 $X2=0 $Y2=0
cc_405 N_A_161_394#_M1009_g N_DE_c_498_n 0.00513217f $X=2.59 $Y=0.775 $X2=0
+ $Y2=0
cc_406 N_A_161_394#_c_380_n N_DE_c_498_n 0.0049143f $X=1.19 $Y=1.615 $X2=0 $Y2=0
cc_407 N_A_161_394#_c_382_n N_DE_c_498_n 0.00568535f $X=1.71 $Y=1.195 $X2=0
+ $Y2=0
cc_408 N_A_161_394#_M1009_g N_A_575_305#_M1001_g 0.0568001f $X=2.59 $Y=0.775
+ $X2=0 $Y2=0
cc_409 N_A_161_394#_c_393_n N_A_575_305#_c_594_n 8.17703e-19 $X=2.335 $Y=2.035
+ $X2=0 $Y2=0
cc_410 N_A_161_394#_c_385_n N_A_575_305#_c_594_n 4.77843e-19 $X=2.5 $Y=1.69
+ $X2=0 $Y2=0
cc_411 N_A_161_394#_c_393_n N_A_575_305#_c_602_n 0.00110012f $X=2.335 $Y=2.035
+ $X2=0 $Y2=0
cc_412 N_A_161_394#_c_385_n N_A_575_305#_c_592_n 0.00115578f $X=2.5 $Y=1.69
+ $X2=0 $Y2=0
cc_413 N_A_161_394#_c_386_n N_A_575_305#_c_592_n 0.0201559f $X=2.5 $Y=1.69 $X2=0
+ $Y2=0
cc_414 N_A_161_394#_c_393_n N_A_575_305#_c_593_n 0.0115373f $X=2.335 $Y=2.035
+ $X2=0 $Y2=0
cc_415 N_A_161_394#_c_385_n N_A_575_305#_c_593_n 0.0274959f $X=2.5 $Y=1.69 $X2=0
+ $Y2=0
cc_416 N_A_161_394#_c_386_n N_A_575_305#_c_593_n 0.00114936f $X=2.5 $Y=1.69
+ $X2=0 $Y2=0
cc_417 N_A_161_394#_c_387_n N_A_27_90#_c_1875_n 0.00180343f $X=0.895 $Y=2.245
+ $X2=0 $Y2=0
cc_418 N_A_161_394#_c_387_n N_A_27_90#_c_1876_n 0.0197185f $X=0.895 $Y=2.245
+ $X2=0 $Y2=0
cc_419 N_A_161_394#_c_388_n N_A_27_90#_c_1876_n 0.00474236f $X=0.895 $Y=2.107
+ $X2=0 $Y2=0
cc_420 N_A_161_394#_c_390_n N_A_27_90#_c_1876_n 0.015789f $X=1.715 $Y=2.035
+ $X2=0 $Y2=0
cc_421 N_A_161_394#_c_391_n N_A_27_90#_c_1876_n 0.0263722f $X=1.355 $Y=2.035
+ $X2=0 $Y2=0
cc_422 N_A_161_394#_c_392_n N_A_27_90#_c_1876_n 0.0141715f $X=1.8 $Y=2.515 $X2=0
+ $Y2=0
cc_423 N_A_161_394#_c_387_n N_A_27_90#_c_1877_n 0.00426176f $X=0.895 $Y=2.245
+ $X2=0 $Y2=0
cc_424 N_A_161_394#_c_392_n N_A_27_90#_c_1877_n 0.0203028f $X=1.8 $Y=2.515 $X2=0
+ $Y2=0
cc_425 N_A_161_394#_M1019_s N_A_27_90#_c_1878_n 0.00480049f $X=1.655 $Y=2.32
+ $X2=0 $Y2=0
cc_426 N_A_161_394#_c_392_n N_A_27_90#_c_1878_n 0.012787f $X=1.8 $Y=2.515 $X2=0
+ $Y2=0
cc_427 N_A_161_394#_c_387_n N_A_27_90#_c_1879_n 6.5162e-19 $X=0.895 $Y=2.245
+ $X2=0 $Y2=0
cc_428 N_A_161_394#_c_392_n N_A_27_90#_c_1908_n 0.0178681f $X=1.8 $Y=2.515 $X2=0
+ $Y2=0
cc_429 N_A_161_394#_c_393_n N_A_27_90#_c_1880_n 0.0309808f $X=2.335 $Y=2.035
+ $X2=0 $Y2=0
cc_430 N_A_161_394#_c_386_n N_A_27_90#_c_1880_n 2.47837e-19 $X=2.5 $Y=1.69 $X2=0
+ $Y2=0
cc_431 N_A_161_394#_c_392_n N_A_27_90#_c_1881_n 0.0133747f $X=1.8 $Y=2.515 $X2=0
+ $Y2=0
cc_432 N_A_161_394#_c_393_n N_A_27_90#_c_1881_n 0.0123833f $X=2.335 $Y=2.035
+ $X2=0 $Y2=0
cc_433 N_A_161_394#_M1009_g N_A_27_90#_c_1870_n 0.00214472f $X=2.59 $Y=0.775
+ $X2=0 $Y2=0
cc_434 N_A_161_394#_M1009_g N_A_27_90#_c_1873_n 8.28834e-19 $X=2.59 $Y=0.775
+ $X2=0 $Y2=0
cc_435 N_A_161_394#_c_387_n N_VPWR_c_1992_n 0.0104537f $X=0.895 $Y=2.245 $X2=0
+ $Y2=0
cc_436 N_A_161_394#_c_387_n N_VPWR_c_2001_n 0.00413917f $X=0.895 $Y=2.245 $X2=0
+ $Y2=0
cc_437 N_A_161_394#_c_387_n N_VPWR_c_1991_n 0.00817239f $X=0.895 $Y=2.245 $X2=0
+ $Y2=0
cc_438 N_A_161_394#_c_381_n N_VGND_c_2397_n 2.29105e-19 $X=1.19 $Y=1.615 $X2=0
+ $Y2=0
cc_439 N_A_161_394#_c_382_n N_VGND_c_2397_n 0.00822581f $X=1.71 $Y=1.195 $X2=0
+ $Y2=0
cc_440 N_A_161_394#_c_383_n N_VGND_c_2397_n 0.0148248f $X=1.355 $Y=1.195 $X2=0
+ $Y2=0
cc_441 N_A_161_394#_c_384_n N_VGND_c_2397_n 0.0232594f $X=1.875 $Y=0.775 $X2=0
+ $Y2=0
cc_442 N_A_161_394#_M1009_g N_VGND_c_2398_n 0.0129412f $X=2.59 $Y=0.775 $X2=0
+ $Y2=0
cc_443 N_A_161_394#_c_384_n N_VGND_c_2398_n 0.0188413f $X=1.875 $Y=0.775 $X2=0
+ $Y2=0
cc_444 N_A_161_394#_c_385_n N_VGND_c_2398_n 0.00760101f $X=2.5 $Y=1.69 $X2=0
+ $Y2=0
cc_445 N_A_161_394#_c_386_n N_VGND_c_2398_n 0.00118383f $X=2.5 $Y=1.69 $X2=0
+ $Y2=0
cc_446 N_A_161_394#_c_384_n N_VGND_c_2405_n 0.00805126f $X=1.875 $Y=0.775 $X2=0
+ $Y2=0
cc_447 N_A_161_394#_M1009_g N_VGND_c_2410_n 0.00372658f $X=2.59 $Y=0.775 $X2=0
+ $Y2=0
cc_448 N_A_161_394#_M1009_g N_VGND_c_2416_n 0.00408518f $X=2.59 $Y=0.775 $X2=0
+ $Y2=0
cc_449 N_A_161_394#_c_384_n N_VGND_c_2416_n 0.0106012f $X=1.875 $Y=0.775 $X2=0
+ $Y2=0
cc_450 N_DE_c_501_n N_A_575_305#_c_594_n 0.00907891f $X=2.63 $Y=2.17 $X2=0 $Y2=0
cc_451 N_DE_c_502_n N_A_575_305#_c_595_n 0.0384652f $X=2.705 $Y=2.245 $X2=0
+ $Y2=0
cc_452 N_DE_c_501_n N_A_575_305#_c_593_n 7.62429e-19 $X=2.63 $Y=2.17 $X2=0 $Y2=0
cc_453 N_DE_c_500_n N_A_27_90#_c_1877_n 0.00326422f $X=2.025 $Y=2.245 $X2=0
+ $Y2=0
cc_454 N_DE_c_500_n N_A_27_90#_c_1878_n 0.0135199f $X=2.025 $Y=2.245 $X2=0 $Y2=0
cc_455 N_DE_c_502_n N_A_27_90#_c_1878_n 4.24321e-19 $X=2.705 $Y=2.245 $X2=0
+ $Y2=0
cc_456 N_DE_c_500_n N_A_27_90#_c_1908_n 0.0113399f $X=2.025 $Y=2.245 $X2=0 $Y2=0
cc_457 N_DE_c_502_n N_A_27_90#_c_1908_n 0.00281561f $X=2.705 $Y=2.245 $X2=0
+ $Y2=0
cc_458 N_DE_c_501_n N_A_27_90#_c_1880_n 0.00748616f $X=2.63 $Y=2.17 $X2=0 $Y2=0
cc_459 N_DE_c_502_n N_A_27_90#_c_1880_n 0.0157312f $X=2.705 $Y=2.245 $X2=0 $Y2=0
cc_460 N_DE_c_500_n N_A_27_90#_c_1881_n 0.00592248f $X=2.025 $Y=2.245 $X2=0
+ $Y2=0
cc_461 N_DE_c_501_n N_A_27_90#_c_1881_n 8.10306e-19 $X=2.63 $Y=2.17 $X2=0 $Y2=0
cc_462 N_DE_M1014_g N_A_27_90#_c_1872_n 9.26497e-19 $X=1.1 $Y=0.66 $X2=0 $Y2=0
cc_463 N_DE_c_502_n N_A_27_90#_c_1884_n 0.00176486f $X=2.705 $Y=2.245 $X2=0
+ $Y2=0
cc_464 N_DE_c_500_n N_VPWR_c_1993_n 0.00154956f $X=2.025 $Y=2.245 $X2=0 $Y2=0
cc_465 N_DE_c_502_n N_VPWR_c_1993_n 0.00971267f $X=2.705 $Y=2.245 $X2=0 $Y2=0
cc_466 N_DE_c_500_n N_VPWR_c_2002_n 0.00278227f $X=2.025 $Y=2.245 $X2=0 $Y2=0
cc_467 N_DE_c_502_n N_VPWR_c_2003_n 0.00413917f $X=2.705 $Y=2.245 $X2=0 $Y2=0
cc_468 N_DE_c_500_n N_VPWR_c_1991_n 0.00360419f $X=2.025 $Y=2.245 $X2=0 $Y2=0
cc_469 N_DE_c_502_n N_VPWR_c_1991_n 0.00416568f $X=2.705 $Y=2.245 $X2=0 $Y2=0
cc_470 N_DE_M1014_g N_VGND_c_2397_n 0.0142649f $X=1.1 $Y=0.66 $X2=0 $Y2=0
cc_471 N_DE_c_492_n N_VGND_c_2397_n 0.00444518f $X=1.755 $Y=1.135 $X2=0 $Y2=0
cc_472 N_DE_c_494_n N_VGND_c_2397_n 0.00346209f $X=2.09 $Y=1.06 $X2=0 $Y2=0
cc_473 N_DE_c_494_n N_VGND_c_2398_n 0.00564371f $X=2.09 $Y=1.06 $X2=0 $Y2=0
cc_474 N_DE_c_494_n N_VGND_c_2405_n 0.00430863f $X=2.09 $Y=1.06 $X2=0 $Y2=0
cc_475 N_DE_M1014_g N_VGND_c_2409_n 0.00432588f $X=1.1 $Y=0.66 $X2=0 $Y2=0
cc_476 N_DE_M1014_g N_VGND_c_2416_n 0.00437282f $X=1.1 $Y=0.66 $X2=0 $Y2=0
cc_477 N_DE_c_494_n N_VGND_c_2416_n 0.00486331f $X=2.09 $Y=1.06 $X2=0 $Y2=0
cc_478 N_A_575_305#_M1001_g N_A_667_87#_c_836_n 0.0180128f $X=2.98 $Y=0.775
+ $X2=0 $Y2=0
cc_479 N_A_575_305#_c_601_n N_A_667_87#_c_843_n 0.00280225f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_480 N_A_575_305#_c_601_n N_A_667_87#_c_840_n 0.00539163f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_481 N_A_575_305#_c_601_n N_A_667_87#_c_846_n 0.0661871f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_482 N_A_575_305#_c_601_n N_A_667_87#_c_847_n 0.0239171f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_483 N_A_575_305#_c_601_n N_A_667_87#_c_848_n 0.00197697f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_484 N_A_575_305#_c_601_n N_A_667_87#_c_849_n 0.0209494f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_485 N_A_575_305#_c_601_n SCD 0.00362617f $X=14.015 $Y=2.035 $X2=0 $Y2=0
cc_486 N_A_575_305#_c_595_n N_SCE_c_978_n 0.00819052f $X=3.125 $Y=2.245
+ $X2=-0.19 $Y2=-0.245
cc_487 N_A_575_305#_c_601_n N_SCE_c_978_n 0.00310516f $X=14.015 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_488 N_A_575_305#_c_595_n N_SCE_c_980_n 0.00291704f $X=3.125 $Y=2.245 $X2=0
+ $Y2=0
cc_489 N_A_575_305#_c_601_n N_SCE_c_977_n 0.00291605f $X=14.015 $Y=2.035 $X2=0
+ $Y2=0
cc_490 N_A_575_305#_c_601_n N_CLK_c_1052_n 0.00513336f $X=14.015 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_491 N_A_575_305#_c_601_n CLK 0.00676205f $X=14.015 $Y=2.035 $X2=0 $Y2=0
cc_492 N_A_575_305#_c_596_n N_A_1549_74#_c_1112_n 0.0202366f $X=13.58 $Y=2.465
+ $X2=0 $Y2=0
cc_493 N_A_575_305#_c_601_n N_A_1549_74#_c_1112_n 0.00258366f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_494 N_A_575_305#_c_606_n N_A_1549_74#_c_1112_n 0.0010662f $X=14.045 $Y=2.15
+ $X2=0 $Y2=0
cc_495 N_A_575_305#_c_596_n N_A_1549_74#_c_1114_n 0.032099f $X=13.58 $Y=2.465
+ $X2=0 $Y2=0
cc_496 N_A_575_305#_c_581_n N_A_1549_74#_c_1088_n 0.0173353f $X=13.68 $Y=2.05
+ $X2=0 $Y2=0
cc_497 N_A_575_305#_c_601_n N_A_1549_74#_c_1088_n 0.00102022f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_498 N_A_575_305#_c_601_n N_A_1549_74#_c_1116_n 0.0543228f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_499 N_A_575_305#_c_601_n N_A_1549_74#_c_1101_n 0.00978658f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_500 N_A_575_305#_c_601_n N_A_1549_74#_c_1119_n 0.0040034f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_501 N_A_575_305#_c_580_n N_A_1549_74#_c_1107_n 0.00221728f $X=13.215 $Y=0.94
+ $X2=0 $Y2=0
cc_502 N_A_575_305#_c_581_n N_A_1549_74#_c_1107_n 0.0029915f $X=13.68 $Y=2.05
+ $X2=0 $Y2=0
cc_503 N_A_575_305#_c_601_n N_A_1549_74#_c_1107_n 9.44933e-19 $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_504 N_A_575_305#_c_580_n N_A_1549_74#_c_1108_n 0.0204694f $X=13.215 $Y=0.94
+ $X2=0 $Y2=0
cc_505 N_A_575_305#_c_581_n N_A_1549_74#_c_1108_n 0.0194145f $X=13.68 $Y=2.05
+ $X2=0 $Y2=0
cc_506 N_A_575_305#_c_601_n N_A_1549_74#_c_1110_n 0.00172851f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_507 N_A_575_305#_c_601_n N_A_1348_368#_c_1333_n 0.00381185f $X=14.015
+ $Y=2.035 $X2=0 $Y2=0
cc_508 N_A_575_305#_c_601_n N_A_1348_368#_c_1336_n 0.00190774f $X=14.015
+ $Y=2.035 $X2=0 $Y2=0
cc_509 N_A_575_305#_c_601_n N_A_1348_368#_c_1322_n 0.0106455f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_510 N_A_575_305#_c_578_n N_A_1348_368#_M1031_g 0.0416832f $X=13.14 $Y=0.865
+ $X2=0 $Y2=0
cc_511 N_A_575_305#_c_601_n N_A_1348_368#_c_1324_n 0.00438916f $X=14.015
+ $Y=2.035 $X2=0 $Y2=0
cc_512 N_A_575_305#_c_601_n N_A_1348_368#_c_1326_n 0.00602409f $X=14.015
+ $Y=2.035 $X2=0 $Y2=0
cc_513 N_A_575_305#_c_601_n N_A_1348_368#_c_1330_n 8.85056e-19 $X=14.015
+ $Y=2.035 $X2=0 $Y2=0
cc_514 N_A_575_305#_c_601_n N_A_1348_368#_c_1341_n 0.0362769f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_515 N_A_575_305#_c_601_n N_A_1348_368#_c_1343_n 0.0711397f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_516 N_A_575_305#_c_601_n N_A_1348_368#_c_1345_n 0.019653f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_517 N_A_575_305#_c_601_n N_A_1348_368#_c_1346_n 0.00127491f $X=14.015
+ $Y=2.035 $X2=0 $Y2=0
cc_518 N_A_575_305#_c_601_n N_A_1348_368#_c_1347_n 0.0166748f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_519 N_A_575_305#_c_601_n N_A_1348_368#_c_1348_n 0.0291663f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_520 N_A_575_305#_c_601_n N_A_1348_368#_c_1331_n 0.0121876f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_521 N_A_575_305#_c_601_n N_A_1972_92#_c_1517_n 0.0061219f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_522 N_A_575_305#_c_601_n N_A_1972_92#_c_1532_n 0.0097408f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_523 N_A_575_305#_c_601_n N_A_1972_92#_c_1521_n 0.00565189f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_524 N_A_575_305#_c_601_n N_A_1972_92#_c_1533_n 0.0161369f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_525 N_A_575_305#_c_601_n N_A_1972_92#_c_1523_n 0.016096f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_526 N_A_575_305#_c_601_n N_A_1972_92#_c_1524_n 0.021913f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_527 N_A_575_305#_c_601_n N_A_1972_92#_c_1525_n 0.0104459f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_528 N_A_575_305#_c_601_n N_A_1747_118#_c_1623_n 0.01184f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_529 N_A_575_305#_c_601_n N_A_1747_118#_c_1631_n 0.0148605f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_530 N_A_575_305#_c_601_n N_A_1747_118#_c_1632_n 0.00582607f $X=14.015
+ $Y=2.035 $X2=0 $Y2=0
cc_531 N_A_575_305#_c_601_n N_A_1747_118#_c_1627_n 0.00930916f $X=14.015
+ $Y=2.035 $X2=0 $Y2=0
cc_532 N_A_575_305#_c_601_n N_A_1747_118#_c_1628_n 0.0243404f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_533 N_A_575_305#_c_601_n N_A_2463_74#_M1030_d 0.0116805f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_534 N_A_575_305#_c_579_n N_A_2463_74#_M1028_g 0.0111968f $X=13.605 $Y=0.94
+ $X2=0 $Y2=0
cc_535 N_A_575_305#_c_584_n N_A_2463_74#_M1028_g 0.0103147f $X=14.37 $Y=0.515
+ $X2=0 $Y2=0
cc_536 N_A_575_305#_c_585_n N_A_2463_74#_M1028_g 0.00374816f $X=14.515 $Y=1.92
+ $X2=0 $Y2=0
cc_537 N_A_575_305#_c_587_n N_A_2463_74#_M1028_g 0.00469426f $X=14.6 $Y=0.34
+ $X2=0 $Y2=0
cc_538 N_A_575_305#_c_591_n N_A_2463_74#_M1028_g 0.0035022f $X=14.402 $Y=1.03
+ $X2=0 $Y2=0
cc_539 N_A_575_305#_c_581_n N_A_2463_74#_c_1715_n 0.00777741f $X=13.68 $Y=2.05
+ $X2=0 $Y2=0
cc_540 N_A_575_305#_c_596_n N_A_2463_74#_c_1727_n 0.0225784f $X=13.58 $Y=2.465
+ $X2=0 $Y2=0
cc_541 N_A_575_305#_c_581_n N_A_2463_74#_c_1727_n 0.00400974f $X=13.68 $Y=2.05
+ $X2=0 $Y2=0
cc_542 N_A_575_305#_c_585_n N_A_2463_74#_c_1727_n 0.00132461f $X=14.515 $Y=1.92
+ $X2=0 $Y2=0
cc_543 N_A_575_305#_c_600_n N_A_2463_74#_c_1727_n 0.00666912f $X=14.515 $Y=2.46
+ $X2=0 $Y2=0
cc_544 N_A_575_305#_c_603_n N_A_2463_74#_c_1727_n 0.00296683f $X=14.16 $Y=2.035
+ $X2=0 $Y2=0
cc_545 N_A_575_305#_c_607_n N_A_2463_74#_c_1727_n 0.0268318f $X=14.515 $Y=2.105
+ $X2=0 $Y2=0
cc_546 N_A_575_305#_c_585_n N_A_2463_74#_c_1716_n 0.0139245f $X=14.515 $Y=1.92
+ $X2=0 $Y2=0
cc_547 N_A_575_305#_c_607_n N_A_2463_74#_c_1716_n 2.69573e-19 $X=14.515 $Y=2.105
+ $X2=0 $Y2=0
cc_548 N_A_575_305#_c_581_n N_A_2463_74#_c_1717_n 0.021392f $X=13.68 $Y=2.05
+ $X2=0 $Y2=0
cc_549 N_A_575_305#_c_585_n N_A_2463_74#_c_1717_n 0.0146711f $X=14.515 $Y=1.92
+ $X2=0 $Y2=0
cc_550 N_A_575_305#_c_591_n N_A_2463_74#_c_1717_n 0.00899313f $X=14.402 $Y=1.03
+ $X2=0 $Y2=0
cc_551 N_A_575_305#_c_601_n N_A_2463_74#_c_1717_n 0.00102393f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_552 N_A_575_305#_c_603_n N_A_2463_74#_c_1717_n 0.00459808f $X=14.16 $Y=2.035
+ $X2=0 $Y2=0
cc_553 N_A_575_305#_c_606_n N_A_2463_74#_c_1717_n 0.00128335f $X=14.045 $Y=2.15
+ $X2=0 $Y2=0
cc_554 N_A_575_305#_c_607_n N_A_2463_74#_c_1717_n 0.00322154f $X=14.515 $Y=2.105
+ $X2=0 $Y2=0
cc_555 N_A_575_305#_M1000_g N_A_2463_74#_c_1718_n 0.00996638f $X=15.825 $Y=0.76
+ $X2=0 $Y2=0
cc_556 N_A_575_305#_c_584_n N_A_2463_74#_c_1718_n 0.00448058f $X=14.37 $Y=0.515
+ $X2=0 $Y2=0
cc_557 N_A_575_305#_c_586_n N_A_2463_74#_c_1718_n 0.0152762f $X=15.185 $Y=0.34
+ $X2=0 $Y2=0
cc_558 N_A_575_305#_c_588_n N_A_2463_74#_c_1718_n 0.0198565f $X=15.27 $Y=1.32
+ $X2=0 $Y2=0
cc_559 N_A_575_305#_c_582_n N_A_2463_74#_c_1719_n 0.0213458f $X=15.8 $Y=1.765
+ $X2=0 $Y2=0
cc_560 N_A_575_305#_M1000_g N_A_2463_74#_c_1719_n 0.00402418f $X=15.825 $Y=0.76
+ $X2=0 $Y2=0
cc_561 N_A_575_305#_c_588_n N_A_2463_74#_c_1719_n 0.00836309f $X=15.27 $Y=1.32
+ $X2=0 $Y2=0
cc_562 N_A_575_305#_c_589_n N_A_2463_74#_c_1719_n 0.00105406f $X=15.355 $Y=1.485
+ $X2=0 $Y2=0
cc_563 N_A_575_305#_c_590_n N_A_2463_74#_c_1719_n 0.00181641f $X=15.765 $Y=1.485
+ $X2=0 $Y2=0
cc_564 N_A_575_305#_c_582_n N_A_2463_74#_c_1720_n 0.00450965f $X=15.8 $Y=1.765
+ $X2=0 $Y2=0
cc_565 N_A_575_305#_c_589_n N_A_2463_74#_c_1720_n 0.0145902f $X=15.355 $Y=1.485
+ $X2=0 $Y2=0
cc_566 N_A_575_305#_c_590_n N_A_2463_74#_c_1720_n 0.00509302f $X=15.765 $Y=1.485
+ $X2=0 $Y2=0
cc_567 N_A_575_305#_c_582_n N_A_2463_74#_c_1729_n 0.0207548f $X=15.8 $Y=1.765
+ $X2=0 $Y2=0
cc_568 N_A_575_305#_c_600_n N_A_2463_74#_c_1729_n 9.02283e-19 $X=14.515 $Y=2.46
+ $X2=0 $Y2=0
cc_569 N_A_575_305#_c_607_n N_A_2463_74#_c_1729_n 9.00246e-19 $X=14.515 $Y=2.105
+ $X2=0 $Y2=0
cc_570 N_A_575_305#_c_578_n N_A_2463_74#_c_1722_n 0.00748201f $X=13.14 $Y=0.865
+ $X2=0 $Y2=0
cc_571 N_A_575_305#_c_579_n N_A_2463_74#_c_1722_n 0.0264434f $X=13.605 $Y=0.94
+ $X2=0 $Y2=0
cc_572 N_A_575_305#_c_580_n N_A_2463_74#_c_1722_n 0.00284486f $X=13.215 $Y=0.94
+ $X2=0 $Y2=0
cc_573 N_A_575_305#_c_584_n N_A_2463_74#_c_1722_n 0.00851476f $X=14.37 $Y=0.515
+ $X2=0 $Y2=0
cc_574 N_A_575_305#_c_596_n N_A_2463_74#_c_1730_n 0.00128259f $X=13.58 $Y=2.465
+ $X2=0 $Y2=0
cc_575 N_A_575_305#_c_581_n N_A_2463_74#_c_1730_n 0.00107747f $X=13.68 $Y=2.05
+ $X2=0 $Y2=0
cc_576 N_A_575_305#_c_601_n N_A_2463_74#_c_1730_n 0.015003f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_577 N_A_575_305#_c_606_n N_A_2463_74#_c_1730_n 0.0165122f $X=14.045 $Y=2.15
+ $X2=0 $Y2=0
cc_578 N_A_575_305#_c_596_n N_A_2463_74#_c_1731_n 0.00326298f $X=13.58 $Y=2.465
+ $X2=0 $Y2=0
cc_579 N_A_575_305#_c_581_n N_A_2463_74#_c_1731_n 0.0127392f $X=13.68 $Y=2.05
+ $X2=0 $Y2=0
cc_580 N_A_575_305#_c_585_n N_A_2463_74#_c_1731_n 0.00624801f $X=14.515 $Y=1.92
+ $X2=0 $Y2=0
cc_581 N_A_575_305#_c_601_n N_A_2463_74#_c_1731_n 0.0237956f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_582 N_A_575_305#_c_606_n N_A_2463_74#_c_1731_n 0.0261817f $X=14.045 $Y=2.15
+ $X2=0 $Y2=0
cc_583 N_A_575_305#_c_579_n N_A_2463_74#_c_1723_n 0.00406672f $X=13.605 $Y=0.94
+ $X2=0 $Y2=0
cc_584 N_A_575_305#_c_581_n N_A_2463_74#_c_1723_n 0.00750619f $X=13.68 $Y=2.05
+ $X2=0 $Y2=0
cc_585 N_A_575_305#_c_585_n N_A_2463_74#_c_1723_n 0.00556876f $X=14.515 $Y=1.92
+ $X2=0 $Y2=0
cc_586 N_A_575_305#_c_591_n N_A_2463_74#_c_1723_n 0.00405365f $X=14.402 $Y=1.03
+ $X2=0 $Y2=0
cc_587 N_A_575_305#_c_581_n N_A_2463_74#_c_1724_n 0.00557048f $X=13.68 $Y=2.05
+ $X2=0 $Y2=0
cc_588 N_A_575_305#_c_585_n N_A_2463_74#_c_1724_n 0.0060599f $X=14.515 $Y=1.92
+ $X2=0 $Y2=0
cc_589 N_A_575_305#_c_596_n N_A_2463_74#_c_1734_n 0.00185207f $X=13.58 $Y=2.465
+ $X2=0 $Y2=0
cc_590 N_A_575_305#_c_601_n N_A_2463_74#_c_1734_n 0.0108136f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_591 N_A_575_305#_c_581_n N_A_2463_74#_c_1725_n 0.00812064f $X=13.68 $Y=2.05
+ $X2=0 $Y2=0
cc_592 N_A_575_305#_c_585_n N_A_2463_74#_c_1725_n 0.0252289f $X=14.515 $Y=1.92
+ $X2=0 $Y2=0
cc_593 N_A_575_305#_c_591_n N_A_2463_74#_c_1725_n 0.00444579f $X=14.402 $Y=1.03
+ $X2=0 $Y2=0
cc_594 N_A_575_305#_c_601_n N_A_2463_74#_c_1725_n 0.00315435f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_595 N_A_575_305#_c_603_n N_A_2463_74#_c_1725_n 0.00568398f $X=14.16 $Y=2.035
+ $X2=0 $Y2=0
cc_596 N_A_575_305#_c_606_n N_A_2463_74#_c_1725_n 0.0032606f $X=14.045 $Y=2.15
+ $X2=0 $Y2=0
cc_597 N_A_575_305#_c_607_n N_A_2463_74#_c_1725_n 0.00580451f $X=14.515 $Y=2.105
+ $X2=0 $Y2=0
cc_598 N_A_575_305#_c_595_n N_A_27_90#_c_1880_n 0.00934852f $X=3.125 $Y=2.245
+ $X2=0 $Y2=0
cc_599 N_A_575_305#_c_602_n N_A_27_90#_c_1880_n 0.00519233f $X=3.265 $Y=2.035
+ $X2=0 $Y2=0
cc_600 N_A_575_305#_c_592_n N_A_27_90#_c_1880_n 5.90449e-19 $X=3.04 $Y=1.69
+ $X2=0 $Y2=0
cc_601 N_A_575_305#_c_593_n N_A_27_90#_c_1880_n 0.0214452f $X=3.04 $Y=1.69 $X2=0
+ $Y2=0
cc_602 N_A_575_305#_M1001_g N_A_27_90#_c_1870_n 0.0138821f $X=2.98 $Y=0.775
+ $X2=0 $Y2=0
cc_603 N_A_575_305#_M1001_g N_A_27_90#_c_1871_n 0.00523715f $X=2.98 $Y=0.775
+ $X2=0 $Y2=0
cc_604 N_A_575_305#_c_595_n N_A_27_90#_c_1871_n 0.00132884f $X=3.125 $Y=2.245
+ $X2=0 $Y2=0
cc_605 N_A_575_305#_c_601_n N_A_27_90#_c_1871_n 0.0222045f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_606 N_A_575_305#_c_602_n N_A_27_90#_c_1871_n 0.00296683f $X=3.265 $Y=2.035
+ $X2=0 $Y2=0
cc_607 N_A_575_305#_c_592_n N_A_27_90#_c_1871_n 0.015199f $X=3.04 $Y=1.69 $X2=0
+ $Y2=0
cc_608 N_A_575_305#_c_593_n N_A_27_90#_c_1871_n 0.0441454f $X=3.04 $Y=1.69 $X2=0
+ $Y2=0
cc_609 N_A_575_305#_M1001_g N_A_27_90#_c_1873_n 0.0069713f $X=2.98 $Y=0.775
+ $X2=0 $Y2=0
cc_610 N_A_575_305#_c_602_n N_A_27_90#_c_1873_n 0.00254272f $X=3.265 $Y=2.035
+ $X2=0 $Y2=0
cc_611 N_A_575_305#_c_592_n N_A_27_90#_c_1873_n 0.00147548f $X=3.04 $Y=1.69
+ $X2=0 $Y2=0
cc_612 N_A_575_305#_c_593_n N_A_27_90#_c_1873_n 0.0127272f $X=3.04 $Y=1.69 $X2=0
+ $Y2=0
cc_613 N_A_575_305#_c_595_n N_A_27_90#_c_1884_n 0.0101556f $X=3.125 $Y=2.245
+ $X2=0 $Y2=0
cc_614 N_A_575_305#_c_601_n N_A_27_90#_c_1884_n 0.00556493f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_615 N_A_575_305#_c_602_n N_A_27_90#_c_1884_n 0.00380336f $X=3.265 $Y=2.035
+ $X2=0 $Y2=0
cc_616 N_A_575_305#_c_593_n N_A_27_90#_c_1884_n 0.00129625f $X=3.04 $Y=1.69
+ $X2=0 $Y2=0
cc_617 N_A_575_305#_c_601_n N_VPWR_M1034_s 0.0137059f $X=14.015 $Y=2.035 $X2=0
+ $Y2=0
cc_618 N_A_575_305#_c_601_n N_VPWR_M1008_s 0.00279283f $X=14.015 $Y=2.035 $X2=0
+ $Y2=0
cc_619 N_A_575_305#_c_601_n N_VPWR_M1041_d 0.00247486f $X=14.015 $Y=2.035 $X2=0
+ $Y2=0
cc_620 N_A_575_305#_c_601_n N_VPWR_M1038_s 0.00857475f $X=14.015 $Y=2.035 $X2=0
+ $Y2=0
cc_621 N_A_575_305#_c_601_n N_VPWR_M1039_d 6.98211e-19 $X=14.015 $Y=2.035 $X2=0
+ $Y2=0
cc_622 N_A_575_305#_c_606_n N_VPWR_M1039_d 0.0035033f $X=14.045 $Y=2.15 $X2=0
+ $Y2=0
cc_623 N_A_575_305#_c_607_n N_VPWR_M1039_d 0.00315433f $X=14.515 $Y=2.105 $X2=0
+ $Y2=0
cc_624 N_A_575_305#_c_595_n N_VPWR_c_1993_n 0.00149818f $X=3.125 $Y=2.245 $X2=0
+ $Y2=0
cc_625 N_A_575_305#_c_601_n N_VPWR_c_1996_n 9.24589e-19 $X=14.015 $Y=2.035 $X2=0
+ $Y2=0
cc_626 N_A_575_305#_c_596_n N_VPWR_c_1999_n 0.01866f $X=13.58 $Y=2.465 $X2=0
+ $Y2=0
cc_627 N_A_575_305#_c_600_n N_VPWR_c_1999_n 0.0225324f $X=14.515 $Y=2.46 $X2=0
+ $Y2=0
cc_628 N_A_575_305#_c_601_n N_VPWR_c_1999_n 0.00193253f $X=14.015 $Y=2.035 $X2=0
+ $Y2=0
cc_629 N_A_575_305#_c_603_n N_VPWR_c_1999_n 0.00116543f $X=14.16 $Y=2.035 $X2=0
+ $Y2=0
cc_630 N_A_575_305#_c_606_n N_VPWR_c_1999_n 0.0275703f $X=14.045 $Y=2.15 $X2=0
+ $Y2=0
cc_631 N_A_575_305#_c_582_n N_VPWR_c_2000_n 0.0113451f $X=15.8 $Y=1.765 $X2=0
+ $Y2=0
cc_632 N_A_575_305#_c_590_n N_VPWR_c_2000_n 0.0215711f $X=15.765 $Y=1.485 $X2=0
+ $Y2=0
cc_633 N_A_575_305#_c_595_n N_VPWR_c_2003_n 0.00445602f $X=3.125 $Y=2.245 $X2=0
+ $Y2=0
cc_634 N_A_575_305#_c_596_n N_VPWR_c_2008_n 0.00413917f $X=13.58 $Y=2.465 $X2=0
+ $Y2=0
cc_635 N_A_575_305#_c_600_n N_VPWR_c_2009_n 0.00742834f $X=14.515 $Y=2.46 $X2=0
+ $Y2=0
cc_636 N_A_575_305#_c_582_n N_VPWR_c_2010_n 0.00445602f $X=15.8 $Y=1.765 $X2=0
+ $Y2=0
cc_637 N_A_575_305#_c_595_n N_VPWR_c_1991_n 0.00455473f $X=3.125 $Y=2.245 $X2=0
+ $Y2=0
cc_638 N_A_575_305#_c_596_n N_VPWR_c_1991_n 0.00852225f $X=13.58 $Y=2.465 $X2=0
+ $Y2=0
cc_639 N_A_575_305#_c_582_n N_VPWR_c_1991_n 0.00860975f $X=15.8 $Y=1.765 $X2=0
+ $Y2=0
cc_640 N_A_575_305#_c_600_n N_VPWR_c_1991_n 0.00617854f $X=14.515 $Y=2.46 $X2=0
+ $Y2=0
cc_641 N_A_575_305#_c_601_n N_A_697_113#_c_2180_n 0.00405912f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_642 N_A_575_305#_c_601_n N_A_697_113#_c_2184_n 0.00136998f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_643 N_A_575_305#_c_601_n N_A_697_113#_c_2173_n 0.0180895f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_644 N_A_575_305#_c_601_n N_A_697_113#_c_2186_n 0.0381577f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_645 N_A_575_305#_c_601_n N_A_697_113#_c_2187_n 0.0143788f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_646 N_A_575_305#_c_601_n N_A_697_113#_c_2174_n 0.00605249f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_647 N_A_575_305#_c_601_n N_A_697_113#_c_2200_n 0.00613078f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_648 N_A_575_305#_M1001_g N_A_697_113#_c_2178_n 6.24512e-19 $X=2.98 $Y=0.775
+ $X2=0 $Y2=0
cc_649 N_A_575_305#_c_601_n N_A_697_113#_c_2178_n 0.0234101f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_650 N_A_575_305#_c_601_n N_A_697_113#_c_2192_n 0.0079778f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_651 N_A_575_305#_c_601_n N_A_697_113#_c_2193_n 0.00847007f $X=14.015 $Y=2.035
+ $X2=0 $Y2=0
cc_652 N_A_575_305#_c_601_n A_2345_392# 0.024037f $X=14.015 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_653 N_A_575_305#_c_586_n N_Q_M1036_s 0.00440738f $X=15.185 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_654 N_A_575_305#_c_584_n N_Q_c_2349_n 0.0379556f $X=14.37 $Y=0.515 $X2=0
+ $Y2=0
cc_655 N_A_575_305#_c_586_n N_Q_c_2349_n 0.0112956f $X=15.185 $Y=0.34 $X2=0
+ $Y2=0
cc_656 N_A_575_305#_c_588_n N_Q_c_2349_n 0.0303369f $X=15.27 $Y=1.32 $X2=0 $Y2=0
cc_657 N_A_575_305#_c_589_n N_Q_c_2349_n 0.0276767f $X=15.355 $Y=1.485 $X2=0
+ $Y2=0
cc_658 N_A_575_305#_c_589_n Q 0.00486469f $X=15.355 $Y=1.485 $X2=0 $Y2=0
cc_659 N_A_575_305#_c_591_n Q 0.0379556f $X=14.402 $Y=1.03 $X2=0 $Y2=0
cc_660 N_A_575_305#_c_603_n Q 0.00102695f $X=14.16 $Y=2.035 $X2=0 $Y2=0
cc_661 N_A_575_305#_c_607_n Q 0.0297348f $X=14.515 $Y=2.105 $X2=0 $Y2=0
cc_662 N_A_575_305#_c_600_n Q 0.0365671f $X=14.515 $Y=2.46 $X2=0 $Y2=0
cc_663 N_A_575_305#_M1000_g N_Q_N_c_2375_n 0.00827903f $X=15.825 $Y=0.76 $X2=0
+ $Y2=0
cc_664 N_A_575_305#_c_582_n N_Q_N_c_2376_n 9.04951e-19 $X=15.8 $Y=1.765 $X2=0
+ $Y2=0
cc_665 N_A_575_305#_M1000_g N_Q_N_c_2376_n 0.0027199f $X=15.825 $Y=0.76 $X2=0
+ $Y2=0
cc_666 N_A_575_305#_c_590_n N_Q_N_c_2376_n 0.00151667f $X=15.765 $Y=1.485 $X2=0
+ $Y2=0
cc_667 N_A_575_305#_c_582_n Q_N 0.00406669f $X=15.8 $Y=1.765 $X2=0 $Y2=0
cc_668 N_A_575_305#_c_590_n Q_N 0.00280403f $X=15.765 $Y=1.485 $X2=0 $Y2=0
cc_669 N_A_575_305#_c_582_n Q_N 0.0108562f $X=15.8 $Y=1.765 $X2=0 $Y2=0
cc_670 N_A_575_305#_c_582_n N_Q_N_c_2377_n 0.0118858f $X=15.8 $Y=1.765 $X2=0
+ $Y2=0
cc_671 N_A_575_305#_M1000_g N_Q_N_c_2377_n 0.00411368f $X=15.825 $Y=0.76 $X2=0
+ $Y2=0
cc_672 N_A_575_305#_c_590_n N_Q_N_c_2377_n 0.0263023f $X=15.765 $Y=1.485 $X2=0
+ $Y2=0
cc_673 N_A_575_305#_c_586_n N_VGND_M1036_d 3.32641e-19 $X=15.185 $Y=0.34 $X2=0
+ $Y2=0
cc_674 N_A_575_305#_c_588_n N_VGND_M1036_d 0.0064283f $X=15.27 $Y=1.32 $X2=0
+ $Y2=0
cc_675 N_A_575_305#_M1001_g N_VGND_c_2398_n 0.0018473f $X=2.98 $Y=0.775 $X2=0
+ $Y2=0
cc_676 N_A_575_305#_c_582_n N_VGND_c_2404_n 0.00218979f $X=15.8 $Y=1.765 $X2=0
+ $Y2=0
cc_677 N_A_575_305#_M1000_g N_VGND_c_2404_n 0.00378095f $X=15.825 $Y=0.76 $X2=0
+ $Y2=0
cc_678 N_A_575_305#_c_586_n N_VGND_c_2404_n 0.0142487f $X=15.185 $Y=0.34 $X2=0
+ $Y2=0
cc_679 N_A_575_305#_c_588_n N_VGND_c_2404_n 0.0526757f $X=15.27 $Y=1.32 $X2=0
+ $Y2=0
cc_680 N_A_575_305#_c_590_n N_VGND_c_2404_n 0.0144735f $X=15.765 $Y=1.485 $X2=0
+ $Y2=0
cc_681 N_A_575_305#_M1001_g N_VGND_c_2410_n 0.00430863f $X=2.98 $Y=0.775 $X2=0
+ $Y2=0
cc_682 N_A_575_305#_c_586_n N_VGND_c_2414_n 0.0498132f $X=15.185 $Y=0.34 $X2=0
+ $Y2=0
cc_683 N_A_575_305#_c_587_n N_VGND_c_2414_n 0.0282284f $X=14.6 $Y=0.34 $X2=0
+ $Y2=0
cc_684 N_A_575_305#_M1000_g N_VGND_c_2415_n 0.00537471f $X=15.825 $Y=0.76 $X2=0
+ $Y2=0
cc_685 N_A_575_305#_M1001_g N_VGND_c_2416_n 0.00486331f $X=2.98 $Y=0.775 $X2=0
+ $Y2=0
cc_686 N_A_575_305#_c_578_n N_VGND_c_2416_n 0.00367447f $X=13.14 $Y=0.865 $X2=0
+ $Y2=0
cc_687 N_A_575_305#_M1000_g N_VGND_c_2416_n 0.00539454f $X=15.825 $Y=0.76 $X2=0
+ $Y2=0
cc_688 N_A_575_305#_c_586_n N_VGND_c_2416_n 0.0285959f $X=15.185 $Y=0.34 $X2=0
+ $Y2=0
cc_689 N_A_575_305#_c_587_n N_VGND_c_2416_n 0.0152423f $X=14.6 $Y=0.34 $X2=0
+ $Y2=0
cc_690 N_A_575_305#_c_578_n N_VGND_c_2422_n 0.00383152f $X=13.14 $Y=0.865 $X2=0
+ $Y2=0
cc_691 N_A_575_305#_c_578_n N_VGND_c_2423_n 0.0105517f $X=13.14 $Y=0.865 $X2=0
+ $Y2=0
cc_692 N_A_575_305#_c_579_n N_VGND_c_2423_n 0.00323484f $X=13.605 $Y=0.94 $X2=0
+ $Y2=0
cc_693 N_A_575_305#_c_587_n N_VGND_c_2423_n 0.0125324f $X=14.6 $Y=0.34 $X2=0
+ $Y2=0
cc_694 N_A_667_87#_c_843_n N_SCD_c_927_n 0.0289443f $X=5.655 $Y=2.235 $X2=0
+ $Y2=0
cc_695 N_A_667_87#_c_846_n N_SCD_c_927_n 0.0135349f $X=5.565 $Y=2.035 $X2=0
+ $Y2=0
cc_696 N_A_667_87#_c_849_n N_SCD_c_927_n 0.00119951f $X=5.73 $Y=1.955 $X2=0
+ $Y2=0
cc_697 N_A_667_87#_c_843_n N_SCD_c_932_n 0.043976f $X=5.655 $Y=2.235 $X2=0 $Y2=0
cc_698 N_A_667_87#_c_842_n N_SCD_M1024_g 3.61896e-19 $X=4.18 $Y=0.737 $X2=0
+ $Y2=0
cc_699 N_A_667_87#_c_843_n SCD 4.20387e-19 $X=5.655 $Y=2.235 $X2=0 $Y2=0
cc_700 N_A_667_87#_c_846_n SCD 0.0145726f $X=5.565 $Y=2.035 $X2=0 $Y2=0
cc_701 N_A_667_87#_c_849_n SCD 0.00333536f $X=5.73 $Y=1.955 $X2=0 $Y2=0
cc_702 N_A_667_87#_c_846_n N_SCD_c_930_n 0.00281188f $X=5.565 $Y=2.035 $X2=0
+ $Y2=0
cc_703 N_A_667_87#_c_848_n N_SCE_c_979_n 0.00173288f $X=4.36 $Y=2.51 $X2=0 $Y2=0
cc_704 N_A_667_87#_c_867_p N_SCE_c_981_n 0.00107941f $X=4.155 $Y=1.255 $X2=0
+ $Y2=0
cc_705 N_A_667_87#_c_840_n N_SCE_c_981_n 0.0178405f $X=4.155 $Y=1.255 $X2=0
+ $Y2=0
cc_706 N_A_667_87#_c_845_n N_SCE_c_981_n 0.00363753f $X=4.22 $Y=2.29 $X2=0 $Y2=0
cc_707 N_A_667_87#_c_846_n N_SCE_c_981_n 0.0139476f $X=5.565 $Y=2.035 $X2=0
+ $Y2=0
cc_708 N_A_667_87#_c_845_n N_SCE_M1003_g 0.00167654f $X=4.22 $Y=2.29 $X2=0 $Y2=0
cc_709 N_A_667_87#_c_848_n N_SCE_M1003_g 0.00903043f $X=4.36 $Y=2.51 $X2=0 $Y2=0
cc_710 N_A_667_87#_c_867_p N_SCE_M1037_g 0.00215718f $X=4.155 $Y=1.255 $X2=0
+ $Y2=0
cc_711 N_A_667_87#_c_841_n N_SCE_M1037_g 0.0263062f $X=4.155 $Y=0.575 $X2=0
+ $Y2=0
cc_712 N_A_667_87#_c_842_n N_SCE_M1037_g 0.00823696f $X=4.18 $Y=0.737 $X2=0
+ $Y2=0
cc_713 N_A_667_87#_c_843_n N_SCE_M1010_g 0.00232566f $X=5.655 $Y=2.235 $X2=0
+ $Y2=0
cc_714 N_A_667_87#_c_849_n N_SCE_M1010_g 8.18203e-19 $X=5.73 $Y=1.955 $X2=0
+ $Y2=0
cc_715 N_A_667_87#_c_867_p N_SCE_c_976_n 3.55703e-19 $X=4.155 $Y=1.255 $X2=0
+ $Y2=0
cc_716 N_A_667_87#_c_840_n N_SCE_c_976_n 0.0199971f $X=4.155 $Y=1.255 $X2=0
+ $Y2=0
cc_717 N_A_667_87#_c_846_n N_SCE_c_976_n 0.00385557f $X=5.565 $Y=2.035 $X2=0
+ $Y2=0
cc_718 N_A_667_87#_c_842_n N_SCE_c_976_n 0.00408345f $X=4.18 $Y=0.737 $X2=0
+ $Y2=0
cc_719 N_A_667_87#_c_867_p N_SCE_c_977_n 0.0259191f $X=4.155 $Y=1.255 $X2=0
+ $Y2=0
cc_720 N_A_667_87#_c_840_n N_SCE_c_977_n 0.00196091f $X=4.155 $Y=1.255 $X2=0
+ $Y2=0
cc_721 N_A_667_87#_c_846_n N_SCE_c_977_n 0.0261529f $X=5.565 $Y=2.035 $X2=0
+ $Y2=0
cc_722 N_A_667_87#_c_842_n N_SCE_c_977_n 0.0119127f $X=4.18 $Y=0.737 $X2=0 $Y2=0
cc_723 N_A_667_87#_c_843_n N_CLK_c_1052_n 0.00400897f $X=5.655 $Y=2.235
+ $X2=-0.19 $Y2=-0.245
cc_724 N_A_667_87#_c_836_n N_A_27_90#_c_1870_n 0.0073934f $X=3.41 $Y=1.06 $X2=0
+ $Y2=0
cc_725 N_A_667_87#_c_838_n N_A_27_90#_c_1870_n 0.00413546f $X=3.485 $Y=1.135
+ $X2=0 $Y2=0
cc_726 N_A_667_87#_c_838_n N_A_27_90#_c_1871_n 9.15581e-19 $X=3.485 $Y=1.135
+ $X2=0 $Y2=0
cc_727 N_A_667_87#_c_837_n N_A_27_90#_c_1873_n 0.00384415f $X=3.99 $Y=1.135
+ $X2=0 $Y2=0
cc_728 N_A_667_87#_c_838_n N_A_27_90#_c_1873_n 0.00908768f $X=3.485 $Y=1.135
+ $X2=0 $Y2=0
cc_729 N_A_667_87#_c_843_n N_VPWR_c_1994_n 0.00149083f $X=5.655 $Y=2.235 $X2=0
+ $Y2=0
cc_730 N_A_667_87#_c_843_n N_VPWR_c_1995_n 0.00334802f $X=5.655 $Y=2.235 $X2=0
+ $Y2=0
cc_731 N_A_667_87#_c_843_n N_VPWR_c_2004_n 0.0055545f $X=5.655 $Y=2.235 $X2=0
+ $Y2=0
cc_732 N_A_667_87#_c_843_n N_VPWR_c_1991_n 0.00542671f $X=5.655 $Y=2.235 $X2=0
+ $Y2=0
cc_733 N_A_667_87#_c_848_n N_A_697_113#_c_2180_n 0.0353494f $X=4.36 $Y=2.51
+ $X2=0 $Y2=0
cc_734 N_A_667_87#_M1003_s N_A_697_113#_c_2182_n 0.00523626f $X=4.215 $Y=2.31
+ $X2=0 $Y2=0
cc_735 N_A_667_87#_c_848_n N_A_697_113#_c_2182_n 0.0229449f $X=4.36 $Y=2.51
+ $X2=0 $Y2=0
cc_736 N_A_667_87#_c_848_n N_A_697_113#_c_2208_n 0.0202406f $X=4.36 $Y=2.51
+ $X2=0 $Y2=0
cc_737 N_A_667_87#_c_846_n N_A_697_113#_c_2184_n 0.0120361f $X=5.565 $Y=2.035
+ $X2=0 $Y2=0
cc_738 N_A_667_87#_c_848_n N_A_697_113#_c_2184_n 0.0139617f $X=4.36 $Y=2.51
+ $X2=0 $Y2=0
cc_739 N_A_667_87#_c_843_n N_A_697_113#_c_2173_n 0.00844496f $X=5.655 $Y=2.235
+ $X2=0 $Y2=0
cc_740 N_A_667_87#_c_849_n N_A_697_113#_c_2173_n 0.0236965f $X=5.73 $Y=1.955
+ $X2=0 $Y2=0
cc_741 N_A_667_87#_c_836_n N_A_697_113#_c_2177_n 0.00336993f $X=3.41 $Y=1.06
+ $X2=0 $Y2=0
cc_742 N_A_667_87#_c_837_n N_A_697_113#_c_2177_n 0.00615128f $X=3.99 $Y=1.135
+ $X2=0 $Y2=0
cc_743 N_A_667_87#_c_841_n N_A_697_113#_c_2177_n 0.0053473f $X=4.155 $Y=0.575
+ $X2=0 $Y2=0
cc_744 N_A_667_87#_c_842_n N_A_697_113#_c_2177_n 0.0431718f $X=4.18 $Y=0.737
+ $X2=0 $Y2=0
cc_745 N_A_667_87#_c_836_n N_A_697_113#_c_2178_n 4.72117e-19 $X=3.41 $Y=1.06
+ $X2=0 $Y2=0
cc_746 N_A_667_87#_c_837_n N_A_697_113#_c_2178_n 0.0149877f $X=3.99 $Y=1.135
+ $X2=0 $Y2=0
cc_747 N_A_667_87#_c_867_p N_A_697_113#_c_2178_n 0.0644749f $X=4.155 $Y=1.255
+ $X2=0 $Y2=0
cc_748 N_A_667_87#_c_840_n N_A_697_113#_c_2178_n 0.0207767f $X=4.155 $Y=1.255
+ $X2=0 $Y2=0
cc_749 N_A_667_87#_c_845_n N_A_697_113#_c_2178_n 0.00975616f $X=4.22 $Y=2.29
+ $X2=0 $Y2=0
cc_750 N_A_667_87#_c_847_n N_A_697_113#_c_2178_n 0.0120785f $X=4.18 $Y=2.035
+ $X2=0 $Y2=0
cc_751 N_A_667_87#_c_848_n N_A_697_113#_c_2178_n 5.1565e-19 $X=4.36 $Y=2.51
+ $X2=0 $Y2=0
cc_752 N_A_667_87#_c_843_n N_A_697_113#_c_2191_n 0.00863242f $X=5.655 $Y=2.235
+ $X2=0 $Y2=0
cc_753 N_A_667_87#_c_843_n N_A_697_113#_c_2192_n 0.0117264f $X=5.655 $Y=2.235
+ $X2=0 $Y2=0
cc_754 N_A_667_87#_c_846_n N_A_697_113#_c_2192_n 0.0521744f $X=5.565 $Y=2.035
+ $X2=0 $Y2=0
cc_755 N_A_667_87#_c_849_n N_A_697_113#_c_2192_n 0.0203965f $X=5.73 $Y=1.955
+ $X2=0 $Y2=0
cc_756 N_A_667_87#_c_843_n N_A_697_113#_c_2193_n 0.00353126f $X=5.655 $Y=2.235
+ $X2=0 $Y2=0
cc_757 N_A_667_87#_c_842_n N_VGND_c_2399_n 0.0236355f $X=4.18 $Y=0.737 $X2=0
+ $Y2=0
cc_758 N_A_667_87#_c_836_n N_VGND_c_2410_n 0.00430863f $X=3.41 $Y=1.06 $X2=0
+ $Y2=0
cc_759 N_A_667_87#_c_841_n N_VGND_c_2410_n 0.00366457f $X=4.155 $Y=0.575 $X2=0
+ $Y2=0
cc_760 N_A_667_87#_c_842_n N_VGND_c_2410_n 0.0173208f $X=4.18 $Y=0.737 $X2=0
+ $Y2=0
cc_761 N_A_667_87#_c_836_n N_VGND_c_2416_n 0.00486331f $X=3.41 $Y=1.06 $X2=0
+ $Y2=0
cc_762 N_A_667_87#_c_841_n N_VGND_c_2416_n 0.00263234f $X=4.155 $Y=0.575 $X2=0
+ $Y2=0
cc_763 N_A_667_87#_c_842_n N_VGND_c_2416_n 0.0217755f $X=4.18 $Y=0.737 $X2=0
+ $Y2=0
cc_764 N_SCD_c_932_n N_SCE_c_979_n 0.00127273f $X=5.265 $Y=2.235 $X2=0 $Y2=0
cc_765 N_SCD_c_927_n N_SCE_c_981_n 0.00704275f $X=5.265 $Y=2.145 $X2=0 $Y2=0
cc_766 N_SCD_c_932_n N_SCE_c_982_n 0.00704275f $X=5.265 $Y=2.235 $X2=0 $Y2=0
cc_767 N_SCD_c_932_n N_SCE_M1003_g 0.0138345f $X=5.265 $Y=2.235 $X2=0 $Y2=0
cc_768 N_SCD_M1024_g N_SCE_M1037_g 0.0150301f $X=5.3 $Y=0.835 $X2=0 $Y2=0
cc_769 SCD N_SCE_M1037_g 0.00178735f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_770 N_SCD_c_930_n N_SCE_M1037_g 0.019939f $X=5.24 $Y=1.345 $X2=0 $Y2=0
cc_771 N_SCD_M1024_g N_SCE_c_973_n 0.00900015f $X=5.3 $Y=0.835 $X2=0 $Y2=0
cc_772 N_SCD_M1024_g N_SCE_M1010_g 0.0347974f $X=5.3 $Y=0.835 $X2=0 $Y2=0
cc_773 SCD N_SCE_M1010_g 7.37715e-19 $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_774 N_SCD_c_927_n N_SCE_c_976_n 0.0100242f $X=5.265 $Y=2.145 $X2=0 $Y2=0
cc_775 N_SCD_c_927_n N_SCE_c_977_n 0.00167639f $X=5.265 $Y=2.145 $X2=0 $Y2=0
cc_776 SCD N_SCE_c_977_n 0.00391033f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_777 N_SCD_c_932_n N_VPWR_c_1994_n 0.00946073f $X=5.265 $Y=2.235 $X2=0 $Y2=0
cc_778 N_SCD_c_932_n N_VPWR_c_2004_n 0.00512473f $X=5.265 $Y=2.235 $X2=0 $Y2=0
cc_779 N_SCD_c_932_n N_VPWR_c_1991_n 0.00492022f $X=5.265 $Y=2.235 $X2=0 $Y2=0
cc_780 N_SCD_c_932_n N_A_697_113#_c_2182_n 4.20814e-19 $X=5.265 $Y=2.235 $X2=0
+ $Y2=0
cc_781 N_SCD_c_932_n N_A_697_113#_c_2208_n 0.00277676f $X=5.265 $Y=2.235 $X2=0
+ $Y2=0
cc_782 N_SCD_c_927_n N_A_697_113#_c_2173_n 0.00575138f $X=5.265 $Y=2.145 $X2=0
+ $Y2=0
cc_783 N_SCD_M1024_g N_A_697_113#_c_2173_n 2.92541e-19 $X=5.3 $Y=0.835 $X2=0
+ $Y2=0
cc_784 SCD N_A_697_113#_c_2173_n 0.0149299f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_785 N_SCD_c_930_n N_A_697_113#_c_2173_n 0.0012913f $X=5.24 $Y=1.345 $X2=0
+ $Y2=0
cc_786 N_SCD_c_932_n N_A_697_113#_c_2191_n 0.00168109f $X=5.265 $Y=2.235 $X2=0
+ $Y2=0
cc_787 N_SCD_c_932_n N_A_697_113#_c_2192_n 0.01578f $X=5.265 $Y=2.235 $X2=0
+ $Y2=0
cc_788 N_SCD_M1024_g N_A_697_113#_c_2179_n 0.00114517f $X=5.3 $Y=0.835 $X2=0
+ $Y2=0
cc_789 N_SCD_M1024_g N_VGND_c_2399_n 0.0104312f $X=5.3 $Y=0.835 $X2=0 $Y2=0
cc_790 SCD N_VGND_c_2399_n 0.0109465f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_791 N_SCD_c_930_n N_VGND_c_2399_n 0.00351787f $X=5.24 $Y=1.345 $X2=0 $Y2=0
cc_792 N_SCD_M1024_g N_VGND_c_2416_n 8.6132e-19 $X=5.3 $Y=0.835 $X2=0 $Y2=0
cc_793 N_SCE_c_978_n N_A_27_90#_c_1871_n 0.00337876f $X=3.575 $Y=3.035 $X2=0
+ $Y2=0
cc_794 N_SCE_c_978_n N_A_27_90#_c_1884_n 0.0089164f $X=3.575 $Y=3.035 $X2=0
+ $Y2=0
cc_795 N_SCE_c_980_n N_A_27_90#_c_1884_n 3.74108e-19 $X=3.65 $Y=3.11 $X2=0 $Y2=0
cc_796 N_SCE_c_979_n N_VPWR_c_1994_n 0.00332747f $X=4.56 $Y=3.11 $X2=0 $Y2=0
cc_797 N_SCE_M1003_g N_VPWR_c_1994_n 0.00131924f $X=4.65 $Y=2.63 $X2=0 $Y2=0
cc_798 N_SCE_c_980_n N_VPWR_c_2003_n 0.0269314f $X=3.65 $Y=3.11 $X2=0 $Y2=0
cc_799 N_SCE_c_979_n N_VPWR_c_1991_n 0.0296321f $X=4.56 $Y=3.11 $X2=0 $Y2=0
cc_800 N_SCE_c_980_n N_VPWR_c_1991_n 0.00967894f $X=3.65 $Y=3.11 $X2=0 $Y2=0
cc_801 N_SCE_M1003_g N_A_697_113#_c_2180_n 0.00291272f $X=4.65 $Y=2.63 $X2=0
+ $Y2=0
cc_802 N_SCE_c_979_n N_A_697_113#_c_2182_n 0.0201879f $X=4.56 $Y=3.11 $X2=0
+ $Y2=0
cc_803 N_SCE_M1003_g N_A_697_113#_c_2182_n 0.00724624f $X=4.65 $Y=2.63 $X2=0
+ $Y2=0
cc_804 N_SCE_c_978_n N_A_697_113#_c_2183_n 0.00317889f $X=3.575 $Y=3.035 $X2=0
+ $Y2=0
cc_805 N_SCE_c_979_n N_A_697_113#_c_2183_n 0.00966106f $X=4.56 $Y=3.11 $X2=0
+ $Y2=0
cc_806 N_SCE_M1003_g N_A_697_113#_c_2208_n 0.0129432f $X=4.65 $Y=2.63 $X2=0
+ $Y2=0
cc_807 N_SCE_c_982_n N_A_697_113#_c_2184_n 4.69291e-19 $X=4.65 $Y=2.235 $X2=0
+ $Y2=0
cc_808 N_SCE_M1003_g N_A_697_113#_c_2184_n 0.00717414f $X=4.65 $Y=2.63 $X2=0
+ $Y2=0
cc_809 N_SCE_M1010_g N_A_697_113#_c_2173_n 0.00504831f $X=5.69 $Y=0.835 $X2=0
+ $Y2=0
cc_810 N_SCE_c_978_n N_A_697_113#_c_2178_n 0.00454961f $X=3.575 $Y=3.035 $X2=0
+ $Y2=0
cc_811 N_SCE_c_981_n N_A_697_113#_c_2178_n 2.37385e-19 $X=4.65 $Y=2.145 $X2=0
+ $Y2=0
cc_812 N_SCE_M1010_g N_A_697_113#_c_2179_n 0.00898259f $X=5.69 $Y=0.835 $X2=0
+ $Y2=0
cc_813 N_SCE_M1037_g N_VGND_c_2399_n 0.0129208f $X=4.79 $Y=0.835 $X2=0 $Y2=0
cc_814 N_SCE_c_973_n N_VGND_c_2399_n 0.0241956f $X=5.615 $Y=0.18 $X2=0 $Y2=0
cc_815 N_SCE_M1010_g N_VGND_c_2399_n 0.00881558f $X=5.69 $Y=0.835 $X2=0 $Y2=0
cc_816 N_SCE_c_973_n N_VGND_c_2400_n 0.00974311f $X=5.615 $Y=0.18 $X2=0 $Y2=0
cc_817 N_SCE_M1010_g N_VGND_c_2400_n 4.47958e-19 $X=5.69 $Y=0.835 $X2=0 $Y2=0
cc_818 N_SCE_c_973_n N_VGND_c_2407_n 0.0191126f $X=5.615 $Y=0.18 $X2=0 $Y2=0
cc_819 N_SCE_c_974_n N_VGND_c_2410_n 0.00729608f $X=4.865 $Y=0.18 $X2=0 $Y2=0
cc_820 N_SCE_c_973_n N_VGND_c_2416_n 0.0312755f $X=5.615 $Y=0.18 $X2=0 $Y2=0
cc_821 N_SCE_c_974_n N_VGND_c_2416_n 0.0106181f $X=4.865 $Y=0.18 $X2=0 $Y2=0
cc_822 N_CLK_c_1052_n N_A_1348_368#_M1004_g 0.00303822f $X=6.665 $Y=1.765 $X2=0
+ $Y2=0
cc_823 N_CLK_c_1052_n N_A_1348_368#_c_1324_n 0.00506913f $X=6.665 $Y=1.765 $X2=0
+ $Y2=0
cc_824 N_CLK_c_1053_n N_A_1348_368#_c_1327_n 0.00636314f $X=6.68 $Y=1.22 $X2=0
+ $Y2=0
cc_825 CLK N_A_1348_368#_c_1328_n 0.00116253f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_826 N_CLK_c_1052_n N_A_1348_368#_c_1329_n 9.01767e-19 $X=6.665 $Y=1.765 $X2=0
+ $Y2=0
cc_827 N_CLK_c_1053_n N_A_1348_368#_c_1329_n 0.00218643f $X=6.68 $Y=1.22 $X2=0
+ $Y2=0
cc_828 CLK N_A_1348_368#_c_1329_n 0.0260568f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_829 N_CLK_c_1052_n N_A_1348_368#_c_1330_n 0.00326261f $X=6.665 $Y=1.765 $X2=0
+ $Y2=0
cc_830 N_CLK_c_1053_n N_A_1348_368#_c_1330_n 0.00279126f $X=6.68 $Y=1.22 $X2=0
+ $Y2=0
cc_831 CLK N_A_1348_368#_c_1330_n 0.0213915f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_832 N_CLK_c_1052_n N_A_1348_368#_c_1346_n 0.00542514f $X=6.665 $Y=1.765 $X2=0
+ $Y2=0
cc_833 N_CLK_c_1052_n N_A_1348_368#_c_1347_n 0.00944601f $X=6.665 $Y=1.765 $X2=0
+ $Y2=0
cc_834 CLK N_A_1348_368#_c_1347_n 0.0170562f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_835 N_CLK_c_1052_n N_A_1348_368#_c_1348_n 2.04342e-19 $X=6.665 $Y=1.765 $X2=0
+ $Y2=0
cc_836 CLK N_A_1348_368#_c_1348_n 0.00111517f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_837 N_CLK_c_1052_n N_VPWR_c_1995_n 0.0217138f $X=6.665 $Y=1.765 $X2=0 $Y2=0
cc_838 N_CLK_c_1052_n N_VPWR_c_2005_n 0.00413917f $X=6.665 $Y=1.765 $X2=0 $Y2=0
cc_839 N_CLK_c_1052_n N_VPWR_c_1991_n 0.00421563f $X=6.665 $Y=1.765 $X2=0 $Y2=0
cc_840 N_CLK_c_1052_n N_A_697_113#_c_2173_n 0.0160947f $X=6.665 $Y=1.765 $X2=0
+ $Y2=0
cc_841 N_CLK_c_1053_n N_A_697_113#_c_2173_n 0.00483239f $X=6.68 $Y=1.22 $X2=0
+ $Y2=0
cc_842 CLK N_A_697_113#_c_2173_n 0.0163434f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_843 N_CLK_c_1052_n N_A_697_113#_c_2186_n 0.016211f $X=6.665 $Y=1.765 $X2=0
+ $Y2=0
cc_844 N_CLK_c_1052_n N_A_697_113#_c_2191_n 0.00448856f $X=6.665 $Y=1.765 $X2=0
+ $Y2=0
cc_845 N_CLK_c_1052_n N_A_697_113#_c_2193_n 6.25071e-19 $X=6.665 $Y=1.765 $X2=0
+ $Y2=0
cc_846 N_CLK_c_1053_n N_VGND_c_2400_n 0.00946865f $X=6.68 $Y=1.22 $X2=0 $Y2=0
cc_847 N_CLK_c_1053_n N_VGND_c_2401_n 0.0033335f $X=6.68 $Y=1.22 $X2=0 $Y2=0
cc_848 N_CLK_c_1053_n N_VGND_c_2411_n 0.00434272f $X=6.68 $Y=1.22 $X2=0 $Y2=0
cc_849 N_CLK_c_1053_n N_VGND_c_2416_n 0.00830282f $X=6.68 $Y=1.22 $X2=0 $Y2=0
cc_850 N_A_1549_74#_c_1089_n N_A_1348_368#_M1004_g 0.00162124f $X=7.885 $Y=0.515
+ $X2=0 $Y2=0
cc_851 N_A_1549_74#_c_1091_n N_A_1348_368#_M1004_g 0.00266901f $X=8.05 $Y=0.34
+ $X2=0 $Y2=0
cc_852 N_A_1549_74#_c_1089_n N_A_1348_368#_c_1319_n 0.001217f $X=7.885 $Y=0.515
+ $X2=0 $Y2=0
cc_853 N_A_1549_74#_c_1116_n N_A_1348_368#_c_1333_n 0.00383185f $X=8.585 $Y=1.98
+ $X2=0 $Y2=0
cc_854 N_A_1549_74#_c_1103_n N_A_1348_368#_c_1333_n 2.47642e-19 $X=8.727 $Y=1.82
+ $X2=0 $Y2=0
cc_855 N_A_1549_74#_c_1119_n N_A_1348_368#_c_1333_n 0.00595778f $X=8.75 $Y=2.215
+ $X2=0 $Y2=0
cc_856 N_A_1549_74#_c_1116_n N_A_1348_368#_c_1320_n 0.0119425f $X=8.585 $Y=1.98
+ $X2=0 $Y2=0
cc_857 N_A_1549_74#_c_1089_n N_A_1348_368#_M1042_g 0.00297897f $X=7.885 $Y=0.515
+ $X2=0 $Y2=0
cc_858 N_A_1549_74#_c_1090_n N_A_1348_368#_M1042_g 0.00551157f $X=8.7 $Y=0.34
+ $X2=0 $Y2=0
cc_859 N_A_1549_74#_c_1103_n N_A_1348_368#_M1042_g 0.0303862f $X=8.727 $Y=1.82
+ $X2=0 $Y2=0
cc_860 N_A_1549_74#_c_1106_n N_A_1348_368#_M1042_g 0.0044439f $X=9.485 $Y=1.285
+ $X2=0 $Y2=0
cc_861 N_A_1549_74#_c_1109_n N_A_1348_368#_M1042_g 0.00631727f $X=9.485 $Y=1.12
+ $X2=0 $Y2=0
cc_862 N_A_1549_74#_c_1116_n N_A_1348_368#_c_1335_n 0.00172181f $X=8.585 $Y=1.98
+ $X2=0 $Y2=0
cc_863 N_A_1549_74#_c_1103_n N_A_1348_368#_c_1335_n 0.00656756f $X=8.727 $Y=1.82
+ $X2=0 $Y2=0
cc_864 N_A_1549_74#_c_1119_n N_A_1348_368#_c_1335_n 0.00776904f $X=8.75 $Y=2.215
+ $X2=0 $Y2=0
cc_865 N_A_1549_74#_c_1106_n N_A_1348_368#_c_1335_n 0.0115914f $X=9.485 $Y=1.285
+ $X2=0 $Y2=0
cc_866 N_A_1549_74#_c_1111_n N_A_1348_368#_c_1336_n 0.0134813f $X=9.08 $Y=2.465
+ $X2=0 $Y2=0
cc_867 N_A_1549_74#_c_1119_n N_A_1348_368#_c_1336_n 0.0130968f $X=8.75 $Y=2.215
+ $X2=0 $Y2=0
cc_868 N_A_1549_74#_c_1106_n N_A_1348_368#_c_1336_n 0.00249028f $X=9.485
+ $Y=1.285 $X2=0 $Y2=0
cc_869 N_A_1549_74#_c_1112_n N_A_1348_368#_c_1322_n 0.0124994f $X=13.16 $Y=2.13
+ $X2=0 $Y2=0
cc_870 N_A_1549_74#_c_1114_n N_A_1348_368#_c_1322_n 0.0131679f $X=13.16 $Y=2.465
+ $X2=0 $Y2=0
cc_871 N_A_1549_74#_c_1088_n N_A_1348_368#_c_1322_n 0.0190226f $X=13.16 $Y=2.04
+ $X2=0 $Y2=0
cc_872 N_A_1549_74#_c_1101_n N_A_1348_368#_c_1322_n 3.05307e-19 $X=12.115
+ $Y=1.635 $X2=0 $Y2=0
cc_873 N_A_1549_74#_c_1102_n N_A_1348_368#_c_1322_n 0.00454447f $X=13.065
+ $Y=1.215 $X2=0 $Y2=0
cc_874 N_A_1549_74#_c_1108_n N_A_1348_368#_c_1322_n 0.00535816f $X=13.23 $Y=1.39
+ $X2=0 $Y2=0
cc_875 N_A_1549_74#_c_1110_n N_A_1348_368#_c_1322_n 0.0206403f $X=12.24 $Y=1.635
+ $X2=0 $Y2=0
cc_876 N_A_1549_74#_M1018_g N_A_1348_368#_M1031_g 0.0293233f $X=12.24 $Y=0.69
+ $X2=0 $Y2=0
cc_877 N_A_1549_74#_c_1101_n N_A_1348_368#_M1031_g 8.90301e-19 $X=12.115
+ $Y=1.635 $X2=0 $Y2=0
cc_878 N_A_1549_74#_c_1102_n N_A_1348_368#_M1031_g 0.0115405f $X=13.065 $Y=1.215
+ $X2=0 $Y2=0
cc_879 N_A_1549_74#_c_1107_n N_A_1348_368#_M1031_g 0.00153298f $X=13.23 $Y=1.215
+ $X2=0 $Y2=0
cc_880 N_A_1549_74#_c_1108_n N_A_1348_368#_M1031_g 0.0135859f $X=13.23 $Y=1.39
+ $X2=0 $Y2=0
cc_881 N_A_1549_74#_c_1116_n N_A_1348_368#_c_1326_n 0.00754546f $X=8.585 $Y=1.98
+ $X2=0 $Y2=0
cc_882 N_A_1549_74#_c_1103_n N_A_1348_368#_c_1326_n 0.00841823f $X=8.727 $Y=1.82
+ $X2=0 $Y2=0
cc_883 N_A_1549_74#_c_1119_n N_A_1348_368#_c_1326_n 0.0214945f $X=8.75 $Y=2.215
+ $X2=0 $Y2=0
cc_884 N_A_1549_74#_c_1089_n N_A_1348_368#_c_1330_n 0.00360221f $X=7.885
+ $Y=0.515 $X2=0 $Y2=0
cc_885 N_A_1549_74#_c_1101_n N_A_1348_368#_c_1343_n 0.00361584f $X=12.115
+ $Y=1.635 $X2=0 $Y2=0
cc_886 N_A_1549_74#_c_1110_n N_A_1348_368#_c_1343_n 0.00318012f $X=12.24
+ $Y=1.635 $X2=0 $Y2=0
cc_887 N_A_1549_74#_c_1112_n N_A_1348_368#_c_1345_n 4.05281e-19 $X=13.16 $Y=2.13
+ $X2=0 $Y2=0
cc_888 N_A_1549_74#_c_1088_n N_A_1348_368#_c_1345_n 2.85345e-19 $X=13.16 $Y=2.04
+ $X2=0 $Y2=0
cc_889 N_A_1549_74#_c_1088_n N_A_1348_368#_c_1331_n 0.00112092f $X=13.16 $Y=2.04
+ $X2=0 $Y2=0
cc_890 N_A_1549_74#_c_1101_n N_A_1348_368#_c_1331_n 0.0264923f $X=12.115
+ $Y=1.635 $X2=0 $Y2=0
cc_891 N_A_1549_74#_c_1102_n N_A_1348_368#_c_1331_n 0.0321686f $X=13.065
+ $Y=1.215 $X2=0 $Y2=0
cc_892 N_A_1549_74#_c_1107_n N_A_1348_368#_c_1331_n 0.00480654f $X=13.23
+ $Y=1.215 $X2=0 $Y2=0
cc_893 N_A_1549_74#_c_1108_n N_A_1348_368#_c_1331_n 3.29048e-19 $X=13.23 $Y=1.39
+ $X2=0 $Y2=0
cc_894 N_A_1549_74#_c_1110_n N_A_1348_368#_c_1331_n 0.00217177f $X=12.24
+ $Y=1.635 $X2=0 $Y2=0
cc_895 N_A_1549_74#_c_1095_n N_A_1972_92#_M1035_d 0.00375374f $X=11.24 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_896 N_A_1549_74#_c_1093_n N_A_1972_92#_M1022_g 0.00578009f $X=9.59 $Y=0.85
+ $X2=0 $Y2=0
cc_897 N_A_1549_74#_c_1094_n N_A_1972_92#_M1022_g 0.0134905f $X=10.56 $Y=0.935
+ $X2=0 $Y2=0
cc_898 N_A_1549_74#_c_1184_p N_A_1972_92#_M1022_g 0.00282878f $X=10.645 $Y=0.85
+ $X2=0 $Y2=0
cc_899 N_A_1549_74#_c_1105_n N_A_1972_92#_M1022_g 0.00386455f $X=9.535 $Y=0.935
+ $X2=0 $Y2=0
cc_900 N_A_1549_74#_c_1106_n N_A_1972_92#_M1022_g 0.0211009f $X=9.485 $Y=1.285
+ $X2=0 $Y2=0
cc_901 N_A_1549_74#_c_1109_n N_A_1972_92#_M1022_g 0.0151737f $X=9.485 $Y=1.12
+ $X2=0 $Y2=0
cc_902 N_A_1549_74#_M1018_g N_A_1972_92#_c_1518_n 0.00531899f $X=12.24 $Y=0.69
+ $X2=0 $Y2=0
cc_903 N_A_1549_74#_c_1100_n N_A_1972_92#_c_1518_n 0.00678101f $X=12.102 $Y=1.3
+ $X2=0 $Y2=0
cc_904 N_A_1549_74#_c_1101_n N_A_1972_92#_c_1518_n 0.00263241f $X=12.115
+ $Y=1.635 $X2=0 $Y2=0
cc_905 N_A_1549_74#_c_1110_n N_A_1972_92#_c_1518_n 0.0218104f $X=12.24 $Y=1.635
+ $X2=0 $Y2=0
cc_906 N_A_1549_74#_M1018_g N_A_1972_92#_c_1520_n 0.0605761f $X=12.24 $Y=0.69
+ $X2=0 $Y2=0
cc_907 N_A_1549_74#_c_1095_n N_A_1972_92#_c_1520_n 6.63977e-19 $X=11.24 $Y=0.34
+ $X2=0 $Y2=0
cc_908 N_A_1549_74#_c_1097_n N_A_1972_92#_c_1520_n 0.004173f $X=11.325 $Y=0.85
+ $X2=0 $Y2=0
cc_909 N_A_1549_74#_c_1098_n N_A_1972_92#_c_1520_n 0.0149517f $X=11.95 $Y=0.935
+ $X2=0 $Y2=0
cc_910 N_A_1549_74#_c_1100_n N_A_1972_92#_c_1520_n 0.0052319f $X=12.102 $Y=1.3
+ $X2=0 $Y2=0
cc_911 N_A_1549_74#_c_1094_n N_A_1972_92#_c_1521_n 0.0139439f $X=10.56 $Y=0.935
+ $X2=0 $Y2=0
cc_912 N_A_1549_74#_c_1094_n N_A_1972_92#_c_1522_n 0.0133748f $X=10.56 $Y=0.935
+ $X2=0 $Y2=0
cc_913 N_A_1549_74#_c_1184_p N_A_1972_92#_c_1522_n 0.0178682f $X=10.645 $Y=0.85
+ $X2=0 $Y2=0
cc_914 N_A_1549_74#_c_1095_n N_A_1972_92#_c_1522_n 0.012787f $X=11.24 $Y=0.34
+ $X2=0 $Y2=0
cc_915 N_A_1549_74#_c_1097_n N_A_1972_92#_c_1522_n 0.0188235f $X=11.325 $Y=0.85
+ $X2=0 $Y2=0
cc_916 N_A_1549_74#_c_1099_n N_A_1972_92#_c_1522_n 0.0141449f $X=11.41 $Y=0.935
+ $X2=0 $Y2=0
cc_917 N_A_1549_74#_M1018_g N_A_1972_92#_c_1524_n 2.45325e-19 $X=12.24 $Y=0.69
+ $X2=0 $Y2=0
cc_918 N_A_1549_74#_c_1098_n N_A_1972_92#_c_1524_n 0.024724f $X=11.95 $Y=0.935
+ $X2=0 $Y2=0
cc_919 N_A_1549_74#_c_1099_n N_A_1972_92#_c_1524_n 0.0143351f $X=11.41 $Y=0.935
+ $X2=0 $Y2=0
cc_920 N_A_1549_74#_c_1100_n N_A_1972_92#_c_1524_n 0.00796281f $X=12.102 $Y=1.3
+ $X2=0 $Y2=0
cc_921 N_A_1549_74#_c_1101_n N_A_1972_92#_c_1524_n 0.0153358f $X=12.115 $Y=1.635
+ $X2=0 $Y2=0
cc_922 N_A_1549_74#_c_1095_n N_A_1972_92#_c_1525_n 0.00385216f $X=11.24 $Y=0.34
+ $X2=0 $Y2=0
cc_923 N_A_1549_74#_c_1098_n N_A_1972_92#_c_1525_n 0.0114772f $X=11.95 $Y=0.935
+ $X2=0 $Y2=0
cc_924 N_A_1549_74#_c_1099_n N_A_1972_92#_c_1525_n 0.00455553f $X=11.41 $Y=0.935
+ $X2=0 $Y2=0
cc_925 N_A_1549_74#_c_1094_n N_A_1972_92#_c_1526_n 0.00457354f $X=10.56 $Y=0.935
+ $X2=0 $Y2=0
cc_926 N_A_1549_74#_c_1105_n N_A_1972_92#_c_1526_n 8.37143e-19 $X=9.535 $Y=0.935
+ $X2=0 $Y2=0
cc_927 N_A_1549_74#_c_1094_n N_A_1972_92#_c_1527_n 0.0515812f $X=10.56 $Y=0.935
+ $X2=0 $Y2=0
cc_928 N_A_1549_74#_c_1105_n N_A_1972_92#_c_1527_n 0.0212635f $X=9.535 $Y=0.935
+ $X2=0 $Y2=0
cc_929 N_A_1549_74#_c_1106_n N_A_1972_92#_c_1527_n 2.95568e-19 $X=9.485 $Y=1.285
+ $X2=0 $Y2=0
cc_930 N_A_1549_74#_c_1103_n N_A_1747_118#_M1042_d 0.00410373f $X=8.727 $Y=1.82
+ $X2=-0.19 $Y2=-0.245
cc_931 N_A_1549_74#_c_1094_n N_A_1747_118#_M1035_g 0.00629676f $X=10.56 $Y=0.935
+ $X2=0 $Y2=0
cc_932 N_A_1549_74#_c_1184_p N_A_1747_118#_M1035_g 0.0122913f $X=10.645 $Y=0.85
+ $X2=0 $Y2=0
cc_933 N_A_1549_74#_c_1095_n N_A_1747_118#_M1035_g 0.0103261f $X=11.24 $Y=0.34
+ $X2=0 $Y2=0
cc_934 N_A_1549_74#_c_1096_n N_A_1747_118#_M1035_g 0.00388648f $X=10.73 $Y=0.34
+ $X2=0 $Y2=0
cc_935 N_A_1549_74#_c_1097_n N_A_1747_118#_M1035_g 0.00321589f $X=11.325 $Y=0.85
+ $X2=0 $Y2=0
cc_936 N_A_1549_74#_c_1105_n N_A_1747_118#_c_1625_n 0.0322508f $X=9.535 $Y=0.935
+ $X2=0 $Y2=0
cc_937 N_A_1549_74#_c_1106_n N_A_1747_118#_c_1625_n 0.00356729f $X=9.485
+ $Y=1.285 $X2=0 $Y2=0
cc_938 N_A_1549_74#_c_1109_n N_A_1747_118#_c_1625_n 0.00161427f $X=9.485 $Y=1.12
+ $X2=0 $Y2=0
cc_939 N_A_1549_74#_c_1111_n N_A_1747_118#_c_1630_n 0.00231881f $X=9.08 $Y=2.465
+ $X2=0 $Y2=0
cc_940 N_A_1549_74#_c_1092_n N_A_1747_118#_c_1650_n 0.0172136f $X=9.49 $Y=0.34
+ $X2=0 $Y2=0
cc_941 N_A_1549_74#_c_1103_n N_A_1747_118#_c_1650_n 0.0751122f $X=8.727 $Y=1.82
+ $X2=0 $Y2=0
cc_942 N_A_1549_74#_c_1103_n N_A_1747_118#_c_1626_n 0.0135293f $X=8.727 $Y=1.82
+ $X2=0 $Y2=0
cc_943 N_A_1549_74#_c_1103_n N_A_1747_118#_c_1631_n 0.0428279f $X=8.727 $Y=1.82
+ $X2=0 $Y2=0
cc_944 N_A_1549_74#_c_1119_n N_A_1747_118#_c_1631_n 0.00858092f $X=8.75 $Y=2.215
+ $X2=0 $Y2=0
cc_945 N_A_1549_74#_c_1111_n N_A_1747_118#_c_1632_n 0.00909944f $X=9.08 $Y=2.465
+ $X2=0 $Y2=0
cc_946 N_A_1549_74#_c_1119_n N_A_1747_118#_c_1632_n 0.00527862f $X=8.75 $Y=2.215
+ $X2=0 $Y2=0
cc_947 N_A_1549_74#_c_1094_n N_A_1747_118#_c_1628_n 0.00531123f $X=10.56
+ $Y=0.935 $X2=0 $Y2=0
cc_948 N_A_1549_74#_c_1105_n N_A_1747_118#_c_1628_n 0.0236282f $X=9.535 $Y=0.935
+ $X2=0 $Y2=0
cc_949 N_A_1549_74#_c_1106_n N_A_1747_118#_c_1628_n 0.00218166f $X=9.485
+ $Y=1.285 $X2=0 $Y2=0
cc_950 N_A_1549_74#_M1018_g N_A_2463_74#_c_1800_n 0.00274767f $X=12.24 $Y=0.69
+ $X2=0 $Y2=0
cc_951 N_A_1549_74#_c_1102_n N_A_2463_74#_c_1800_n 0.0224089f $X=13.065 $Y=1.215
+ $X2=0 $Y2=0
cc_952 N_A_1549_74#_M1018_g N_A_2463_74#_c_1721_n 0.00726238f $X=12.24 $Y=0.69
+ $X2=0 $Y2=0
cc_953 N_A_1549_74#_c_1102_n N_A_2463_74#_c_1722_n 0.0298078f $X=13.065 $Y=1.215
+ $X2=0 $Y2=0
cc_954 N_A_1549_74#_c_1107_n N_A_2463_74#_c_1722_n 0.0233024f $X=13.23 $Y=1.215
+ $X2=0 $Y2=0
cc_955 N_A_1549_74#_c_1108_n N_A_2463_74#_c_1722_n 3.0538e-19 $X=13.23 $Y=1.39
+ $X2=0 $Y2=0
cc_956 N_A_1549_74#_c_1112_n N_A_2463_74#_c_1730_n 0.00274086f $X=13.16 $Y=2.13
+ $X2=0 $Y2=0
cc_957 N_A_1549_74#_c_1113_n N_A_2463_74#_c_1730_n 0.00630729f $X=13.16 $Y=2.375
+ $X2=0 $Y2=0
cc_958 N_A_1549_74#_c_1114_n N_A_2463_74#_c_1730_n 0.00529243f $X=13.16 $Y=2.465
+ $X2=0 $Y2=0
cc_959 N_A_1549_74#_c_1088_n N_A_2463_74#_c_1730_n 0.00502906f $X=13.16 $Y=2.04
+ $X2=0 $Y2=0
cc_960 N_A_1549_74#_c_1088_n N_A_2463_74#_c_1731_n 0.00473287f $X=13.16 $Y=2.04
+ $X2=0 $Y2=0
cc_961 N_A_1549_74#_c_1107_n N_A_2463_74#_c_1731_n 0.0143348f $X=13.23 $Y=1.215
+ $X2=0 $Y2=0
cc_962 N_A_1549_74#_c_1108_n N_A_2463_74#_c_1731_n 0.00330283f $X=13.23 $Y=1.39
+ $X2=0 $Y2=0
cc_963 N_A_1549_74#_c_1088_n N_A_2463_74#_c_1732_n 0.00388667f $X=13.16 $Y=2.04
+ $X2=0 $Y2=0
cc_964 N_A_1549_74#_c_1102_n N_A_2463_74#_c_1732_n 0.00181925f $X=13.065
+ $Y=1.215 $X2=0 $Y2=0
cc_965 N_A_1549_74#_c_1107_n N_A_2463_74#_c_1732_n 0.0102143f $X=13.23 $Y=1.215
+ $X2=0 $Y2=0
cc_966 N_A_1549_74#_c_1108_n N_A_2463_74#_c_1732_n 4.28385e-19 $X=13.23 $Y=1.39
+ $X2=0 $Y2=0
cc_967 N_A_1549_74#_c_1107_n N_A_2463_74#_c_1723_n 0.003386f $X=13.23 $Y=1.215
+ $X2=0 $Y2=0
cc_968 N_A_1549_74#_c_1088_n N_A_2463_74#_c_1724_n 7.89853e-19 $X=13.16 $Y=2.04
+ $X2=0 $Y2=0
cc_969 N_A_1549_74#_c_1107_n N_A_2463_74#_c_1724_n 6.62355e-19 $X=13.23 $Y=1.215
+ $X2=0 $Y2=0
cc_970 N_A_1549_74#_c_1114_n N_A_2463_74#_c_1734_n 0.0178544f $X=13.16 $Y=2.465
+ $X2=0 $Y2=0
cc_971 N_A_1549_74#_c_1107_n N_A_2463_74#_c_1725_n 0.0159969f $X=13.23 $Y=1.215
+ $X2=0 $Y2=0
cc_972 N_A_1549_74#_c_1108_n N_A_2463_74#_c_1725_n 9.10574e-19 $X=13.23 $Y=1.39
+ $X2=0 $Y2=0
cc_973 N_A_1549_74#_c_1114_n N_VPWR_c_1999_n 0.00145136f $X=13.16 $Y=2.465 $X2=0
+ $Y2=0
cc_974 N_A_1549_74#_c_1111_n N_VPWR_c_2006_n 0.00444483f $X=9.08 $Y=2.465 $X2=0
+ $Y2=0
cc_975 N_A_1549_74#_c_1114_n N_VPWR_c_2008_n 0.00336933f $X=13.16 $Y=2.465 $X2=0
+ $Y2=0
cc_976 N_A_1549_74#_c_1111_n N_VPWR_c_1991_n 0.00508527f $X=9.08 $Y=2.465 $X2=0
+ $Y2=0
cc_977 N_A_1549_74#_c_1114_n N_VPWR_c_1991_n 0.00543715f $X=13.16 $Y=2.465 $X2=0
+ $Y2=0
cc_978 N_A_1549_74#_c_1116_n N_A_697_113#_c_2187_n 0.0169707f $X=8.585 $Y=1.98
+ $X2=0 $Y2=0
cc_979 N_A_1549_74#_c_1089_n N_A_697_113#_c_2174_n 0.00529576f $X=7.885 $Y=0.515
+ $X2=0 $Y2=0
cc_980 N_A_1549_74#_c_1116_n N_A_697_113#_c_2174_n 0.0311276f $X=8.585 $Y=1.98
+ $X2=0 $Y2=0
cc_981 N_A_1549_74#_c_1103_n N_A_697_113#_c_2174_n 0.0135227f $X=8.727 $Y=1.82
+ $X2=0 $Y2=0
cc_982 N_A_1549_74#_c_1089_n N_A_697_113#_c_2175_n 0.00815189f $X=7.885 $Y=0.515
+ $X2=0 $Y2=0
cc_983 N_A_1549_74#_M1008_d N_A_697_113#_c_2200_n 0.00439762f $X=8.13 $Y=1.84
+ $X2=0 $Y2=0
cc_984 N_A_1549_74#_c_1111_n N_A_697_113#_c_2200_n 3.58206e-19 $X=9.08 $Y=2.465
+ $X2=0 $Y2=0
cc_985 N_A_1549_74#_c_1116_n N_A_697_113#_c_2200_n 0.0166025f $X=8.585 $Y=1.98
+ $X2=0 $Y2=0
cc_986 N_A_1549_74#_c_1119_n N_A_697_113#_c_2200_n 0.00283414f $X=8.75 $Y=2.215
+ $X2=0 $Y2=0
cc_987 N_A_1549_74#_M1008_d N_A_697_113#_c_2265_n 0.00519937f $X=8.13 $Y=1.84
+ $X2=0 $Y2=0
cc_988 N_A_1549_74#_c_1111_n N_A_697_113#_c_2265_n 0.00398193f $X=9.08 $Y=2.465
+ $X2=0 $Y2=0
cc_989 N_A_1549_74#_c_1089_n N_A_697_113#_c_2176_n 0.0345841f $X=7.885 $Y=0.515
+ $X2=0 $Y2=0
cc_990 N_A_1549_74#_c_1090_n N_A_697_113#_c_2176_n 0.0191962f $X=8.7 $Y=0.34
+ $X2=0 $Y2=0
cc_991 N_A_1549_74#_c_1103_n N_A_697_113#_c_2176_n 0.0486628f $X=8.727 $Y=1.82
+ $X2=0 $Y2=0
cc_992 N_A_1549_74#_M1008_d N_A_697_113#_c_2188_n 0.00188412f $X=8.13 $Y=1.84
+ $X2=0 $Y2=0
cc_993 N_A_1549_74#_M1008_d N_A_697_113#_c_2189_n 0.00290816f $X=8.13 $Y=1.84
+ $X2=0 $Y2=0
cc_994 N_A_1549_74#_c_1111_n N_A_697_113#_c_2189_n 0.0035695f $X=9.08 $Y=2.465
+ $X2=0 $Y2=0
cc_995 N_A_1549_74#_c_1116_n N_A_697_113#_c_2189_n 0.0214293f $X=8.585 $Y=1.98
+ $X2=0 $Y2=0
cc_996 N_A_1549_74#_c_1119_n N_A_697_113#_c_2189_n 0.00483701f $X=8.75 $Y=2.215
+ $X2=0 $Y2=0
cc_997 N_A_1549_74#_c_1094_n N_VGND_M1022_d 0.00955404f $X=10.56 $Y=0.935 $X2=0
+ $Y2=0
cc_998 N_A_1549_74#_c_1184_p N_VGND_M1022_d 0.00519548f $X=10.645 $Y=0.85 $X2=0
+ $Y2=0
cc_999 N_A_1549_74#_c_1096_n N_VGND_M1022_d 6.10141e-19 $X=10.73 $Y=0.34 $X2=0
+ $Y2=0
cc_1000 N_A_1549_74#_c_1098_n N_VGND_M1016_s 0.00391333f $X=11.95 $Y=0.935 $X2=0
+ $Y2=0
cc_1001 N_A_1549_74#_c_1091_n N_VGND_c_2401_n 0.0112234f $X=8.05 $Y=0.34 $X2=0
+ $Y2=0
cc_1002 N_A_1549_74#_c_1092_n N_VGND_c_2402_n 0.00867558f $X=9.49 $Y=0.34 $X2=0
+ $Y2=0
cc_1003 N_A_1549_74#_c_1093_n N_VGND_c_2402_n 0.00945189f $X=9.59 $Y=0.85 $X2=0
+ $Y2=0
cc_1004 N_A_1549_74#_c_1094_n N_VGND_c_2402_n 0.025645f $X=10.56 $Y=0.935 $X2=0
+ $Y2=0
cc_1005 N_A_1549_74#_c_1184_p N_VGND_c_2402_n 0.0194279f $X=10.645 $Y=0.85 $X2=0
+ $Y2=0
cc_1006 N_A_1549_74#_c_1096_n N_VGND_c_2402_n 0.0148401f $X=10.73 $Y=0.34 $X2=0
+ $Y2=0
cc_1007 N_A_1549_74#_M1018_g N_VGND_c_2403_n 0.00147043f $X=12.24 $Y=0.69 $X2=0
+ $Y2=0
cc_1008 N_A_1549_74#_c_1095_n N_VGND_c_2403_n 0.0146661f $X=11.24 $Y=0.34 $X2=0
+ $Y2=0
cc_1009 N_A_1549_74#_c_1097_n N_VGND_c_2403_n 0.0193741f $X=11.325 $Y=0.85 $X2=0
+ $Y2=0
cc_1010 N_A_1549_74#_c_1098_n N_VGND_c_2403_n 0.015048f $X=11.95 $Y=0.935 $X2=0
+ $Y2=0
cc_1011 N_A_1549_74#_c_1090_n N_VGND_c_2412_n 0.0418136f $X=8.7 $Y=0.34 $X2=0
+ $Y2=0
cc_1012 N_A_1549_74#_c_1091_n N_VGND_c_2412_n 0.0179217f $X=8.05 $Y=0.34 $X2=0
+ $Y2=0
cc_1013 N_A_1549_74#_c_1092_n N_VGND_c_2412_n 0.0542184f $X=9.49 $Y=0.34 $X2=0
+ $Y2=0
cc_1014 N_A_1549_74#_c_1104_n N_VGND_c_2412_n 0.0121867f $X=8.785 $Y=0.34 $X2=0
+ $Y2=0
cc_1015 N_A_1549_74#_c_1095_n N_VGND_c_2413_n 0.0446936f $X=11.24 $Y=0.34 $X2=0
+ $Y2=0
cc_1016 N_A_1549_74#_c_1096_n N_VGND_c_2413_n 0.012011f $X=10.73 $Y=0.34 $X2=0
+ $Y2=0
cc_1017 N_A_1549_74#_M1018_g N_VGND_c_2416_n 0.00821463f $X=12.24 $Y=0.69 $X2=0
+ $Y2=0
cc_1018 N_A_1549_74#_c_1090_n N_VGND_c_2416_n 0.0244305f $X=8.7 $Y=0.34 $X2=0
+ $Y2=0
cc_1019 N_A_1549_74#_c_1091_n N_VGND_c_2416_n 0.00971942f $X=8.05 $Y=0.34 $X2=0
+ $Y2=0
cc_1020 N_A_1549_74#_c_1092_n N_VGND_c_2416_n 0.0310781f $X=9.49 $Y=0.34 $X2=0
+ $Y2=0
cc_1021 N_A_1549_74#_c_1094_n N_VGND_c_2416_n 0.0192226f $X=10.56 $Y=0.935 $X2=0
+ $Y2=0
cc_1022 N_A_1549_74#_c_1095_n N_VGND_c_2416_n 0.0253215f $X=11.24 $Y=0.34 $X2=0
+ $Y2=0
cc_1023 N_A_1549_74#_c_1096_n N_VGND_c_2416_n 0.00638043f $X=10.73 $Y=0.34 $X2=0
+ $Y2=0
cc_1024 N_A_1549_74#_c_1098_n N_VGND_c_2416_n 0.00988673f $X=11.95 $Y=0.935
+ $X2=0 $Y2=0
cc_1025 N_A_1549_74#_c_1100_n N_VGND_c_2416_n 0.00660638f $X=12.102 $Y=1.3 $X2=0
+ $Y2=0
cc_1026 N_A_1549_74#_c_1104_n N_VGND_c_2416_n 0.00660921f $X=8.785 $Y=0.34 $X2=0
+ $Y2=0
cc_1027 N_A_1549_74#_M1018_g N_VGND_c_2422_n 0.00434272f $X=12.24 $Y=0.69 $X2=0
+ $Y2=0
cc_1028 N_A_1549_74#_c_1093_n A_1895_118# 0.00521187f $X=9.59 $Y=0.85 $X2=-0.19
+ $Y2=-0.245
cc_1029 N_A_1549_74#_c_1094_n A_1895_118# 0.00227085f $X=10.56 $Y=0.935
+ $X2=-0.19 $Y2=-0.245
cc_1030 N_A_1549_74#_c_1105_n A_1895_118# 7.37266e-19 $X=9.535 $Y=0.935
+ $X2=-0.19 $Y2=-0.245
cc_1031 N_A_1549_74#_c_1100_n A_2391_74# 0.00229931f $X=12.102 $Y=1.3 $X2=-0.19
+ $Y2=-0.245
cc_1032 N_A_1348_368#_c_1343_n N_A_1972_92#_M1005_d 0.00779702f $X=12.425
+ $Y=2.475 $X2=0 $Y2=0
cc_1033 N_A_1348_368#_c_1336_n N_A_1972_92#_c_1517_n 0.0385867f $X=9.58 $Y=2.465
+ $X2=0 $Y2=0
cc_1034 N_A_1348_368#_c_1341_n N_A_1972_92#_c_1517_n 0.00643117f $X=9.69 $Y=2.09
+ $X2=0 $Y2=0
cc_1035 N_A_1348_368#_c_1342_n N_A_1972_92#_c_1517_n 0.00392779f $X=9.775
+ $Y=2.39 $X2=0 $Y2=0
cc_1036 N_A_1348_368#_c_1336_n N_A_1972_92#_c_1530_n 0.0267627f $X=9.58 $Y=2.465
+ $X2=0 $Y2=0
cc_1037 N_A_1348_368#_c_1343_n N_A_1972_92#_c_1530_n 0.0147368f $X=12.425
+ $Y=2.475 $X2=0 $Y2=0
cc_1038 N_A_1348_368#_c_1343_n N_A_1972_92#_c_1532_n 0.0163341f $X=12.425
+ $Y=2.475 $X2=0 $Y2=0
cc_1039 N_A_1348_368#_c_1345_n N_A_1972_92#_c_1532_n 0.0017491f $X=12.51 $Y=2.39
+ $X2=0 $Y2=0
cc_1040 N_A_1348_368#_c_1343_n N_A_1972_92#_c_1533_n 0.0285202f $X=12.425
+ $Y=2.475 $X2=0 $Y2=0
cc_1041 N_A_1348_368#_c_1343_n N_A_1747_118#_c_1623_n 0.0165356f $X=12.425
+ $Y=2.475 $X2=0 $Y2=0
cc_1042 N_A_1348_368#_c_1326_n N_A_1747_118#_c_1625_n 0.0016426f $X=8.66
+ $Y=1.727 $X2=0 $Y2=0
cc_1043 N_A_1348_368#_c_1336_n N_A_1747_118#_c_1630_n 0.00782963f $X=9.58
+ $Y=2.465 $X2=0 $Y2=0
cc_1044 N_A_1348_368#_M1042_g N_A_1747_118#_c_1650_n 0.0016426f $X=8.66 $Y=0.8
+ $X2=0 $Y2=0
cc_1045 N_A_1348_368#_c_1335_n N_A_1747_118#_c_1626_n 0.00714571f $X=9.38
+ $Y=1.765 $X2=0 $Y2=0
cc_1046 N_A_1348_368#_c_1326_n N_A_1747_118#_c_1626_n 3.95135e-19 $X=8.66
+ $Y=1.727 $X2=0 $Y2=0
cc_1047 N_A_1348_368#_c_1335_n N_A_1747_118#_c_1631_n 0.00629732f $X=9.38
+ $Y=1.765 $X2=0 $Y2=0
cc_1048 N_A_1348_368#_c_1336_n N_A_1747_118#_c_1631_n 0.00682785f $X=9.58
+ $Y=2.465 $X2=0 $Y2=0
cc_1049 N_A_1348_368#_c_1341_n N_A_1747_118#_c_1631_n 0.0187531f $X=9.69 $Y=2.09
+ $X2=0 $Y2=0
cc_1050 N_A_1348_368#_c_1342_n N_A_1747_118#_c_1631_n 0.00602345f $X=9.775
+ $Y=2.39 $X2=0 $Y2=0
cc_1051 N_A_1348_368#_c_1335_n N_A_1747_118#_c_1632_n 0.00269406f $X=9.38
+ $Y=1.765 $X2=0 $Y2=0
cc_1052 N_A_1348_368#_c_1336_n N_A_1747_118#_c_1632_n 0.00764087f $X=9.58
+ $Y=2.465 $X2=0 $Y2=0
cc_1053 N_A_1348_368#_c_1341_n N_A_1747_118#_c_1632_n 0.0103858f $X=9.69 $Y=2.09
+ $X2=0 $Y2=0
cc_1054 N_A_1348_368#_c_1344_n N_A_1747_118#_c_1632_n 0.0136934f $X=9.86
+ $Y=2.475 $X2=0 $Y2=0
cc_1055 N_A_1348_368#_c_1343_n N_A_1747_118#_c_1627_n 0.00207969f $X=12.425
+ $Y=2.475 $X2=0 $Y2=0
cc_1056 N_A_1348_368#_c_1335_n N_A_1747_118#_c_1628_n 0.00602187f $X=9.38
+ $Y=1.765 $X2=0 $Y2=0
cc_1057 N_A_1348_368#_c_1336_n N_A_1747_118#_c_1628_n 0.00824036f $X=9.58
+ $Y=2.465 $X2=0 $Y2=0
cc_1058 N_A_1348_368#_c_1341_n N_A_1747_118#_c_1628_n 0.0331302f $X=9.69 $Y=2.09
+ $X2=0 $Y2=0
cc_1059 N_A_1348_368#_c_1343_n N_A_1747_118#_c_1628_n 0.0061485f $X=12.425
+ $Y=2.475 $X2=0 $Y2=0
cc_1060 N_A_1348_368#_M1031_g N_A_2463_74#_c_1721_n 0.00236994f $X=12.75 $Y=0.58
+ $X2=0 $Y2=0
cc_1061 N_A_1348_368#_M1031_g N_A_2463_74#_c_1722_n 0.0118688f $X=12.75 $Y=0.58
+ $X2=0 $Y2=0
cc_1062 N_A_1348_368#_c_1322_n N_A_2463_74#_c_1730_n 0.00416226f $X=12.625
+ $Y=1.885 $X2=0 $Y2=0
cc_1063 N_A_1348_368#_c_1343_n N_A_2463_74#_c_1730_n 0.0051562f $X=12.425
+ $Y=2.475 $X2=0 $Y2=0
cc_1064 N_A_1348_368#_c_1345_n N_A_2463_74#_c_1730_n 0.0163192f $X=12.51 $Y=2.39
+ $X2=0 $Y2=0
cc_1065 N_A_1348_368#_c_1322_n N_A_2463_74#_c_1732_n 0.0010855f $X=12.625
+ $Y=1.885 $X2=0 $Y2=0
cc_1066 N_A_1348_368#_c_1345_n N_A_2463_74#_c_1732_n 0.00344187f $X=12.51
+ $Y=2.39 $X2=0 $Y2=0
cc_1067 N_A_1348_368#_c_1331_n N_A_2463_74#_c_1732_n 0.00724947f $X=12.69
+ $Y=1.635 $X2=0 $Y2=0
cc_1068 N_A_1348_368#_c_1322_n N_A_2463_74#_c_1734_n 0.010605f $X=12.625
+ $Y=1.885 $X2=0 $Y2=0
cc_1069 N_A_1348_368#_c_1343_n N_A_2463_74#_c_1734_n 0.00329319f $X=12.425
+ $Y=2.475 $X2=0 $Y2=0
cc_1070 N_A_1348_368#_c_1343_n N_VPWR_M1041_d 0.00677866f $X=12.425 $Y=2.475
+ $X2=0 $Y2=0
cc_1071 N_A_1348_368#_c_1343_n N_VPWR_M1038_s 0.0100777f $X=12.425 $Y=2.475
+ $X2=0 $Y2=0
cc_1072 N_A_1348_368#_c_1333_n N_VPWR_c_1996_n 0.0109611f $X=8.055 $Y=1.765
+ $X2=0 $Y2=0
cc_1073 N_A_1348_368#_c_1336_n N_VPWR_c_1997_n 0.00124671f $X=9.58 $Y=2.465
+ $X2=0 $Y2=0
cc_1074 N_A_1348_368#_c_1343_n N_VPWR_c_1997_n 0.0213705f $X=12.425 $Y=2.475
+ $X2=0 $Y2=0
cc_1075 N_A_1348_368#_c_1343_n N_VPWR_c_1998_n 0.0259982f $X=12.425 $Y=2.475
+ $X2=0 $Y2=0
cc_1076 N_A_1348_368#_c_1333_n N_VPWR_c_2006_n 0.00413917f $X=8.055 $Y=1.765
+ $X2=0 $Y2=0
cc_1077 N_A_1348_368#_c_1336_n N_VPWR_c_2006_n 0.00445602f $X=9.58 $Y=2.465
+ $X2=0 $Y2=0
cc_1078 N_A_1348_368#_c_1322_n N_VPWR_c_2008_n 0.00461464f $X=12.625 $Y=1.885
+ $X2=0 $Y2=0
cc_1079 N_A_1348_368#_c_1333_n N_VPWR_c_1991_n 0.00421563f $X=8.055 $Y=1.765
+ $X2=0 $Y2=0
cc_1080 N_A_1348_368#_c_1336_n N_VPWR_c_1991_n 0.0089489f $X=9.58 $Y=2.465 $X2=0
+ $Y2=0
cc_1081 N_A_1348_368#_c_1322_n N_VPWR_c_1991_n 0.00776565f $X=12.625 $Y=1.885
+ $X2=0 $Y2=0
cc_1082 N_A_1348_368#_c_1343_n N_VPWR_c_1991_n 0.0765599f $X=12.425 $Y=2.475
+ $X2=0 $Y2=0
cc_1083 N_A_1348_368#_c_1344_n N_VPWR_c_1991_n 0.00704359f $X=9.86 $Y=2.475
+ $X2=0 $Y2=0
cc_1084 N_A_1348_368#_c_1347_n N_A_697_113#_c_2173_n 0.00867645f $X=7.055
+ $Y=1.975 $X2=0 $Y2=0
cc_1085 N_A_1348_368#_M1034_d N_A_697_113#_c_2186_n 0.00821192f $X=6.74 $Y=1.84
+ $X2=0 $Y2=0
cc_1086 N_A_1348_368#_c_1324_n N_A_697_113#_c_2186_n 0.00446176f $X=7.47 $Y=1.69
+ $X2=0 $Y2=0
cc_1087 N_A_1348_368#_c_1346_n N_A_697_113#_c_2186_n 0.00814455f $X=7.36
+ $Y=1.975 $X2=0 $Y2=0
cc_1088 N_A_1348_368#_c_1347_n N_A_697_113#_c_2186_n 0.0517307f $X=7.055
+ $Y=1.975 $X2=0 $Y2=0
cc_1089 N_A_1348_368#_c_1319_n N_A_697_113#_c_2187_n 0.0114826f $X=7.98 $Y=1.69
+ $X2=0 $Y2=0
cc_1090 N_A_1348_368#_c_1333_n N_A_697_113#_c_2187_n 0.00702413f $X=8.055
+ $Y=1.765 $X2=0 $Y2=0
cc_1091 N_A_1348_368#_c_1330_n N_A_697_113#_c_2187_n 0.00809291f $X=7.44 $Y=1.81
+ $X2=0 $Y2=0
cc_1092 N_A_1348_368#_c_1346_n N_A_697_113#_c_2187_n 0.00150572f $X=7.36
+ $Y=1.975 $X2=0 $Y2=0
cc_1093 N_A_1348_368#_c_1348_n N_A_697_113#_c_2187_n 0.017236f $X=7.44 $Y=1.975
+ $X2=0 $Y2=0
cc_1094 N_A_1348_368#_c_1319_n N_A_697_113#_c_2174_n 0.00152648f $X=7.98 $Y=1.69
+ $X2=0 $Y2=0
cc_1095 N_A_1348_368#_c_1320_n N_A_697_113#_c_2174_n 0.0127033f $X=8.585 $Y=1.69
+ $X2=0 $Y2=0
cc_1096 N_A_1348_368#_M1042_g N_A_697_113#_c_2174_n 0.00309069f $X=8.66 $Y=0.8
+ $X2=0 $Y2=0
cc_1097 N_A_1348_368#_c_1325_n N_A_697_113#_c_2174_n 0.00674941f $X=8.055
+ $Y=1.69 $X2=0 $Y2=0
cc_1098 N_A_1348_368#_M1004_g N_A_697_113#_c_2175_n 0.00342028f $X=7.67 $Y=0.74
+ $X2=0 $Y2=0
cc_1099 N_A_1348_368#_c_1319_n N_A_697_113#_c_2175_n 0.00305869f $X=7.98 $Y=1.69
+ $X2=0 $Y2=0
cc_1100 N_A_1348_368#_c_1330_n N_A_697_113#_c_2175_n 0.0106446f $X=7.44 $Y=1.81
+ $X2=0 $Y2=0
cc_1101 N_A_1348_368#_c_1333_n N_A_697_113#_c_2200_n 0.0160314f $X=8.055
+ $Y=1.765 $X2=0 $Y2=0
cc_1102 N_A_1348_368#_M1004_g N_A_697_113#_c_2176_n 0.0094266f $X=7.67 $Y=0.74
+ $X2=0 $Y2=0
cc_1103 N_A_1348_368#_M1042_g N_A_697_113#_c_2176_n 0.0109029f $X=8.66 $Y=0.8
+ $X2=0 $Y2=0
cc_1104 N_A_1348_368#_c_1333_n N_A_697_113#_c_2188_n 0.00497744f $X=8.055
+ $Y=1.765 $X2=0 $Y2=0
cc_1105 N_A_1348_368#_c_1343_n A_1931_508# 3.21084e-19 $X=12.425 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_1106 N_A_1348_368#_c_1344_n A_1931_508# 0.00328363f $X=9.86 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_1107 N_A_1348_368#_c_1343_n A_2345_392# 0.0269035f $X=12.425 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_1108 N_A_1348_368#_c_1345_n A_2345_392# 0.0134123f $X=12.51 $Y=2.39 $X2=-0.19
+ $Y2=-0.245
cc_1109 N_A_1348_368#_c_1328_n N_VGND_M1004_s 0.00675916f $X=7.355 $Y=0.925
+ $X2=0 $Y2=0
cc_1110 N_A_1348_368#_c_1330_n N_VGND_M1004_s 0.00355875f $X=7.44 $Y=1.81 $X2=0
+ $Y2=0
cc_1111 N_A_1348_368#_c_1327_n N_VGND_c_2400_n 0.018213f $X=6.895 $Y=0.515 $X2=0
+ $Y2=0
cc_1112 N_A_1348_368#_M1004_g N_VGND_c_2401_n 0.00936698f $X=7.67 $Y=0.74 $X2=0
+ $Y2=0
cc_1113 N_A_1348_368#_c_1327_n N_VGND_c_2401_n 0.0215739f $X=6.895 $Y=0.515
+ $X2=0 $Y2=0
cc_1114 N_A_1348_368#_c_1328_n N_VGND_c_2401_n 0.020074f $X=7.355 $Y=0.925 $X2=0
+ $Y2=0
cc_1115 N_A_1348_368#_c_1327_n N_VGND_c_2411_n 0.0145323f $X=6.895 $Y=0.515
+ $X2=0 $Y2=0
cc_1116 N_A_1348_368#_M1004_g N_VGND_c_2412_n 0.00383152f $X=7.67 $Y=0.74 $X2=0
+ $Y2=0
cc_1117 N_A_1348_368#_M1042_g N_VGND_c_2412_n 2.67369e-19 $X=8.66 $Y=0.8 $X2=0
+ $Y2=0
cc_1118 N_A_1348_368#_M1004_g N_VGND_c_2416_n 0.00762539f $X=7.67 $Y=0.74 $X2=0
+ $Y2=0
cc_1119 N_A_1348_368#_M1031_g N_VGND_c_2416_n 0.00447595f $X=12.75 $Y=0.58 $X2=0
+ $Y2=0
cc_1120 N_A_1348_368#_c_1327_n N_VGND_c_2416_n 0.0119861f $X=6.895 $Y=0.515
+ $X2=0 $Y2=0
cc_1121 N_A_1348_368#_c_1328_n N_VGND_c_2416_n 0.00878953f $X=7.355 $Y=0.925
+ $X2=0 $Y2=0
cc_1122 N_A_1348_368#_M1031_g N_VGND_c_2422_n 0.00461464f $X=12.75 $Y=0.58 $X2=0
+ $Y2=0
cc_1123 N_A_1348_368#_M1031_g N_VGND_c_2423_n 0.00128745f $X=12.75 $Y=0.58 $X2=0
+ $Y2=0
cc_1124 N_A_1972_92#_c_1517_n N_A_1747_118#_c_1623_n 0.0356437f $X=10.01
+ $Y=2.375 $X2=0 $Y2=0
cc_1125 N_A_1972_92#_c_1530_n N_A_1747_118#_c_1623_n 0.00936349f $X=10.01
+ $Y=2.465 $X2=0 $Y2=0
cc_1126 N_A_1972_92#_c_1521_n N_A_1747_118#_c_1623_n 0.00714712f $X=10.9
+ $Y=1.275 $X2=0 $Y2=0
cc_1127 N_A_1972_92#_c_1533_n N_A_1747_118#_c_1623_n 0.00953376f $X=10.9
+ $Y=2.135 $X2=0 $Y2=0
cc_1128 N_A_1972_92#_c_1523_n N_A_1747_118#_c_1623_n 0.0139157f $X=10.985
+ $Y=2.05 $X2=0 $Y2=0
cc_1129 N_A_1972_92#_M1022_g N_A_1747_118#_M1035_g 0.00896516f $X=9.935 $Y=0.8
+ $X2=0 $Y2=0
cc_1130 N_A_1972_92#_c_1517_n N_A_1747_118#_M1035_g 3.69694e-19 $X=10.01
+ $Y=2.375 $X2=0 $Y2=0
cc_1131 N_A_1972_92#_c_1521_n N_A_1747_118#_M1035_g 0.0150675f $X=10.9 $Y=1.275
+ $X2=0 $Y2=0
cc_1132 N_A_1972_92#_c_1522_n N_A_1747_118#_M1035_g 0.00704904f $X=10.985
+ $Y=0.81 $X2=0 $Y2=0
cc_1133 N_A_1972_92#_c_1525_n N_A_1747_118#_M1035_g 0.0212503f $X=11.575
+ $Y=1.355 $X2=0 $Y2=0
cc_1134 N_A_1972_92#_c_1526_n N_A_1747_118#_M1035_g 0.00747304f $X=10.025
+ $Y=1.32 $X2=0 $Y2=0
cc_1135 N_A_1972_92#_c_1527_n N_A_1747_118#_M1035_g 4.80678e-19 $X=10.19 $Y=1.32
+ $X2=0 $Y2=0
cc_1136 N_A_1972_92#_c_1528_n N_A_1747_118#_M1035_g 0.00490245f $X=10.985
+ $Y=1.355 $X2=0 $Y2=0
cc_1137 N_A_1972_92#_c_1526_n N_A_1747_118#_c_1625_n 8.02253e-19 $X=10.025
+ $Y=1.32 $X2=0 $Y2=0
cc_1138 N_A_1972_92#_c_1530_n N_A_1747_118#_c_1632_n 0.00166172f $X=10.01
+ $Y=2.465 $X2=0 $Y2=0
cc_1139 N_A_1972_92#_c_1517_n N_A_1747_118#_c_1627_n 8.06641e-19 $X=10.01
+ $Y=2.375 $X2=0 $Y2=0
cc_1140 N_A_1972_92#_c_1521_n N_A_1747_118#_c_1627_n 0.0238486f $X=10.9 $Y=1.275
+ $X2=0 $Y2=0
cc_1141 N_A_1972_92#_c_1533_n N_A_1747_118#_c_1627_n 0.00475756f $X=10.9
+ $Y=2.135 $X2=0 $Y2=0
cc_1142 N_A_1972_92#_c_1523_n N_A_1747_118#_c_1627_n 0.0232504f $X=10.985
+ $Y=2.05 $X2=0 $Y2=0
cc_1143 N_A_1972_92#_c_1517_n N_A_1747_118#_c_1628_n 0.0149344f $X=10.01
+ $Y=2.375 $X2=0 $Y2=0
cc_1144 N_A_1972_92#_c_1521_n N_A_1747_118#_c_1628_n 0.0109136f $X=10.9 $Y=1.275
+ $X2=0 $Y2=0
cc_1145 N_A_1972_92#_c_1526_n N_A_1747_118#_c_1628_n 0.0037499f $X=10.025
+ $Y=1.32 $X2=0 $Y2=0
cc_1146 N_A_1972_92#_c_1527_n N_A_1747_118#_c_1628_n 0.0228829f $X=10.19 $Y=1.32
+ $X2=0 $Y2=0
cc_1147 N_A_1972_92#_c_1520_n N_A_2463_74#_c_1800_n 4.65641e-19 $X=11.88 $Y=1.11
+ $X2=0 $Y2=0
cc_1148 N_A_1972_92#_c_1520_n N_A_2463_74#_c_1721_n 0.00134647f $X=11.88 $Y=1.11
+ $X2=0 $Y2=0
cc_1149 N_A_1972_92#_c_1530_n N_VPWR_c_1997_n 0.0086591f $X=10.01 $Y=2.465 $X2=0
+ $Y2=0
cc_1150 N_A_1972_92#_c_1532_n N_VPWR_c_1998_n 0.0148532f $X=11.65 $Y=1.885 $X2=0
+ $Y2=0
cc_1151 N_A_1972_92#_c_1530_n N_VPWR_c_2006_n 0.00444681f $X=10.01 $Y=2.465
+ $X2=0 $Y2=0
cc_1152 N_A_1972_92#_c_1532_n N_VPWR_c_2008_n 0.00461464f $X=11.65 $Y=1.885
+ $X2=0 $Y2=0
cc_1153 N_A_1972_92#_c_1530_n N_VPWR_c_1991_n 0.00427716f $X=10.01 $Y=2.465
+ $X2=0 $Y2=0
cc_1154 N_A_1972_92#_c_1532_n N_VPWR_c_1991_n 0.0045644f $X=11.65 $Y=1.885 $X2=0
+ $Y2=0
cc_1155 N_A_1972_92#_M1022_g N_VGND_c_2402_n 0.00272252f $X=9.935 $Y=0.8 $X2=0
+ $Y2=0
cc_1156 N_A_1972_92#_c_1520_n N_VGND_c_2403_n 0.010393f $X=11.88 $Y=1.11 $X2=0
+ $Y2=0
cc_1157 N_A_1972_92#_M1022_g N_VGND_c_2412_n 0.00434252f $X=9.935 $Y=0.8 $X2=0
+ $Y2=0
cc_1158 N_A_1972_92#_M1022_g N_VGND_c_2416_n 0.00479212f $X=9.935 $Y=0.8 $X2=0
+ $Y2=0
cc_1159 N_A_1972_92#_c_1520_n N_VGND_c_2416_n 0.0038545f $X=11.88 $Y=1.11 $X2=0
+ $Y2=0
cc_1160 N_A_1972_92#_c_1520_n N_VGND_c_2422_n 0.00383152f $X=11.88 $Y=1.11 $X2=0
+ $Y2=0
cc_1161 N_A_1747_118#_c_1623_n N_VPWR_c_1997_n 0.00644269f $X=10.555 $Y=1.915
+ $X2=0 $Y2=0
cc_1162 N_A_1747_118#_c_1630_n N_VPWR_c_1997_n 0.00703659f $X=9.355 $Y=2.75
+ $X2=0 $Y2=0
cc_1163 N_A_1747_118#_c_1623_n N_VPWR_c_1998_n 0.0057683f $X=10.555 $Y=1.915
+ $X2=0 $Y2=0
cc_1164 N_A_1747_118#_c_1630_n N_VPWR_c_2006_n 0.014453f $X=9.355 $Y=2.75 $X2=0
+ $Y2=0
cc_1165 N_A_1747_118#_c_1623_n N_VPWR_c_2007_n 0.00487664f $X=10.555 $Y=1.915
+ $X2=0 $Y2=0
cc_1166 N_A_1747_118#_c_1623_n N_VPWR_c_1991_n 0.00505379f $X=10.555 $Y=1.915
+ $X2=0 $Y2=0
cc_1167 N_A_1747_118#_c_1630_n N_VPWR_c_1991_n 0.011992f $X=9.355 $Y=2.75 $X2=0
+ $Y2=0
cc_1168 N_A_1747_118#_c_1632_n N_VPWR_c_1991_n 0.00536095f $X=9.28 $Y=2.56 $X2=0
+ $Y2=0
cc_1169 N_A_1747_118#_c_1630_n N_A_697_113#_c_2189_n 0.0111988f $X=9.355 $Y=2.75
+ $X2=0 $Y2=0
cc_1170 N_A_1747_118#_M1035_g N_VGND_c_2402_n 0.0023268f $X=10.755 $Y=0.69 $X2=0
+ $Y2=0
cc_1171 N_A_1747_118#_M1035_g N_VGND_c_2413_n 0.00278223f $X=10.755 $Y=0.69
+ $X2=0 $Y2=0
cc_1172 N_A_1747_118#_M1035_g N_VGND_c_2416_n 0.00363422f $X=10.755 $Y=0.69
+ $X2=0 $Y2=0
cc_1173 N_A_2463_74#_c_1727_n N_VPWR_c_1999_n 0.0172212f $X=14.29 $Y=1.885 $X2=0
+ $Y2=0
cc_1174 N_A_2463_74#_c_1734_n N_VPWR_c_1999_n 0.0121119f $X=13.11 $Y=2.75 $X2=0
+ $Y2=0
cc_1175 N_A_2463_74#_c_1729_n N_VPWR_c_2000_n 0.00731351f $X=15.3 $Y=1.765 $X2=0
+ $Y2=0
cc_1176 N_A_2463_74#_c_1734_n N_VPWR_c_2008_n 0.018246f $X=13.11 $Y=2.75 $X2=0
+ $Y2=0
cc_1177 N_A_2463_74#_c_1727_n N_VPWR_c_2009_n 0.00413917f $X=14.29 $Y=1.885
+ $X2=0 $Y2=0
cc_1178 N_A_2463_74#_c_1729_n N_VPWR_c_2009_n 0.00445602f $X=15.3 $Y=1.765 $X2=0
+ $Y2=0
cc_1179 N_A_2463_74#_c_1727_n N_VPWR_c_1991_n 0.00822528f $X=14.29 $Y=1.885
+ $X2=0 $Y2=0
cc_1180 N_A_2463_74#_c_1729_n N_VPWR_c_1991_n 0.00862905f $X=15.3 $Y=1.765 $X2=0
+ $Y2=0
cc_1181 N_A_2463_74#_c_1734_n N_VPWR_c_1991_n 0.0151301f $X=13.11 $Y=2.75 $X2=0
+ $Y2=0
cc_1182 N_A_2463_74#_M1028_g N_Q_c_2349_n 6.05976e-19 $X=14.155 $Y=0.69 $X2=0
+ $Y2=0
cc_1183 N_A_2463_74#_c_1716_n N_Q_c_2349_n 0.01483f $X=15.07 $Y=1.28 $X2=0 $Y2=0
cc_1184 N_A_2463_74#_c_1718_n N_Q_c_2349_n 0.00388121f $X=15.145 $Y=1.205 $X2=0
+ $Y2=0
cc_1185 N_A_2463_74#_c_1720_n N_Q_c_2349_n 0.00584749f $X=15.3 $Y=1.675 $X2=0
+ $Y2=0
cc_1186 N_A_2463_74#_c_1729_n N_Q_c_2349_n 0.00177084f $X=15.3 $Y=1.765 $X2=0
+ $Y2=0
cc_1187 N_A_2463_74#_c_1727_n Q 0.00115341f $X=14.29 $Y=1.885 $X2=0 $Y2=0
cc_1188 N_A_2463_74#_c_1716_n Q 0.00341878f $X=15.07 $Y=1.28 $X2=0 $Y2=0
cc_1189 N_A_2463_74#_c_1729_n Q 0.00308602f $X=15.3 $Y=1.765 $X2=0 $Y2=0
cc_1190 N_A_2463_74#_c_1729_n Q 0.0114593f $X=15.3 $Y=1.765 $X2=0 $Y2=0
cc_1191 N_A_2463_74#_c_1722_n N_VGND_M1032_d 0.00829009f $X=13.705 $Y=0.855
+ $X2=0 $Y2=0
cc_1192 N_A_2463_74#_c_1723_n N_VGND_M1032_d 7.68198e-19 $X=13.79 $Y=1.2 $X2=0
+ $Y2=0
cc_1193 N_A_2463_74#_c_1721_n N_VGND_c_2403_n 0.010811f $X=12.455 $Y=0.515 $X2=0
+ $Y2=0
cc_1194 N_A_2463_74#_c_1718_n N_VGND_c_2404_n 0.00244473f $X=15.145 $Y=1.205
+ $X2=0 $Y2=0
cc_1195 N_A_2463_74#_M1028_g N_VGND_c_2414_n 0.00430908f $X=14.155 $Y=0.69 $X2=0
+ $Y2=0
cc_1196 N_A_2463_74#_c_1718_n N_VGND_c_2414_n 9.78499e-19 $X=15.145 $Y=1.205
+ $X2=0 $Y2=0
cc_1197 N_A_2463_74#_M1028_g N_VGND_c_2416_n 0.00825434f $X=14.155 $Y=0.69 $X2=0
+ $Y2=0
cc_1198 N_A_2463_74#_c_1721_n N_VGND_c_2416_n 0.0119404f $X=12.455 $Y=0.515
+ $X2=0 $Y2=0
cc_1199 N_A_2463_74#_c_1722_n N_VGND_c_2416_n 0.021428f $X=13.705 $Y=0.855 $X2=0
+ $Y2=0
cc_1200 N_A_2463_74#_c_1721_n N_VGND_c_2422_n 0.014415f $X=12.455 $Y=0.515 $X2=0
+ $Y2=0
cc_1201 N_A_2463_74#_M1028_g N_VGND_c_2423_n 0.00777377f $X=14.155 $Y=0.69 $X2=0
+ $Y2=0
cc_1202 N_A_2463_74#_c_1717_n N_VGND_c_2423_n 0.00115735f $X=14.38 $Y=1.28 $X2=0
+ $Y2=0
cc_1203 N_A_2463_74#_c_1721_n N_VGND_c_2423_n 0.00419512f $X=12.455 $Y=0.515
+ $X2=0 $Y2=0
cc_1204 N_A_2463_74#_c_1722_n N_VGND_c_2423_n 0.0501494f $X=13.705 $Y=0.855
+ $X2=0 $Y2=0
cc_1205 N_A_2463_74#_c_1725_n N_VGND_c_2423_n 0.00507997f $X=14.13 $Y=1.365
+ $X2=0 $Y2=0
cc_1206 N_A_2463_74#_c_1722_n A_2565_74# 0.0023798f $X=13.705 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_1207 N_A_27_90#_c_1876_n A_116_464# 0.0048076f $X=1.375 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_1208 N_A_27_90#_c_1876_n N_VPWR_M1029_d 0.00509381f $X=1.375 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_1209 N_A_27_90#_c_1878_n N_VPWR_M1019_d 5.2468e-19 $X=2.055 $Y=2.99 $X2=0
+ $Y2=0
cc_1210 N_A_27_90#_c_1908_n N_VPWR_M1019_d 0.00471831f $X=2.14 $Y=2.905 $X2=0
+ $Y2=0
cc_1211 N_A_27_90#_c_1880_n N_VPWR_M1019_d 0.00680034f $X=3.185 $Y=2.395 $X2=0
+ $Y2=0
cc_1212 N_A_27_90#_c_1875_n N_VPWR_c_1992_n 0.0104837f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_1213 N_A_27_90#_c_1876_n N_VPWR_c_1992_n 0.0154248f $X=1.375 $Y=2.375 $X2=0
+ $Y2=0
cc_1214 N_A_27_90#_c_1877_n N_VPWR_c_1992_n 0.0208967f $X=1.46 $Y=2.905 $X2=0
+ $Y2=0
cc_1215 N_A_27_90#_c_1879_n N_VPWR_c_1992_n 0.0146662f $X=1.545 $Y=2.99 $X2=0
+ $Y2=0
cc_1216 N_A_27_90#_c_1878_n N_VPWR_c_1993_n 0.0145682f $X=2.055 $Y=2.99 $X2=0
+ $Y2=0
cc_1217 N_A_27_90#_c_1908_n N_VPWR_c_1993_n 0.0190357f $X=2.14 $Y=2.905 $X2=0
+ $Y2=0
cc_1218 N_A_27_90#_c_1880_n N_VPWR_c_1993_n 0.0150987f $X=3.185 $Y=2.395 $X2=0
+ $Y2=0
cc_1219 N_A_27_90#_c_1884_n N_VPWR_c_1993_n 0.00946102f $X=3.35 $Y=2.475 $X2=0
+ $Y2=0
cc_1220 N_A_27_90#_c_1875_n N_VPWR_c_2001_n 0.0146013f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_1221 N_A_27_90#_c_1878_n N_VPWR_c_2002_n 0.0445209f $X=2.055 $Y=2.99 $X2=0
+ $Y2=0
cc_1222 N_A_27_90#_c_1879_n N_VPWR_c_2002_n 0.0121867f $X=1.545 $Y=2.99 $X2=0
+ $Y2=0
cc_1223 N_A_27_90#_c_1884_n N_VPWR_c_2003_n 0.0157912f $X=3.35 $Y=2.475 $X2=0
+ $Y2=0
cc_1224 N_A_27_90#_c_1875_n N_VPWR_c_1991_n 0.0120495f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_1225 N_A_27_90#_c_1878_n N_VPWR_c_1991_n 0.0250929f $X=2.055 $Y=2.99 $X2=0
+ $Y2=0
cc_1226 N_A_27_90#_c_1879_n N_VPWR_c_1991_n 0.00660921f $X=1.545 $Y=2.99 $X2=0
+ $Y2=0
cc_1227 N_A_27_90#_c_1880_n N_VPWR_c_1991_n 0.0232051f $X=3.185 $Y=2.395 $X2=0
+ $Y2=0
cc_1228 N_A_27_90#_c_1884_n N_VPWR_c_1991_n 0.0128787f $X=3.35 $Y=2.475 $X2=0
+ $Y2=0
cc_1229 N_A_27_90#_c_1880_n A_556_464# 0.00316297f $X=3.185 $Y=2.395 $X2=-0.19
+ $Y2=-0.245
cc_1230 N_A_27_90#_c_1884_n N_A_697_113#_c_2180_n 0.0137059f $X=3.35 $Y=2.475
+ $X2=0 $Y2=0
cc_1231 N_A_27_90#_c_1884_n N_A_697_113#_c_2181_n 0.0324354f $X=3.35 $Y=2.475
+ $X2=0 $Y2=0
cc_1232 N_A_27_90#_c_1884_n N_A_697_113#_c_2183_n 0.00626619f $X=3.35 $Y=2.475
+ $X2=0 $Y2=0
cc_1233 N_A_27_90#_c_1870_n N_A_697_113#_c_2177_n 0.0188588f $X=3.195 $Y=0.775
+ $X2=0 $Y2=0
cc_1234 N_A_27_90#_c_1873_n N_A_697_113#_c_2177_n 0.00109257f $X=3.46 $Y=1.26
+ $X2=0 $Y2=0
cc_1235 N_A_27_90#_c_1870_n N_A_697_113#_c_2178_n 0.00689028f $X=3.195 $Y=0.775
+ $X2=0 $Y2=0
cc_1236 N_A_27_90#_c_1871_n N_A_697_113#_c_2178_n 0.0712086f $X=3.46 $Y=2.31
+ $X2=0 $Y2=0
cc_1237 N_A_27_90#_c_1873_n N_A_697_113#_c_2178_n 0.0135923f $X=3.46 $Y=1.26
+ $X2=0 $Y2=0
cc_1238 N_A_27_90#_c_1872_n N_VGND_c_2397_n 0.0108279f $X=0.495 $Y=0.645 $X2=0
+ $Y2=0
cc_1239 N_A_27_90#_c_1870_n N_VGND_c_2398_n 0.0145731f $X=3.195 $Y=0.775 $X2=0
+ $Y2=0
cc_1240 N_A_27_90#_c_1872_n N_VGND_c_2409_n 0.0138602f $X=0.495 $Y=0.645 $X2=0
+ $Y2=0
cc_1241 N_A_27_90#_c_1870_n N_VGND_c_2410_n 0.00794834f $X=3.195 $Y=0.775 $X2=0
+ $Y2=0
cc_1242 N_A_27_90#_c_1870_n N_VGND_c_2416_n 0.0105391f $X=3.195 $Y=0.775 $X2=0
+ $Y2=0
cc_1243 N_A_27_90#_c_1872_n N_VGND_c_2416_n 0.0179195f $X=0.495 $Y=0.645 $X2=0
+ $Y2=0
cc_1244 N_VPWR_M1003_d N_A_697_113#_c_2182_n 4.29284e-19 $X=4.725 $Y=2.31 $X2=0
+ $Y2=0
cc_1245 N_VPWR_c_1994_n N_A_697_113#_c_2182_n 0.0145995f $X=5.04 $Y=2.8 $X2=0
+ $Y2=0
cc_1246 N_VPWR_c_2003_n N_A_697_113#_c_2182_n 0.0516485f $X=4.955 $Y=3.33 $X2=0
+ $Y2=0
cc_1247 N_VPWR_c_1991_n N_A_697_113#_c_2182_n 0.027478f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1248 N_VPWR_c_2003_n N_A_697_113#_c_2183_n 0.0170431f $X=4.955 $Y=3.33 $X2=0
+ $Y2=0
cc_1249 N_VPWR_c_1991_n N_A_697_113#_c_2183_n 0.00857552f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1250 N_VPWR_M1003_d N_A_697_113#_c_2208_n 0.00490162f $X=4.725 $Y=2.31 $X2=0
+ $Y2=0
cc_1251 N_VPWR_c_1994_n N_A_697_113#_c_2208_n 0.0205314f $X=5.04 $Y=2.8 $X2=0
+ $Y2=0
cc_1252 N_VPWR_M1034_s N_A_697_113#_c_2186_n 0.00676213f $X=6.295 $Y=1.84 $X2=0
+ $Y2=0
cc_1253 N_VPWR_M1008_s N_A_697_113#_c_2186_n 0.00225423f $X=7.685 $Y=1.84 $X2=0
+ $Y2=0
cc_1254 N_VPWR_c_1995_n N_A_697_113#_c_2186_n 0.02081f $X=6.44 $Y=2.815 $X2=0
+ $Y2=0
cc_1255 N_VPWR_c_1996_n N_A_697_113#_c_2186_n 0.00841219f $X=7.83 $Y=2.815 $X2=0
+ $Y2=0
cc_1256 N_VPWR_c_1991_n N_A_697_113#_c_2186_n 0.0367827f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1257 N_VPWR_M1008_s N_A_697_113#_c_2187_n 0.0107829f $X=7.685 $Y=1.84 $X2=0
+ $Y2=0
cc_1258 N_VPWR_c_1996_n N_A_697_113#_c_2200_n 9.6946e-19 $X=7.83 $Y=2.815 $X2=0
+ $Y2=0
cc_1259 N_VPWR_c_1991_n N_A_697_113#_c_2200_n 0.0050195f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1260 N_VPWR_c_1996_n N_A_697_113#_c_2188_n 0.0103109f $X=7.83 $Y=2.815 $X2=0
+ $Y2=0
cc_1261 N_VPWR_c_2006_n N_A_697_113#_c_2188_n 0.00757735f $X=10.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1262 N_VPWR_c_1991_n N_A_697_113#_c_2188_n 0.00627549f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1263 N_VPWR_c_2006_n N_A_697_113#_c_2189_n 0.0283027f $X=10.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1264 N_VPWR_c_1991_n N_A_697_113#_c_2189_n 0.0244128f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1265 N_VPWR_c_1994_n N_A_697_113#_c_2191_n 0.0101841f $X=5.04 $Y=2.8 $X2=0
+ $Y2=0
cc_1266 N_VPWR_c_1995_n N_A_697_113#_c_2191_n 0.021574f $X=6.44 $Y=2.815 $X2=0
+ $Y2=0
cc_1267 N_VPWR_c_2004_n N_A_697_113#_c_2191_n 0.0137032f $X=6.275 $Y=3.33 $X2=0
+ $Y2=0
cc_1268 N_VPWR_c_1991_n N_A_697_113#_c_2191_n 0.0118961f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1269 N_VPWR_M1003_d N_A_697_113#_c_2192_n 0.00923394f $X=4.725 $Y=2.31 $X2=0
+ $Y2=0
cc_1270 N_VPWR_c_1994_n N_A_697_113#_c_2192_n 0.0148828f $X=5.04 $Y=2.8 $X2=0
+ $Y2=0
cc_1271 N_VPWR_c_1991_n N_A_697_113#_c_2193_n 0.0080067f $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1272 N_VPWR_M1008_s N_A_697_113#_c_2333_n 0.00184106f $X=7.685 $Y=1.84 $X2=0
+ $Y2=0
cc_1273 N_VPWR_c_1996_n N_A_697_113#_c_2333_n 0.0126027f $X=7.83 $Y=2.815 $X2=0
+ $Y2=0
cc_1274 N_VPWR_c_1991_n N_A_697_113#_c_2333_n 6.0606e-19 $X=16.08 $Y=3.33 $X2=0
+ $Y2=0
cc_1275 N_VPWR_c_2000_n Q 0.0788705f $X=15.525 $Y=1.985 $X2=0 $Y2=0
cc_1276 N_VPWR_c_2009_n Q 0.0174942f $X=15.44 $Y=3.33 $X2=0 $Y2=0
cc_1277 N_VPWR_c_1991_n Q 0.0144473f $X=16.08 $Y=3.33 $X2=0 $Y2=0
cc_1278 N_VPWR_c_2000_n Q_N 0.0458635f $X=15.525 $Y=1.985 $X2=0 $Y2=0
cc_1279 N_VPWR_c_2010_n Q_N 0.0166018f $X=16.08 $Y=3.33 $X2=0 $Y2=0
cc_1280 N_VPWR_c_1991_n Q_N 0.0137086f $X=16.08 $Y=3.33 $X2=0 $Y2=0
cc_1281 N_A_697_113#_c_2192_n A_1068_462# 0.0048076f $X=5.715 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_1282 N_A_697_113#_c_2179_n N_VGND_c_2399_n 0.0129196f $X=6.125 $Y=0.807 $X2=0
+ $Y2=0
cc_1283 N_A_697_113#_c_2179_n N_VGND_c_2400_n 0.0324845f $X=6.125 $Y=0.807 $X2=0
+ $Y2=0
cc_1284 N_A_697_113#_c_2179_n N_VGND_c_2407_n 0.00967672f $X=6.125 $Y=0.807
+ $X2=0 $Y2=0
cc_1285 N_A_697_113#_c_2177_n N_VGND_c_2410_n 0.00859936f $X=3.695 $Y=0.775
+ $X2=0 $Y2=0
cc_1286 N_A_697_113#_c_2177_n N_VGND_c_2416_n 0.0113392f $X=3.695 $Y=0.775 $X2=0
+ $Y2=0
cc_1287 N_A_697_113#_c_2179_n N_VGND_c_2416_n 0.0141076f $X=6.125 $Y=0.807 $X2=0
+ $Y2=0
cc_1288 N_Q_N_c_2375_n N_VGND_c_2404_n 0.0296679f $X=16.04 $Y=0.535 $X2=0 $Y2=0
cc_1289 N_Q_N_c_2375_n N_VGND_c_2415_n 0.0147163f $X=16.04 $Y=0.535 $X2=0 $Y2=0
cc_1290 N_Q_N_c_2375_n N_VGND_c_2416_n 0.0130412f $X=16.04 $Y=0.535 $X2=0 $Y2=0
