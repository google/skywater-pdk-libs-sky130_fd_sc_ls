# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ls__o32a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__o32a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845000 1.120000 7.295000 1.410000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.075000 1.130000 6.405000 1.580000 ;
        RECT 6.075000 1.580000 8.035000 1.780000 ;
        RECT 6.075000 1.780000 6.405000 1.800000 ;
        RECT 7.565000 1.450000 8.035000 1.580000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.065000 1.180000 5.735000 1.510000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.450000 2.855000 1.780000 ;
        RECT 2.685000 1.780000 2.855000 2.360000 ;
        RECT 2.685000 2.360000 5.905000 2.530000 ;
        RECT 4.495000 1.450000 4.825000 1.680000 ;
        RECT 4.495000 1.680000 5.905000 1.850000 ;
        RECT 5.735000 1.850000 5.905000 2.360000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.925000 1.270000 4.255000 1.780000 ;
    END
  END B2
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 8.160000 0.245000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 8.350000 3.520000 ;
    END
  END VPB
  PIN X
    ANTENNADIFFAREA  1.313300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.140000 1.015000 1.310000 ;
        RECT 0.125000 1.310000 0.355000 1.480000 ;
        RECT 0.125000 1.480000 0.895000 1.650000 ;
        RECT 0.565000 1.650000 0.895000 1.780000 ;
        RECT 0.565000 1.780000 1.895000 1.950000 ;
        RECT 0.565000 1.950000 0.895000 2.980000 ;
        RECT 0.685000 0.350000 1.015000 0.940000 ;
        RECT 0.685000 0.940000 2.015000 1.110000 ;
        RECT 0.685000 1.110000 1.015000 1.140000 ;
        RECT 1.565000 1.950000 1.895000 2.980000 ;
        RECT 1.685000 0.350000 2.015000 0.940000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.185000  0.085000 0.515000 0.970000 ;
      RECT 1.065000  2.120000 1.395000 3.245000 ;
      RECT 1.185000  0.085000 1.515000 0.770000 ;
      RECT 1.255000  1.280000 2.355000 1.610000 ;
      RECT 2.085000  1.950000 2.415000 3.245000 ;
      RECT 2.185000  1.110000 3.560000 1.280000 ;
      RECT 2.240000  0.085000 2.570000 0.940000 ;
      RECT 2.655000  2.700000 4.025000 2.960000 ;
      RECT 2.800000  0.255000 5.060000 0.425000 ;
      RECT 2.800000  0.425000 3.130000 0.940000 ;
      RECT 3.230000  1.280000 3.560000 1.920000 ;
      RECT 3.230000  1.920000 3.575000 2.020000 ;
      RECT 3.230000  2.020000 5.565000 2.190000 ;
      RECT 3.300000  0.595000 3.560000 0.930000 ;
      RECT 3.300000  0.930000 4.560000 1.100000 ;
      RECT 3.300000  1.100000 3.560000 1.110000 ;
      RECT 3.730000  0.425000 4.060000 0.760000 ;
      RECT 4.195000  2.700000 4.525000 3.245000 ;
      RECT 4.230000  0.595000 4.560000 0.930000 ;
      RECT 4.730000  0.425000 5.060000 0.790000 ;
      RECT 4.730000  0.790000 8.045000 0.950000 ;
      RECT 4.730000  0.950000 6.060000 0.960000 ;
      RECT 4.730000  0.960000 5.060000 1.010000 ;
      RECT 4.785000  2.700000 6.245000 2.980000 ;
      RECT 5.230000  0.085000 5.560000 0.620000 ;
      RECT 5.730000  0.350000 6.060000 0.780000 ;
      RECT 5.730000  0.780000 8.045000 0.790000 ;
      RECT 6.075000  2.390000 8.045000 2.560000 ;
      RECT 6.075000  2.560000 6.245000 2.700000 ;
      RECT 6.155000  1.970000 7.595000 2.200000 ;
      RECT 6.155000  2.200000 6.675000 2.220000 ;
      RECT 6.230000  0.085000 6.560000 0.610000 ;
      RECT 6.740000  0.350000 6.990000 0.780000 ;
      RECT 6.805000  2.730000 7.135000 3.245000 ;
      RECT 7.160000  0.085000 7.545000 0.600000 ;
      RECT 7.265000  1.950000 7.595000 1.970000 ;
      RECT 7.715000  0.350000 8.045000 0.780000 ;
      RECT 7.715000  0.950000 8.045000 1.030000 ;
      RECT 7.715000  2.560000 8.045000 2.980000 ;
      RECT 7.765000  1.950000 8.045000 2.390000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_ls__o32a_4
END LIBRARY
