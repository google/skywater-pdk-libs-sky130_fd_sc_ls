* File: sky130_fd_sc_ls__o2111a_4.pex.spice
* Created: Wed Sep  2 11:16:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O2111A_4%D1 3 5 7 8 12 14 16 17 19 23
c57 17 0 7.68806e-20 $X=0.93 $Y=1.757
r58 22 24 13.2661 $w=3.27e-07 $l=9e-08 $layer=POLY_cond $X=0.407 $Y=1.615
+ $X2=0.407 $Y2=1.705
r59 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.615 $X2=0.385 $Y2=1.615
r60 19 23 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.385 $Y2=1.615
r61 17 18 28.0233 $w=2.15e-07 $l=1.25e-07 $layer=POLY_cond $X=0.93 $Y=1.757
+ $X2=1.055 $Y2=1.757
r62 14 18 11.2427 $w=1.5e-07 $l=1.28e-07 $layer=POLY_cond $X=1.055 $Y=1.885
+ $X2=1.055 $Y2=1.757
r63 14 16 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.055 $Y=1.885
+ $X2=1.055 $Y2=2.38
r64 10 17 11.2427 $w=1.5e-07 $l=1.27e-07 $layer=POLY_cond $X=0.93 $Y=1.63
+ $X2=0.93 $Y2=1.757
r65 10 12 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=0.93 $Y=1.63
+ $X2=0.93 $Y2=0.74
r66 9 24 21.0057 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=0.595 $Y=1.705
+ $X2=0.407 $Y2=1.705
r67 8 17 21.2711 $w=2.15e-07 $l=9.75961e-08 $layer=POLY_cond $X=0.855 $Y=1.705
+ $X2=0.93 $Y2=1.757
r68 8 9 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=0.855 $Y=1.705
+ $X2=0.595 $Y2=1.705
r69 5 24 40.7928 $w=3.27e-07 $l=2.23696e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.407 $Y2=1.705
r70 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.38
r71 1 22 38.5818 $w=3.27e-07 $l=2.06325e-07 $layer=POLY_cond $X=0.5 $Y=1.45
+ $X2=0.407 $Y2=1.615
r72 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.5 $Y=1.45 $X2=0.5
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_4%C1 1 3 4 6 7 9 10 12 13 14 22
r52 22 23 20.9354 $w=4.95e-07 $l=2.15e-07 $layer=POLY_cond $X=1.79 $Y=1.535
+ $X2=2.005 $Y2=1.535
r53 20 22 20.4485 $w=4.95e-07 $l=2.1e-07 $layer=POLY_cond $X=1.58 $Y=1.535
+ $X2=1.79 $Y2=1.535
r54 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.58
+ $Y=1.615 $X2=1.58 $Y2=1.615
r55 18 20 7.30303 $w=4.95e-07 $l=7.5e-08 $layer=POLY_cond $X=1.505 $Y=1.535
+ $X2=1.58 $Y2=1.535
r56 14 21 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.68 $Y=1.615 $X2=1.58
+ $Y2=1.615
r57 13 21 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.58 $Y2=1.615
r58 10 23 31.1543 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.005 $Y=1.885
+ $X2=2.005 $Y2=1.535
r59 10 12 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.005 $Y=1.885
+ $X2=2.005 $Y2=2.38
r60 7 22 31.1543 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.79 $Y=1.185
+ $X2=1.79 $Y2=1.535
r61 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.79 $Y=1.185
+ $X2=1.79 $Y2=0.74
r62 4 18 31.1543 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.505 $Y=1.885
+ $X2=1.505 $Y2=1.535
r63 4 6 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.505 $Y=1.885
+ $X2=1.505 $Y2=2.38
r64 1 18 14.1192 $w=4.95e-07 $l=4.16233e-07 $layer=POLY_cond $X=1.36 $Y=1.185
+ $X2=1.505 $Y2=1.535
r65 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.36 $Y=1.185
+ $X2=1.36 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_4%B1 1 3 6 8 10 13 15 21
c50 13 0 2.37497e-19 $X=3.255 $Y=0.91
r51 21 23 15.4299 $w=3.28e-07 $l=1.05e-07 $layer=POLY_cond $X=3.15 $Y=1.667
+ $X2=3.255 $Y2=1.667
r52 19 21 11.0213 $w=3.28e-07 $l=7.5e-08 $layer=POLY_cond $X=3.075 $Y=1.667
+ $X2=3.15 $Y2=1.667
r53 18 19 36.7378 $w=3.28e-07 $l=2.5e-07 $layer=POLY_cond $X=2.825 $Y=1.667
+ $X2=3.075 $Y2=1.667
r54 17 18 29.3902 $w=3.28e-07 $l=2e-07 $layer=POLY_cond $X=2.625 $Y=1.667
+ $X2=2.825 $Y2=1.667
r55 15 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.15
+ $Y=1.615 $X2=3.15 $Y2=1.615
r56 11 23 21.0783 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=3.255 $Y=1.45
+ $X2=3.255 $Y2=1.667
r57 11 13 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=3.255 $Y=1.45
+ $X2=3.255 $Y2=0.91
r58 8 19 21.0783 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=3.075 $Y=1.885
+ $X2=3.075 $Y2=1.667
r59 8 10 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.075 $Y=1.885
+ $X2=3.075 $Y2=2.38
r60 4 18 21.0783 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=2.825 $Y=1.45
+ $X2=2.825 $Y2=1.667
r61 4 6 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.825 $Y=1.45
+ $X2=2.825 $Y2=0.91
r62 1 17 21.0783 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=2.625 $Y=1.885
+ $X2=2.625 $Y2=1.667
r63 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.625 $Y=1.885
+ $X2=2.625 $Y2=2.38
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_4%A2 1 3 6 8 10 13 15 16 17 18 28
r51 28 29 1.87792 $w=3.85e-07 $l=1.5e-08 $layer=POLY_cond $X=4.16 $Y=1.667
+ $X2=4.175 $Y2=1.667
r52 26 28 10.6416 $w=3.85e-07 $l=8.5e-08 $layer=POLY_cond $X=4.075 $Y=1.667
+ $X2=4.16 $Y2=1.667
r53 24 26 48.826 $w=3.85e-07 $l=3.9e-07 $layer=POLY_cond $X=3.685 $Y=1.667
+ $X2=4.075 $Y2=1.667
r54 23 24 3.12987 $w=3.85e-07 $l=2.5e-08 $layer=POLY_cond $X=3.66 $Y=1.667
+ $X2=3.685 $Y2=1.667
r55 17 18 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.615
+ $X2=5.04 $Y2=1.615
r56 16 17 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=4.075 $Y=1.615
+ $X2=4.56 $Y2=1.615
r57 16 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.075
+ $Y=1.615 $X2=4.075 $Y2=1.615
r58 15 16 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=3.6 $Y=1.615
+ $X2=4.075 $Y2=1.615
r59 11 29 24.9301 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=4.175 $Y=1.45
+ $X2=4.175 $Y2=1.667
r60 11 13 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=4.175 $Y=1.45
+ $X2=4.175 $Y2=0.91
r61 8 28 24.9301 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=4.16 $Y=1.885
+ $X2=4.16 $Y2=1.667
r62 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.16 $Y=1.885
+ $X2=4.16 $Y2=2.46
r63 4 24 24.9301 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=3.685 $Y=1.45
+ $X2=3.685 $Y2=1.667
r64 4 6 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=3.685 $Y=1.45
+ $X2=3.685 $Y2=0.91
r65 1 23 24.9301 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=3.66 $Y=1.885
+ $X2=3.66 $Y2=1.667
r66 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.66 $Y=1.885
+ $X2=3.66 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_4%A1 3 5 7 10 12 14 15 22
c48 15 0 1.3655e-20 $X=5.52 $Y=1.665
c49 10 0 3.86387e-19 $X=5.635 $Y=0.74
r50 22 23 4.43947 $w=3.8e-07 $l=3.5e-08 $layer=POLY_cond $X=5.635 $Y=1.667
+ $X2=5.67 $Y2=1.667
r51 20 22 18.3921 $w=3.8e-07 $l=1.45e-07 $layer=POLY_cond $X=5.49 $Y=1.667
+ $X2=5.635 $Y2=1.667
r52 18 20 34.2474 $w=3.8e-07 $l=2.7e-07 $layer=POLY_cond $X=5.22 $Y=1.667
+ $X2=5.49 $Y2=1.667
r53 17 18 1.90263 $w=3.8e-07 $l=1.5e-08 $layer=POLY_cond $X=5.205 $Y=1.667
+ $X2=5.22 $Y2=1.667
r54 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.49
+ $Y=1.615 $X2=5.49 $Y2=1.615
r55 12 23 24.6126 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=5.67 $Y=1.885
+ $X2=5.67 $Y2=1.667
r56 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.67 $Y=1.885
+ $X2=5.67 $Y2=2.46
r57 8 22 24.6126 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=5.635 $Y=1.45
+ $X2=5.635 $Y2=1.667
r58 8 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.635 $Y=1.45
+ $X2=5.635 $Y2=0.74
r59 5 18 24.6126 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=5.22 $Y=1.885
+ $X2=5.22 $Y2=1.667
r60 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.22 $Y=1.885
+ $X2=5.22 $Y2=2.46
r61 1 17 24.6126 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=5.205 $Y=1.45
+ $X2=5.205 $Y2=1.667
r62 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.205 $Y=1.45
+ $X2=5.205 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_4%A_27_392# 1 2 3 4 5 6 21 23 25 28 30 32 35
+ 37 39 40 41 44 47 48 50 51 54 57 58 62 66 71 72 74 75 77 78 83 87 89 92 94 96
+ 98 100
c223 78 0 1.58594e-19 $X=6.145 $Y=1.515
c224 23 0 1.5326e-19 $X=6.205 $Y=1.765
r225 110 111 2.67778 $w=3.6e-07 $l=2e-08 $layer=POLY_cond $X=7.135 $Y=1.557
+ $X2=7.155 $Y2=1.557
r226 107 108 18.7444 $w=3.6e-07 $l=1.4e-07 $layer=POLY_cond $X=6.565 $Y=1.557
+ $X2=6.705 $Y2=1.557
r227 104 105 9.37222 $w=3.6e-07 $l=7e-08 $layer=POLY_cond $X=6.135 $Y=1.557
+ $X2=6.205 $Y2=1.557
r228 100 102 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.385 $Y=2.805
+ $X2=4.385 $Y2=2.99
r229 89 91 8.98035 $w=3.38e-07 $l=1.8e-07 $layer=LI1_cond $X=0.72 $Y=0.95
+ $X2=0.72 $Y2=1.13
r230 84 110 23.4306 $w=3.6e-07 $l=1.75e-07 $layer=POLY_cond $X=6.96 $Y=1.557
+ $X2=7.135 $Y2=1.557
r231 84 108 34.1417 $w=3.6e-07 $l=2.55e-07 $layer=POLY_cond $X=6.96 $Y=1.557
+ $X2=6.705 $Y2=1.557
r232 83 84 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.96
+ $Y=1.515 $X2=6.96 $Y2=1.515
r233 81 107 38.1583 $w=3.6e-07 $l=2.85e-07 $layer=POLY_cond $X=6.28 $Y=1.557
+ $X2=6.565 $Y2=1.557
r234 81 105 10.0417 $w=3.6e-07 $l=7.5e-08 $layer=POLY_cond $X=6.28 $Y=1.557
+ $X2=6.205 $Y2=1.557
r235 80 83 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.28 $Y=1.515
+ $X2=6.96 $Y2=1.515
r236 80 81 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.28
+ $Y=1.515 $X2=6.28 $Y2=1.515
r237 78 80 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.145 $Y=1.515
+ $X2=6.28 $Y2=1.515
r238 76 78 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.06 $Y=1.68
+ $X2=6.145 $Y2=1.515
r239 76 77 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.06 $Y=1.68
+ $X2=6.06 $Y2=1.95
r240 74 102 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.22 $Y=2.99
+ $X2=4.385 $Y2=2.99
r241 74 75 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.22 $Y=2.99
+ $X2=3.55 $Y2=2.99
r242 73 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=2.035
+ $X2=3.385 $Y2=2.035
r243 72 77 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.975 $Y=2.035
+ $X2=6.06 $Y2=1.95
r244 72 73 158.209 $w=1.68e-07 $l=2.425e-06 $layer=LI1_cond $X=5.975 $Y=2.035
+ $X2=3.55 $Y2=2.035
r245 69 75 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.385 $Y=2.905
+ $X2=3.55 $Y2=2.99
r246 69 71 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.385 $Y=2.905
+ $X2=3.385 $Y2=2.815
r247 68 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=2.12
+ $X2=3.385 $Y2=2.035
r248 68 71 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.385 $Y=2.12
+ $X2=3.385 $Y2=2.815
r249 67 96 8.61065 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=2.48 $Y=2.035
+ $X2=2.315 $Y2=2.03
r250 66 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.22 $Y=2.035
+ $X2=3.385 $Y2=2.035
r251 66 67 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.22 $Y=2.035
+ $X2=2.48 $Y2=2.035
r252 63 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=2.035
+ $X2=1.28 $Y2=2.035
r253 62 96 8.61065 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=2.15 $Y=2.035
+ $X2=2.315 $Y2=2.03
r254 62 63 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.15 $Y=2.035
+ $X2=1.445 $Y2=2.035
r255 59 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=2.035
+ $X2=0.805 $Y2=2.035
r256 58 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=2.035
+ $X2=1.28 $Y2=2.035
r257 58 59 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.115 $Y=2.035
+ $X2=0.89 $Y2=2.035
r258 57 92 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=1.95
+ $X2=0.805 $Y2=2.035
r259 57 91 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.805 $Y=1.95
+ $X2=0.805 $Y2=1.13
r260 55 87 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r261 54 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.035
+ $X2=0.805 $Y2=2.035
r262 54 55 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.72 $Y=2.035
+ $X2=0.445 $Y2=2.035
r263 48 50 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.605 $Y=1.765
+ $X2=7.605 $Y2=2.4
r264 47 48 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.605 $Y=1.675
+ $X2=7.605 $Y2=1.765
r265 46 51 18.8402 $w=1.65e-07 $l=8.12404e-08 $layer=POLY_cond $X=7.605 $Y=1.5
+ $X2=7.592 $Y2=1.425
r266 46 47 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=7.605 $Y=1.5
+ $X2=7.605 $Y2=1.675
r267 42 51 18.8402 $w=1.65e-07 $l=8.74643e-08 $layer=POLY_cond $X=7.565 $Y=1.35
+ $X2=7.592 $Y2=1.425
r268 42 44 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.565 $Y=1.35
+ $X2=7.565 $Y2=0.74
r269 41 111 28.8686 $w=3.6e-07 $l=1.71184e-07 $layer=POLY_cond $X=7.245 $Y=1.425
+ $X2=7.155 $Y2=1.557
r270 40 51 6.66866 $w=1.5e-07 $l=1.02e-07 $layer=POLY_cond $X=7.49 $Y=1.425
+ $X2=7.592 $Y2=1.425
r271 40 41 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=7.49 $Y=1.425
+ $X2=7.245 $Y2=1.425
r272 37 111 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.155 $Y=1.765
+ $X2=7.155 $Y2=1.557
r273 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.155 $Y=1.765
+ $X2=7.155 $Y2=2.4
r274 33 110 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.135 $Y=1.35
+ $X2=7.135 $Y2=1.557
r275 33 35 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.135 $Y=1.35
+ $X2=7.135 $Y2=0.74
r276 30 108 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.705 $Y=1.765
+ $X2=6.705 $Y2=1.557
r277 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.705 $Y=1.765
+ $X2=6.705 $Y2=2.4
r278 26 107 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.565 $Y=1.35
+ $X2=6.565 $Y2=1.557
r279 26 28 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.565 $Y=1.35
+ $X2=6.565 $Y2=0.74
r280 23 105 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.205 $Y=1.765
+ $X2=6.205 $Y2=1.557
r281 23 25 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.205 $Y=1.765
+ $X2=6.205 $Y2=2.4
r282 19 104 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.135 $Y=1.35
+ $X2=6.135 $Y2=1.557
r283 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.135 $Y=1.35
+ $X2=6.135 $Y2=0.74
r284 6 100 600 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=4.235
+ $Y=1.96 $X2=4.385 $Y2=2.805
r285 5 98 300 $w=1.7e-07 $l=3.02738e-07 $layer=licon1_PDIFF $count=2 $X=3.15
+ $Y=1.96 $X2=3.385 $Y2=2.115
r286 5 71 600 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=3.15
+ $Y=1.96 $X2=3.385 $Y2=2.815
r287 4 96 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=2.08
+ $Y=1.96 $X2=2.315 $Y2=2.105
r288 3 94 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=1.13
+ $Y=1.96 $X2=1.28 $Y2=2.115
r289 2 87 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
r290 1 89 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.37 $X2=0.715 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_4%VPWR 1 2 3 4 5 6 7 24 26 30 34 38 42 46 48
+ 50 55 56 58 59 60 62 77 81 86 92 95 98 101 105
c123 24 0 7.68806e-20 $X=0.78 $Y=2.48
r124 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r125 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r126 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r127 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r128 93 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r129 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r130 90 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r131 90 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r132 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r133 87 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.095 $Y=3.33
+ $X2=6.93 $Y2=3.33
r134 87 89 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.095 $Y=3.33
+ $X2=7.44 $Y2=3.33
r135 86 104 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.937 $Y2=3.33
r136 86 89 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.44 $Y2=3.33
r137 85 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r138 85 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r139 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r140 82 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=3.33
+ $X2=5.98 $Y2=3.33
r141 82 84 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.145 $Y=3.33
+ $X2=6.48 $Y2=3.33
r142 81 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.765 $Y=3.33
+ $X2=6.93 $Y2=3.33
r143 81 84 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.765 $Y=3.33
+ $X2=6.48 $Y2=3.33
r144 80 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r145 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r146 77 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=3.33
+ $X2=5.98 $Y2=3.33
r147 77 79 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.815 $Y=3.33
+ $X2=5.52 $Y2=3.33
r148 76 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r149 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r150 72 75 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r151 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r152 70 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r153 70 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r154 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r155 67 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=1.78 $Y2=3.33
r156 67 69 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=2.64 $Y2=3.33
r157 65 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r158 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r159 62 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r160 62 64 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r161 60 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r162 60 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r163 58 75 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.78 $Y=3.33
+ $X2=4.56 $Y2=3.33
r164 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.78 $Y=3.33
+ $X2=4.945 $Y2=3.33
r165 57 79 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=5.11 $Y=3.33
+ $X2=5.52 $Y2=3.33
r166 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.11 $Y=3.33
+ $X2=4.945 $Y2=3.33
r167 55 69 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.685 $Y=3.33
+ $X2=2.64 $Y2=3.33
r168 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=3.33
+ $X2=2.85 $Y2=3.33
r169 54 72 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.015 $Y=3.33
+ $X2=3.12 $Y2=3.33
r170 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=3.33
+ $X2=2.85 $Y2=3.33
r171 50 53 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.88 $Y=1.985
+ $X2=7.88 $Y2=2.815
r172 48 104 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.88 $Y=3.245
+ $X2=7.937 $Y2=3.33
r173 48 53 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.88 $Y=3.245
+ $X2=7.88 $Y2=2.815
r174 44 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.93 $Y=3.245
+ $X2=6.93 $Y2=3.33
r175 44 46 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=6.93 $Y=3.245
+ $X2=6.93 $Y2=2.435
r176 40 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.98 $Y=3.245
+ $X2=5.98 $Y2=3.33
r177 40 42 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=5.98 $Y=3.245
+ $X2=5.98 $Y2=2.455
r178 36 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.945 $Y=3.245
+ $X2=4.945 $Y2=3.33
r179 36 38 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=4.945 $Y=3.245
+ $X2=4.945 $Y2=2.805
r180 32 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=3.245
+ $X2=2.85 $Y2=3.33
r181 32 34 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=2.85 $Y=3.245
+ $X2=2.85 $Y2=2.48
r182 28 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=3.245
+ $X2=1.78 $Y2=3.33
r183 28 30 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=1.78 $Y=3.245
+ $X2=1.78 $Y2=2.48
r184 27 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r185 26 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=3.33
+ $X2=1.78 $Y2=3.33
r186 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=3.33
+ $X2=0.945 $Y2=3.33
r187 22 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r188 22 24 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.48
r189 7 53 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=7.68
+ $Y=1.84 $X2=7.88 $Y2=2.815
r190 7 50 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=7.68
+ $Y=1.84 $X2=7.88 $Y2=1.985
r191 6 46 300 $w=1.7e-07 $l=6.65789e-07 $layer=licon1_PDIFF $count=2 $X=6.78
+ $Y=1.84 $X2=6.93 $Y2=2.435
r192 5 42 300 $w=1.7e-07 $l=6.01124e-07 $layer=licon1_PDIFF $count=2 $X=5.745
+ $Y=1.96 $X2=5.98 $Y2=2.455
r193 4 38 600 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=4.8
+ $Y=1.96 $X2=4.945 $Y2=2.805
r194 3 34 600 $w=1.7e-07 $l=5.90254e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.96 $X2=2.85 $Y2=2.48
r195 2 30 600 $w=1.7e-07 $l=6.11882e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.96 $X2=1.78 $Y2=2.48
r196 1 24 600 $w=1.7e-07 $l=6.11882e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.96 $X2=0.78 $Y2=2.48
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_4%A_747_392# 1 2 7 11 17
c23 17 0 1.39605e-19 $X=5.445 $Y=2.455
r24 11 14 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.885 $Y=2.375
+ $X2=3.885 $Y2=2.51
r25 8 11 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=2.375
+ $X2=3.885 $Y2=2.375
r26 7 17 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.28 $Y=2.375
+ $X2=5.445 $Y2=2.375
r27 7 8 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=5.28 $Y=2.375 $X2=4.05
+ $Y2=2.375
r28 2 17 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=5.295
+ $Y=1.96 $X2=5.445 $Y2=2.455
r29 1 14 600 $w=1.7e-07 $l=6.20484e-07 $layer=licon1_PDIFF $count=1 $X=3.735
+ $Y=1.96 $X2=3.885 $Y2=2.51
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_4%X 1 2 3 4 15 17 19 21 22 23 27 30 33 35 37
+ 38 41 43 46
c82 30 0 5.23076e-20 $X=7.42 $Y=1.85
c83 22 0 1.93862e-19 $X=6.515 $Y=1.095
c84 15 0 1.92524e-19 $X=6.35 $Y=0.515
r85 45 46 9.26965 $w=2.28e-07 $l=1.85e-07 $layer=LI1_cond $X=7.92 $Y=1.48
+ $X2=7.92 $Y2=1.295
r86 44 46 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=7.92 $Y=1.18
+ $X2=7.92 $Y2=1.295
r87 37 45 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.805 $Y=1.565
+ $X2=7.92 $Y2=1.48
r88 37 38 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.805 $Y=1.565
+ $X2=7.545 $Y2=1.565
r89 36 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.515 $Y=1.095
+ $X2=7.35 $Y2=1.095
r90 35 44 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.805 $Y=1.095
+ $X2=7.92 $Y2=1.18
r91 35 36 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.805 $Y=1.095
+ $X2=7.515 $Y2=1.095
r92 31 43 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=7.42 $Y=2.18
+ $X2=7.42 $Y2=2.015
r93 31 33 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=7.42 $Y=2.18
+ $X2=7.42 $Y2=2.4
r94 30 43 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=7.42 $Y=1.85
+ $X2=7.42 $Y2=2.015
r95 29 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.42 $Y=1.65
+ $X2=7.545 $Y2=1.565
r96 29 30 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=7.42 $Y=1.65 $X2=7.42
+ $Y2=1.85
r97 25 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.35 $Y=1.01 $X2=7.35
+ $Y2=1.095
r98 25 27 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=7.35 $Y=1.01
+ $X2=7.35 $Y2=0.515
r99 24 40 3.13803 $w=3.3e-07 $l=1.38e-07 $layer=LI1_cond $X=6.59 $Y=2.015
+ $X2=6.452 $Y2=2.015
r100 23 43 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=7.295 $Y=2.015
+ $X2=7.42 $Y2=2.015
r101 23 24 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=7.295 $Y=2.015
+ $X2=6.59 $Y2=2.015
r102 21 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.185 $Y=1.095
+ $X2=7.35 $Y2=1.095
r103 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.185 $Y=1.095
+ $X2=6.515 $Y2=1.095
r104 17 40 3.75199 $w=2.75e-07 $l=1.65e-07 $layer=LI1_cond $X=6.452 $Y=2.18
+ $X2=6.452 $Y2=2.015
r105 17 19 9.21954 $w=2.73e-07 $l=2.2e-07 $layer=LI1_cond $X=6.452 $Y=2.18
+ $X2=6.452 $Y2=2.4
r106 13 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.35 $Y=1.01
+ $X2=6.515 $Y2=1.095
r107 13 15 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=6.35 $Y=1.01
+ $X2=6.35 $Y2=0.515
r108 4 43 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=1.84 $X2=7.38 $Y2=1.985
r109 4 33 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=7.23
+ $Y=1.84 $X2=7.38 $Y2=2.4
r110 3 40 600 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.84 $X2=6.48 $Y2=2.015
r111 3 19 300 $w=1.7e-07 $l=6.5238e-07 $layer=licon1_PDIFF $count=2 $X=6.28
+ $Y=1.84 $X2=6.48 $Y2=2.4
r112 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.21
+ $Y=0.37 $X2=7.35 $Y2=0.515
r113 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.21
+ $Y=0.37 $X2=6.35 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_4%A_27_74# 1 2 3 10 12 14 18 25 27 28
r39 27 28 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=2.085 $Y=0.397
+ $X2=1.92 $Y2=0.397
r40 21 25 3.6114 $w=2.57e-07 $l=1.22327e-07 $layer=LI1_cond $X=1.23 $Y=0.34
+ $X2=1.145 $Y2=0.427
r41 21 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.23 $Y=0.34 $X2=1.92
+ $Y2=0.34
r42 16 25 2.87242 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=1.145 $Y=0.6
+ $X2=1.145 $Y2=0.427
r43 16 18 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.145 $Y=0.6
+ $X2=1.145 $Y2=0.965
r44 15 23 3.02949 $w=3.45e-07 $l=1.33e-07 $layer=LI1_cond $X=0.38 $Y=0.427
+ $X2=0.247 $Y2=0.427
r45 14 25 3.6114 $w=2.57e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=0.427
+ $X2=1.145 $Y2=0.427
r46 14 15 22.7148 $w=3.43e-07 $l=6.8e-07 $layer=LI1_cond $X=1.06 $Y=0.427
+ $X2=0.38 $Y2=0.427
r47 10 23 3.94061 $w=2.65e-07 $l=1.73e-07 $layer=LI1_cond $X=0.247 $Y=0.6
+ $X2=0.247 $Y2=0.427
r48 10 12 15.2209 $w=2.63e-07 $l=3.5e-07 $layer=LI1_cond $X=0.247 $Y=0.6
+ $X2=0.247 $Y2=0.95
r49 3 27 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.37 $X2=2.085 $Y2=0.375
r50 2 25 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.37 $X2=1.145 $Y2=0.515
r51 2 18 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.37 $X2=1.145 $Y2=0.965
r52 1 23 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
r53 1 12 182 $w=1.7e-07 $l=6.4846e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_4%A_287_74# 1 2 7 12 14
c29 14 0 1.44963e-19 $X=3.04 $Y=0.7
r30 14 16 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=3 $Y=0.7 $X2=3
+ $Y2=0.795
r31 10 12 9.7361 $w=5.33e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=0.862
+ $X2=1.74 $Y2=0.862
r32 7 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.875 $Y=0.795 $X2=3
+ $Y2=0.795
r33 7 12 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=2.875 $Y=0.795
+ $X2=1.74 $Y2=0.795
r34 2 14 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=2.9
+ $Y=0.54 $X2=3.04 $Y2=0.7
r35 1 10 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.37 $X2=1.575 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_4%A_477_198# 1 2 3 4 13 17 21 23 27 29 33 35
+ 36 37
c64 35 0 9.25343e-20 $X=2.775 $Y=1.175
r65 31 33 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.42 $Y=1.11
+ $X2=5.42 $Y2=0.515
r66 30 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.565 $Y=1.195
+ $X2=4.4 $Y2=1.195
r67 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.335 $Y=1.195
+ $X2=5.42 $Y2=1.11
r68 29 30 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.335 $Y=1.195
+ $X2=4.565 $Y2=1.195
r69 25 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.4 $Y=1.11 $X2=4.4
+ $Y2=1.195
r70 25 27 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=4.4 $Y=1.11 $X2=4.4
+ $Y2=0.685
r71 24 36 6.19399 $w=2e-07 $l=1.39194e-07 $layer=LI1_cond $X=3.555 $Y=1.195
+ $X2=3.43 $Y2=1.165
r72 23 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.235 $Y=1.195
+ $X2=4.4 $Y2=1.195
r73 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.235 $Y=1.195
+ $X2=3.555 $Y2=1.195
r74 19 36 0.552779 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=3.43 $Y=1.05
+ $X2=3.43 $Y2=1.165
r75 19 21 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=3.43 $Y=1.05
+ $X2=3.43 $Y2=0.685
r76 17 36 6.19399 $w=2e-07 $l=1.25e-07 $layer=LI1_cond $X=3.305 $Y=1.165
+ $X2=3.43 $Y2=1.165
r77 17 35 26.5563 $w=2.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.305 $Y=1.165
+ $X2=2.775 $Y2=1.165
r78 13 35 5.85606 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.65 $Y=1.175
+ $X2=2.775 $Y2=1.175
r79 13 15 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.65 $Y=1.175 $X2=2.57
+ $Y2=1.175
r80 4 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.28
+ $Y=0.37 $X2=5.42 $Y2=0.515
r81 3 27 91 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=2 $X=4.25
+ $Y=0.54 $X2=4.4 $Y2=0.685
r82 2 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.33
+ $Y=0.54 $X2=3.47 $Y2=0.685
r83 1 15 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.385
+ $Y=0.99 $X2=2.57 $Y2=1.135
.ends

.subckt PM_SKY130_FD_SC_LS__O2111A_4%VGND 1 2 3 4 5 18 22 26 30 32 34 37 38 40
+ 41 43 44 45 54 65 70 74
r99 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r100 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r101 68 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r102 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r103 65 73 4.67153 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=7.685 $Y=0
+ $X2=7.922 $Y2=0
r104 65 67 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.685 $Y=0 $X2=7.44
+ $Y2=0
r105 64 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r106 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r107 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r108 61 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r109 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r110 58 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.155 $Y=0 $X2=4.99
+ $Y2=0
r111 58 60 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.155 $Y=0
+ $X2=5.52 $Y2=0
r112 57 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r113 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r114 54 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.825 $Y=0 $X2=4.99
+ $Y2=0
r115 54 56 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.825 $Y=0
+ $X2=4.56 $Y2=0
r116 52 53 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r117 49 53 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=3.6
+ $Y2=0
r118 48 52 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.6
+ $Y2=0
r119 48 49 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r120 45 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r121 45 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r122 43 63 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.685 $Y=0
+ $X2=6.48 $Y2=0
r123 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.685 $Y=0 $X2=6.85
+ $Y2=0
r124 42 67 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=7.015 $Y=0
+ $X2=7.44 $Y2=0
r125 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.015 $Y=0 $X2=6.85
+ $Y2=0
r126 40 60 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=0
+ $X2=5.52 $Y2=0
r127 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=0 $X2=5.85
+ $Y2=0
r128 39 63 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=6.015 $Y=0
+ $X2=6.48 $Y2=0
r129 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.015 $Y=0 $X2=5.85
+ $Y2=0
r130 37 52 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=3.6
+ $Y2=0
r131 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=3.9
+ $Y2=0
r132 36 56 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=4.065 $Y=0
+ $X2=4.56 $Y2=0
r133 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.065 $Y=0 $X2=3.9
+ $Y2=0
r134 32 73 3.09464 $w=3.3e-07 $l=1.15521e-07 $layer=LI1_cond $X=7.85 $Y=0.085
+ $X2=7.922 $Y2=0
r135 32 34 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=7.85 $Y=0.085
+ $X2=7.85 $Y2=0.65
r136 28 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.85 $Y=0.085
+ $X2=6.85 $Y2=0
r137 28 30 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=6.85 $Y=0.085
+ $X2=6.85 $Y2=0.65
r138 24 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.85 $Y=0.085
+ $X2=5.85 $Y2=0
r139 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.85 $Y=0.085
+ $X2=5.85 $Y2=0.515
r140 20 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=0.085
+ $X2=4.99 $Y2=0
r141 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.99 $Y=0.085
+ $X2=4.99 $Y2=0.515
r142 16 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.9 $Y=0.085 $X2=3.9
+ $Y2=0
r143 16 18 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=3.9 $Y=0.085
+ $X2=3.9 $Y2=0.73
r144 5 34 182 $w=1.7e-07 $l=3.70405e-07 $layer=licon1_NDIFF $count=1 $X=7.64
+ $Y=0.37 $X2=7.85 $Y2=0.65
r145 4 30 182 $w=1.7e-07 $l=3.70405e-07 $layer=licon1_NDIFF $count=1 $X=6.64
+ $Y=0.37 $X2=6.85 $Y2=0.65
r146 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.71
+ $Y=0.37 $X2=5.85 $Y2=0.515
r147 2 22 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.845
+ $Y=0.37 $X2=4.99 $Y2=0.515
r148 1 18 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=3.76
+ $Y=0.54 $X2=3.9 $Y2=0.73
.ends

