* File: sky130_fd_sc_ls__or4_2.spice
* Created: Wed Sep  2 11:25:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__or4_2.pex.spice"
.subckt sky130_fd_sc_ls__or4_2  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1004 N_A_85_392#_M1004_d N_D_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.284075 PD=0.92 PS=2.19 NRD=0 NRS=21.552 M=1 R=4.26667
+ SA=75000.4 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1007_d N_C_M1007_g N_A_85_392#_M1004_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1943 AS=0.0896 PD=1.255 PS=0.92 NRD=29.052 NRS=0 M=1 R=4.26667 SA=75000.8
+ SB=75002.5 A=0.096 P=1.58 MULT=1
MM1001 N_A_85_392#_M1001_d N_B_M1001_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1943 PD=0.92 PS=1.255 NRD=0 NRS=29.052 M=1 R=4.26667 SA=75001.5
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_A_M1006_g N_A_85_392#_M1001_d VNB NSHORT L=0.15 W=0.64
+ AD=0.16742 AS=0.0896 PD=1.17333 PS=0.92 NRD=24.372 NRS=0 M=1 R=4.26667
+ SA=75002 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1002 N_X_M1002_d N_A_85_392#_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.19358 PD=1.02 PS=1.35667 NRD=0 NRS=18.648 M=1 R=4.93333
+ SA=75002.3 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1008 N_X_M1002_d N_A_85_392#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 A_174_392# N_D_M1000_g N_A_85_392#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1011 A_258_392# N_C_M1011_g A_174_392# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=15.7403 NRS=15.7403 M=1 R=6.66667 SA=75000.6
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1009 A_342_392# N_B_M1009_g A_258_392# VPB PHIGHVT L=0.15 W=1 AD=0.215
+ AS=0.135 PD=1.43 PS=1.27 NRD=31.5003 NRS=15.7403 M=1 R=6.66667 SA=75001.1
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g A_342_392# VPB PHIGHVT L=0.15 W=1 AD=0.224717
+ AS=0.215 PD=1.46698 PS=1.43 NRD=18.715 NRS=31.5003 M=1 R=6.66667 SA=75001.6
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1005_d N_A_85_392#_M1005_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.251683 PD=1.42 PS=1.64302 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1010 N_X_M1005_d N_A_85_392#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.5 SB=75000.3 A=0.168 P=2.54 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ls__or4_2.pxi.spice"
*
.ends
*
*
