# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__o2bb2a_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__o2bb2a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.415000 1.350000 4.745000 1.780000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.845000 1.350000 4.195000 1.780000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.260000 1.115000 1.770000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.470000 1.450000 2.275000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.311300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.255000 0.350000 5.585000 0.810000 ;
        RECT 5.255000 0.810000 6.585000 1.050000 ;
        RECT 5.255000 1.720000 6.585000 1.890000 ;
        RECT 5.255000 1.890000 5.585000 2.980000 ;
        RECT 6.255000 0.350000 6.585000 0.810000 ;
        RECT 6.255000 1.050000 6.585000 1.720000 ;
        RECT 6.255000 1.890000 6.585000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.200000 0.085000 ;
        RECT 0.615000  0.085000 0.945000 0.750000 ;
        RECT 1.615000  0.085000 1.945000 0.610000 ;
        RECT 4.540000  0.085000 5.080000 0.780000 ;
        RECT 5.755000  0.085000 6.085000 0.640000 ;
        RECT 6.755000  0.085000 7.085000 1.130000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.200000 3.415000 ;
        RECT 0.715000 2.290000 0.885000 3.245000 ;
        RECT 2.545000 2.320000 2.875000 3.245000 ;
        RECT 3.600000 2.790000 3.930000 3.245000 ;
        RECT 4.670000 2.790000 5.000000 3.245000 ;
        RECT 5.755000 2.060000 6.085000 3.245000 ;
        RECT 6.755000 1.820000 7.085000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.350000 0.445000 0.920000 ;
      RECT 0.115000 0.920000 3.335000 1.090000 ;
      RECT 0.185000 1.940000 0.515000 1.950000 ;
      RECT 0.185000 1.950000 1.415000 2.120000 ;
      RECT 0.185000 2.120000 0.515000 2.980000 ;
      RECT 1.085000 2.120000 1.415000 2.905000 ;
      RECT 1.085000 2.905000 2.315000 3.075000 ;
      RECT 1.115000 0.350000 1.445000 0.780000 ;
      RECT 1.115000 0.780000 3.335000 0.920000 ;
      RECT 1.615000 1.950000 3.335000 2.120000 ;
      RECT 1.615000 2.120000 1.785000 2.735000 ;
      RECT 1.985000 2.290000 2.315000 2.905000 ;
      RECT 2.490000 1.300000 3.675000 1.630000 ;
      RECT 2.505000 0.255000 4.370000 0.425000 ;
      RECT 2.505000 0.425000 2.835000 0.610000 ;
      RECT 2.995000 1.820000 3.335000 1.950000 ;
      RECT 2.995000 2.120000 3.335000 2.150000 ;
      RECT 3.005000 0.595000 3.335000 0.780000 ;
      RECT 3.165000 2.150000 3.335000 2.450000 ;
      RECT 3.165000 2.450000 5.085000 2.620000 ;
      RECT 3.505000 0.960000 4.030000 1.130000 ;
      RECT 3.505000 1.130000 3.675000 1.300000 ;
      RECT 3.505000 1.630000 3.675000 1.950000 ;
      RECT 3.505000 1.950000 4.465000 2.280000 ;
      RECT 3.700000 0.635000 4.030000 0.960000 ;
      RECT 4.200000 0.425000 4.370000 0.950000 ;
      RECT 4.200000 0.950000 5.085000 1.120000 ;
      RECT 4.915000 1.120000 5.085000 1.220000 ;
      RECT 4.915000 1.220000 6.065000 1.550000 ;
      RECT 4.915000 1.550000 5.085000 2.450000 ;
  END
END sky130_fd_sc_ls__o2bb2a_4
