* NGSPICE file created from sky130_fd_sc_ls__or2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__or2b_2 A B_N VGND VNB VPB VPWR X
M1000 VPWR a_187_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=8.614e+11p pd=6.09e+06u as=5.768e+11p ps=3.27e+06u
M1001 VGND B_N a_27_368# VNB nshort w=550000u l=150000u
+  ad=9.5555e+11p pd=7.08e+06u as=1.5675e+11p ps=1.67e+06u
M1002 a_187_48# A VGND VNB nshort w=640000u l=150000u
+  ad=2.208e+11p pd=1.97e+06u as=0p ps=0u
M1003 X a_187_48# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1004 VGND a_187_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_27_368# a_187_48# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR B_N a_27_368# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1007 a_187_48# a_27_368# a_470_368# VPB phighvt w=1e+06u l=150000u
+  ad=4.15e+11p pd=2.83e+06u as=2.7e+11p ps=2.54e+06u
M1008 X a_187_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_470_368# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

