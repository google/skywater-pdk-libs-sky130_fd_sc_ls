* NGSPICE file created from sky130_fd_sc_ls__o311ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 a_670_74# B1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=5.18e+11p pd=4.36e+06u as=1.1174e+12p ps=1.042e+07u
M1001 VPWR B1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=1.0192e+12p pd=8.54e+06u as=1.3328e+12p ps=1.134e+07u
M1002 VGND A3 a_27_74# VNB nshort w=740000u l=150000u
+  ad=6.956e+11p pd=6.32e+06u as=0p ps=0u
M1003 a_28_368# A1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=1.0416e+12p pd=8.58e+06u as=0p ps=0u
M1004 Y B1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y C1 a_670_74# VNB nshort w=740000u l=150000u
+  ad=4.218e+11p pd=4.1e+06u as=0p ps=0u
M1006 a_28_368# A2 a_307_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=7.504e+11p ps=5.82e+06u
M1007 VGND A2 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# A2 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_28_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# B1 a_670_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR C1 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_307_368# A3 Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y C1 VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_307_368# A2 a_28_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_74# A3 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A1 a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y A3 a_307_368# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_74# A1 VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_670_74# C1 Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

