# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__a41oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 1.430000 1.795000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.665000 1.300000 3.715000 1.630000 ;
        RECT 3.005000 1.630000 3.715000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.350000 4.675000 1.780000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.350000 5.635000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.085000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.810100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 0.400000 0.945000 1.010000 ;
        RECT 0.615000 1.010000 1.935000 1.090000 ;
        RECT 0.615000 1.090000 2.275000 1.180000 ;
        RECT 0.615000 1.950000 2.135000 2.120000 ;
        RECT 0.615000 2.120000 0.945000 2.735000 ;
        RECT 1.685000 0.595000 1.935000 1.010000 ;
        RECT 1.685000 1.180000 2.275000 1.260000 ;
        RECT 1.965000 1.260000 2.275000 1.650000 ;
        RECT 1.965000 1.650000 2.135000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.180000 ;
      RECT 0.115000  1.950000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 1.445000 3.075000 ;
      RECT 1.115000  2.290000 2.635000 2.460000 ;
      RECT 1.115000  2.460000 1.445000 2.905000 ;
      RECT 1.175000  0.255000 2.355000 0.425000 ;
      RECT 1.175000  0.425000 1.505000 0.840000 ;
      RECT 1.615000  2.650000 2.135000 3.245000 ;
      RECT 2.105000  0.425000 2.355000 0.750000 ;
      RECT 2.105000  0.750000 3.295000 0.920000 ;
      RECT 2.305000  1.820000 2.635000 1.950000 ;
      RECT 2.305000  1.950000 5.645000 2.120000 ;
      RECT 2.305000  2.120000 2.635000 2.290000 ;
      RECT 2.305000  2.460000 2.635000 2.980000 ;
      RECT 2.535000  0.330000 4.285000 0.580000 ;
      RECT 2.805000  2.290000 3.135000 3.245000 ;
      RECT 2.965000  0.920000 3.295000 1.080000 ;
      RECT 3.305000  2.120000 3.635000 2.980000 ;
      RECT 3.525000  0.850000 4.635000 1.010000 ;
      RECT 3.525000  1.010000 5.645000 1.130000 ;
      RECT 3.805000  2.290000 4.135000 3.245000 ;
      RECT 3.955000  0.580000 4.285000 0.680000 ;
      RECT 4.305000  2.120000 4.670000 3.000000 ;
      RECT 4.465000  0.350000 4.635000 0.850000 ;
      RECT 4.465000  1.130000 5.645000 1.180000 ;
      RECT 4.815000  0.085000 5.145000 0.840000 ;
      RECT 4.840000  2.290000 5.170000 3.245000 ;
      RECT 5.315000  0.350000 5.645000 1.010000 ;
      RECT 5.340000  2.120000 5.645000 3.000000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_ls__a41oi_2
END LIBRARY
