* File: sky130_fd_sc_ls__dfrtp_2.pxi.spice
* Created: Fri Aug 28 13:14:39 2020
* 
x_PM_SKY130_FD_SC_LS__DFRTP_2%D N_D_c_243_n N_D_c_248_n N_D_c_249_n N_D_M1022_g
+ N_D_M1025_g D D D N_D_c_245_n N_D_c_246_n N_D_c_251_n
+ PM_SKY130_FD_SC_LS__DFRTP_2%D
x_PM_SKY130_FD_SC_LS__DFRTP_2%CLK N_CLK_c_278_n N_CLK_M1027_g N_CLK_c_279_n
+ N_CLK_M1015_g CLK PM_SKY130_FD_SC_LS__DFRTP_2%CLK
x_PM_SKY130_FD_SC_LS__DFRTP_2%A_495_390# N_A_495_390#_M1012_d
+ N_A_495_390#_M1004_d N_A_495_390#_c_323_n N_A_495_390#_M1008_g
+ N_A_495_390#_c_343_n N_A_495_390#_c_324_n N_A_495_390#_M1014_g
+ N_A_495_390#_c_326_n N_A_495_390#_M1003_g N_A_495_390#_c_327_n
+ N_A_495_390#_c_328_n N_A_495_390#_c_345_n N_A_495_390#_M1002_g
+ N_A_495_390#_c_329_n N_A_495_390#_c_330_n N_A_495_390#_c_331_n
+ N_A_495_390#_c_375_p N_A_495_390#_c_332_n N_A_495_390#_c_333_n
+ N_A_495_390#_c_334_n N_A_495_390#_c_347_n N_A_495_390#_c_335_n
+ N_A_495_390#_c_336_n N_A_495_390#_c_337_n N_A_495_390#_c_338_n
+ N_A_495_390#_c_339_n N_A_495_390#_c_340_n
+ PM_SKY130_FD_SC_LS__DFRTP_2%A_495_390#
x_PM_SKY130_FD_SC_LS__DFRTP_2%A_839_359# N_A_839_359#_M1020_d
+ N_A_839_359#_M1028_d N_A_839_359#_c_521_n N_A_839_359#_M1010_g
+ N_A_839_359#_M1006_g N_A_839_359#_c_517_n N_A_839_359#_c_518_n
+ N_A_839_359#_c_539_n N_A_839_359#_c_542_n N_A_839_359#_c_524_n
+ N_A_839_359#_c_519_n N_A_839_359#_c_520_n
+ PM_SKY130_FD_SC_LS__DFRTP_2%A_839_359#
x_PM_SKY130_FD_SC_LS__DFRTP_2%RESET_B N_RESET_B_M1009_g N_RESET_B_c_604_n
+ N_RESET_B_c_614_n N_RESET_B_M1023_g N_RESET_B_c_605_n N_RESET_B_c_606_n
+ N_RESET_B_M1001_g N_RESET_B_c_608_n N_RESET_B_c_616_n N_RESET_B_M1007_g
+ N_RESET_B_c_617_n N_RESET_B_M1000_g N_RESET_B_M1017_g N_RESET_B_c_619_n
+ N_RESET_B_c_610_n N_RESET_B_c_620_n N_RESET_B_c_621_n N_RESET_B_c_622_n
+ N_RESET_B_c_623_n N_RESET_B_c_624_n N_RESET_B_c_625_n RESET_B
+ N_RESET_B_c_611_n N_RESET_B_c_612_n N_RESET_B_c_627_n N_RESET_B_c_628_n
+ PM_SKY130_FD_SC_LS__DFRTP_2%RESET_B
x_PM_SKY130_FD_SC_LS__DFRTP_2%A_697_463# N_A_697_463#_M1016_d
+ N_A_697_463#_M1008_d N_A_697_463#_M1007_d N_A_697_463#_M1020_g
+ N_A_697_463#_c_814_n N_A_697_463#_M1028_g N_A_697_463#_c_815_n
+ N_A_697_463#_c_822_n N_A_697_463#_c_847_n N_A_697_463#_c_823_n
+ N_A_697_463#_c_816_n N_A_697_463#_c_817_n N_A_697_463#_c_825_n
+ N_A_697_463#_c_818_n N_A_697_463#_c_826_n N_A_697_463#_c_819_n
+ N_A_697_463#_c_864_n PM_SKY130_FD_SC_LS__DFRTP_2%A_697_463#
x_PM_SKY130_FD_SC_LS__DFRTP_2%A_309_390# N_A_309_390#_M1015_s
+ N_A_309_390#_M1027_s N_A_309_390#_c_949_n N_A_309_390#_M1004_g
+ N_A_309_390#_c_939_n N_A_309_390#_M1012_g N_A_309_390#_c_950_n
+ N_A_309_390#_c_951_n N_A_309_390#_c_952_n N_A_309_390#_c_940_n
+ N_A_309_390#_c_941_n N_A_309_390#_c_942_n N_A_309_390#_M1016_g
+ N_A_309_390#_M1011_g N_A_309_390#_c_955_n N_A_309_390#_M1013_g
+ N_A_309_390#_c_943_n N_A_309_390#_c_958_n N_A_309_390#_M1031_g
+ N_A_309_390#_c_959_n N_A_309_390#_c_960_n N_A_309_390#_c_945_n
+ N_A_309_390#_c_946_n N_A_309_390#_c_975_n N_A_309_390#_c_947_n
+ N_A_309_390#_c_948_n N_A_309_390#_c_962_n
+ PM_SKY130_FD_SC_LS__DFRTP_2%A_309_390#
x_PM_SKY130_FD_SC_LS__DFRTP_2%A_1525_212# N_A_1525_212#_M1018_d
+ N_A_1525_212#_M1000_d N_A_1525_212#_M1005_g N_A_1525_212#_c_1126_n
+ N_A_1525_212#_c_1127_n N_A_1525_212#_c_1128_n N_A_1525_212#_M1026_g
+ N_A_1525_212#_c_1118_n N_A_1525_212#_c_1119_n N_A_1525_212#_c_1130_n
+ N_A_1525_212#_c_1120_n N_A_1525_212#_c_1131_n N_A_1525_212#_c_1132_n
+ N_A_1525_212#_c_1133_n N_A_1525_212#_c_1121_n N_A_1525_212#_c_1122_n
+ N_A_1525_212#_c_1123_n N_A_1525_212#_c_1124_n N_A_1525_212#_c_1125_n
+ PM_SKY130_FD_SC_LS__DFRTP_2%A_1525_212#
x_PM_SKY130_FD_SC_LS__DFRTP_2%A_1271_74# N_A_1271_74#_M1003_d
+ N_A_1271_74#_M1013_d N_A_1271_74#_M1018_g N_A_1271_74#_c_1245_n
+ N_A_1271_74#_c_1246_n N_A_1271_74#_M1033_g N_A_1271_74#_c_1236_n
+ N_A_1271_74#_c_1237_n N_A_1271_74#_c_1249_n N_A_1271_74#_c_1250_n
+ N_A_1271_74#_M1024_g N_A_1271_74#_M1019_g N_A_1271_74#_c_1239_n
+ N_A_1271_74#_c_1259_n N_A_1271_74#_c_1240_n N_A_1271_74#_c_1252_n
+ N_A_1271_74#_c_1241_n N_A_1271_74#_c_1273_n N_A_1271_74#_c_1367_p
+ N_A_1271_74#_c_1253_n N_A_1271_74#_c_1242_n N_A_1271_74#_c_1243_n
+ N_A_1271_74#_c_1244_n N_A_1271_74#_c_1257_n
+ PM_SKY130_FD_SC_LS__DFRTP_2%A_1271_74#
x_PM_SKY130_FD_SC_LS__DFRTP_2%A_1921_409# N_A_1921_409#_M1019_d
+ N_A_1921_409#_M1024_d N_A_1921_409#_c_1383_n N_A_1921_409#_c_1384_n
+ N_A_1921_409#_c_1396_n N_A_1921_409#_M1021_g N_A_1921_409#_M1029_g
+ N_A_1921_409#_c_1386_n N_A_1921_409#_c_1387_n N_A_1921_409#_c_1398_n
+ N_A_1921_409#_M1030_g N_A_1921_409#_M1032_g N_A_1921_409#_c_1389_n
+ N_A_1921_409#_c_1390_n N_A_1921_409#_c_1399_n N_A_1921_409#_c_1391_n
+ N_A_1921_409#_c_1392_n N_A_1921_409#_c_1393_n N_A_1921_409#_c_1394_n
+ PM_SKY130_FD_SC_LS__DFRTP_2%A_1921_409#
x_PM_SKY130_FD_SC_LS__DFRTP_2%VPWR N_VPWR_M1022_s N_VPWR_M1023_d N_VPWR_M1027_d
+ N_VPWR_M1010_d N_VPWR_M1028_s N_VPWR_M1026_d N_VPWR_M1033_d N_VPWR_M1021_s
+ N_VPWR_M1030_s N_VPWR_c_1456_n N_VPWR_c_1457_n N_VPWR_c_1458_n N_VPWR_c_1459_n
+ N_VPWR_c_1460_n N_VPWR_c_1461_n N_VPWR_c_1462_n N_VPWR_c_1463_n
+ N_VPWR_c_1464_n N_VPWR_c_1465_n N_VPWR_c_1466_n N_VPWR_c_1467_n
+ N_VPWR_c_1468_n N_VPWR_c_1469_n VPWR N_VPWR_c_1470_n N_VPWR_c_1471_n
+ N_VPWR_c_1472_n N_VPWR_c_1473_n N_VPWR_c_1474_n N_VPWR_c_1475_n
+ N_VPWR_c_1476_n N_VPWR_c_1477_n N_VPWR_c_1478_n N_VPWR_c_1479_n
+ N_VPWR_c_1480_n N_VPWR_c_1481_n N_VPWR_c_1455_n
+ PM_SKY130_FD_SC_LS__DFRTP_2%VPWR
x_PM_SKY130_FD_SC_LS__DFRTP_2%A_30_78# N_A_30_78#_M1025_s N_A_30_78#_M1016_s
+ N_A_30_78#_M1022_d N_A_30_78#_M1008_s N_A_30_78#_c_1614_n N_A_30_78#_c_1621_n
+ N_A_30_78#_c_1615_n N_A_30_78#_c_1623_n N_A_30_78#_c_1624_n
+ N_A_30_78#_c_1616_n N_A_30_78#_c_1625_n N_A_30_78#_c_1617_n
+ N_A_30_78#_c_1618_n N_A_30_78#_c_1627_n N_A_30_78#_c_1628_n
+ N_A_30_78#_c_1619_n N_A_30_78#_c_1620_n PM_SKY130_FD_SC_LS__DFRTP_2%A_30_78#
x_PM_SKY130_FD_SC_LS__DFRTP_2%Q N_Q_M1029_d N_Q_M1021_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LS__DFRTP_2%Q
x_PM_SKY130_FD_SC_LS__DFRTP_2%VGND N_VGND_M1009_d N_VGND_M1015_d N_VGND_M1001_d
+ N_VGND_M1005_d N_VGND_M1019_s N_VGND_M1029_s N_VGND_M1032_s N_VGND_c_1769_n
+ N_VGND_c_1770_n N_VGND_c_1771_n N_VGND_c_1772_n N_VGND_c_1773_n
+ N_VGND_c_1774_n N_VGND_c_1775_n N_VGND_c_1776_n VGND N_VGND_c_1777_n
+ N_VGND_c_1778_n N_VGND_c_1779_n N_VGND_c_1780_n N_VGND_c_1781_n
+ N_VGND_c_1782_n N_VGND_c_1783_n N_VGND_c_1784_n N_VGND_c_1785_n
+ N_VGND_c_1786_n N_VGND_c_1787_n N_VGND_c_1788_n
+ PM_SKY130_FD_SC_LS__DFRTP_2%VGND
cc_1 VNB N_D_c_243_n 0.040598f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.828
cc_2 VNB N_D_M1025_g 0.0286444f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_3 VNB N_D_c_245_n 0.0216261f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_4 VNB N_D_c_246_n 0.0279969f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_5 VNB N_CLK_c_278_n 0.0225612f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.182
cc_6 VNB N_CLK_c_279_n 0.0155569f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_7 VNB CLK 0.00281093f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1
cc_8 VNB N_A_495_390#_c_323_n 0.00226217f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.75
cc_9 VNB N_A_495_390#_c_324_n 0.0146344f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB N_A_495_390#_M1014_g 0.0252137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_495_390#_c_326_n 0.0178063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_495_390#_c_327_n 0.0205353f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_13 VNB N_A_495_390#_c_328_n 0.010064f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1
cc_14 VNB N_A_495_390#_c_329_n 0.0082862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_495_390#_c_330_n 0.0342757f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.295
cc_16 VNB N_A_495_390#_c_331_n 0.00299032f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.665
cc_17 VNB N_A_495_390#_c_332_n 0.0145916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_495_390#_c_333_n 0.00228045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_495_390#_c_334_n 0.0036821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_495_390#_c_335_n 0.00197952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_495_390#_c_336_n 0.00264192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_495_390#_c_337_n 0.0129363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_495_390#_c_338_n 0.00711318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_495_390#_c_339_n 0.0318573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_495_390#_c_340_n 0.00728799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_839_359#_M1006_g 0.0276542f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_27 VNB N_A_839_359#_c_517_n 0.00256007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_839_359#_c_518_n 0.0099177f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_29 VNB N_A_839_359#_c_519_n 0.00239189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_839_359#_c_520_n 0.00880031f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.845
cc_31 VNB N_RESET_B_M1009_g 0.0210204f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.375
cc_32 VNB N_RESET_B_c_604_n 0.0235199f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.75
cc_33 VNB N_RESET_B_c_605_n 0.280594f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_34 VNB N_RESET_B_c_606_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_35 VNB N_RESET_B_M1001_g 0.0342254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_RESET_B_c_608_n 0.0104399f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_37 VNB N_RESET_B_M1017_g 0.0519208f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.295
cc_38 VNB N_RESET_B_c_610_n 0.0156921f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=2.035
cc_39 VNB N_RESET_B_c_611_n 0.0389069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_RESET_B_c_612_n 0.00329735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_697_463#_M1020_g 0.0236184f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_42 VNB N_A_697_463#_c_814_n 0.0170235f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_43 VNB N_A_697_463#_c_815_n 0.026897f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.165
cc_44 VNB N_A_697_463#_c_816_n 0.00249866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_697_463#_c_817_n 0.00408962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_697_463#_c_818_n 0.00211346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_697_463#_c_819_n 0.00233475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_309_390#_c_939_n 0.0146915f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_49 VNB N_A_309_390#_c_940_n 0.0333154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_309_390#_c_941_n 0.0608621f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.165
cc_51 VNB N_A_309_390#_c_942_n 0.0172403f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_52 VNB N_A_309_390#_c_943_n 0.0126064f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.845
cc_53 VNB N_A_309_390#_M1031_g 0.0521291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_309_390#_c_945_n 0.013578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_309_390#_c_946_n 0.00805872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_309_390#_c_947_n 9.72279e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_309_390#_c_948_n 0.00351963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1525_212#_M1005_g 0.0235036f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_59 VNB N_A_1525_212#_c_1118_n 0.013872f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.165
cc_60 VNB N_A_1525_212#_c_1119_n 0.0150411f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_61 VNB N_A_1525_212#_c_1120_n 0.0124228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1525_212#_c_1121_n 0.0141072f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=2.035
cc_63 VNB N_A_1525_212#_c_1122_n 0.00326635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1525_212#_c_1123_n 0.00415979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1525_212#_c_1124_n 0.031534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1525_212#_c_1125_n 0.00288865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1271_74#_M1018_g 0.0561848f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_68 VNB N_A_1271_74#_c_1236_n 0.0155616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1271_74#_c_1237_n 0.0127478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1271_74#_M1019_g 0.0397312f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=2.01
cc_71 VNB N_A_1271_74#_c_1239_n 0.00459979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1271_74#_c_1240_n 0.00477322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1271_74#_c_1241_n 0.00415183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1271_74#_c_1242_n 0.00523477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1271_74#_c_1243_n 0.00751489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1271_74#_c_1244_n 0.00236307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1921_409#_c_1383_n 0.0140421f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=2.75
cc_78 VNB N_A_1921_409#_c_1384_n 0.0102109f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_79 VNB N_A_1921_409#_M1029_g 0.0229651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1921_409#_c_1386_n 0.00938445f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.165
cc_81 VNB N_A_1921_409#_c_1387_n 0.0167069f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1
cc_82 VNB N_A_1921_409#_M1032_g 0.0260342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1921_409#_c_1389_n 0.00591123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1921_409#_c_1390_n 0.0111562f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=1.665
cc_85 VNB N_A_1921_409#_c_1391_n 0.0124224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1921_409#_c_1392_n 0.00109385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1921_409#_c_1393_n 0.00157695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1921_409#_c_1394_n 0.0465967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VPWR_c_1455_n 0.48212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_30_78#_c_1614_n 0.00271393f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_91 VNB N_A_30_78#_c_1615_n 0.00538705f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_92 VNB N_A_30_78#_c_1616_n 9.52573e-19 $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.165
cc_93 VNB N_A_30_78#_c_1617_n 0.0032682f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.665
cc_94 VNB N_A_30_78#_c_1618_n 0.0223919f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.845
cc_95 VNB N_A_30_78#_c_1619_n 0.00159616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_30_78#_c_1620_n 0.00571698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB Q 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.75
cc_98 VNB N_VGND_c_1769_n 0.00871111f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_99 VNB N_VGND_c_1770_n 0.0203532f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.165
cc_100 VNB N_VGND_c_1771_n 0.0116406f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.665
cc_101 VNB N_VGND_c_1772_n 0.00612754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1773_n 0.0164559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1774_n 0.0191664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1775_n 0.0105185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1776_n 0.0507342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1777_n 0.0290143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1778_n 0.0773321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1779_n 0.0578377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1780_n 0.0306389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1781_n 0.0209223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1782_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1783_n 0.00372873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1784_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1785_n 0.0080786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1786_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1787_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1788_n 0.608208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VPB N_D_c_243_n 0.0142136f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.828
cc_119 VPB N_D_c_248_n 0.0278558f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.375
cc_120 VPB N_D_c_249_n 0.0277349f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.465
cc_121 VPB N_D_c_246_n 0.0227717f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_122 VPB N_D_c_251_n 0.0207699f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_123 VPB N_CLK_c_278_n 0.0127766f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.182
cc_124 VPB N_CLK_M1027_g 0.0221764f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.01
cc_125 VPB CLK 0.00342379f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_126 VPB N_A_495_390#_c_323_n 0.0287832f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_127 VPB N_A_495_390#_M1008_g 0.0287256f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_128 VPB N_A_495_390#_c_343_n 0.0223188f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_495_390#_c_324_n 0.0177812f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_130 VPB N_A_495_390#_c_345_n 0.0194137f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_131 VPB N_A_495_390#_c_334_n 0.006052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_495_390#_c_347_n 0.0479926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_495_390#_c_336_n 0.0103833f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_839_359#_c_521_n 0.0626503f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_135 VPB N_A_839_359#_M1006_g 0.0125375f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_136 VPB N_A_839_359#_c_517_n 0.00243408f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_839_359#_c_524_n 5.83759e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_839_359#_c_520_n 0.00377881f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.845
cc_139 VPB N_RESET_B_c_604_n 0.0208082f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_140 VPB N_RESET_B_c_614_n 0.017748f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_141 VPB N_RESET_B_c_608_n 0.0181282f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_142 VPB N_RESET_B_c_616_n 0.0715955f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_143 VPB N_RESET_B_c_617_n 0.0571202f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_144 VPB N_RESET_B_M1017_g 0.0162636f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.295
cc_145 VPB N_RESET_B_c_619_n 0.0262718f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.665
cc_146 VPB N_RESET_B_c_620_n 0.0192355f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_RESET_B_c_621_n 0.00199327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_RESET_B_c_622_n 0.020195f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_RESET_B_c_623_n 0.00143938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_RESET_B_c_624_n 0.00397837f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_RESET_B_c_625_n 0.0019787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_RESET_B_c_612_n 7.70379e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_RESET_B_c_627_n 0.0332067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_RESET_B_c_628_n 0.00930396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_697_463#_c_814_n 0.0288648f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_156 VPB N_A_697_463#_c_815_n 0.0122975f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.165
cc_157 VPB N_A_697_463#_c_822_n 0.00334632f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_158 VPB N_A_697_463#_c_823_n 0.0117494f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.295
cc_159 VPB N_A_697_463#_c_817_n 0.00331109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_697_463#_c_825_n 0.00255206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_697_463#_c_826_n 0.00208187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_697_463#_c_819_n 0.0067815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_309_390#_c_949_n 0.0155222f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_164 VPB N_A_309_390#_c_950_n 0.0692226f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_165 VPB N_A_309_390#_c_951_n 0.059821f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_309_390#_c_952_n 0.0125215f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_309_390#_c_941_n 0.0236807f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.165
cc_168 VPB N_A_309_390#_M1011_g 0.035005f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_169 VPB N_A_309_390#_c_955_n 0.171666f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.165
cc_170 VPB N_A_309_390#_M1013_g 0.0107276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_309_390#_c_943_n 0.0397359f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.845
cc_172 VPB N_A_309_390#_c_958_n 0.00832634f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=2.035
cc_173 VPB N_A_309_390#_c_959_n 0.00749069f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_309_390#_c_960_n 0.0335383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_309_390#_c_946_n 0.00488299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_309_390#_c_962_n 0.00936754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_1525_212#_c_1126_n 0.00452844f $X=-0.19 $Y=1.66 $X2=0.155
+ $Y2=1.58
cc_178 VPB N_A_1525_212#_c_1127_n 0.0112203f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_179 VPB N_A_1525_212#_c_1128_n 0.0209833f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_1525_212#_c_1118_n 0.0172903f $X=-0.19 $Y=1.66 $X2=0.402
+ $Y2=1.165
cc_181 VPB N_A_1525_212#_c_1130_n 0.0123021f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1
cc_182 VPB N_A_1525_212#_c_1131_n 0.00195592f $X=-0.19 $Y=1.66 $X2=0.31
+ $Y2=1.665
cc_183 VPB N_A_1525_212#_c_1132_n 0.00467452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1525_212#_c_1133_n 0.00234171f $X=-0.19 $Y=1.66 $X2=0.31
+ $Y2=1.845
cc_185 VPB N_A_1525_212#_c_1122_n 0.00587125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1271_74#_c_1245_n 0.0253818f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_187 VPB N_A_1271_74#_c_1246_n 0.0240491f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_188 VPB N_A_1271_74#_c_1236_n 0.00814854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_1271_74#_c_1237_n 0.0260612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1271_74#_c_1249_n 0.010774f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_191 VPB N_A_1271_74#_c_1250_n 0.0240694f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_192 VPB N_A_1271_74#_c_1239_n 0.00430295f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_1271_74#_c_1252_n 0.00135315f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1271_74#_c_1253_n 0.0127664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_1271_74#_c_1242_n 0.0140489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_1271_74#_c_1243_n 4.13852e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1271_74#_c_1244_n 4.64263e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_1271_74#_c_1257_n 0.00154868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1921_409#_c_1384_n 8.65682e-19 $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_200 VPB N_A_1921_409#_c_1396_n 0.023821f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_1921_409#_c_1387_n 0.00111912f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1
cc_202 VPB N_A_1921_409#_c_1398_n 0.0258791f $X=-0.19 $Y=1.66 $X2=0.402
+ $Y2=1.845
cc_203 VPB N_A_1921_409#_c_1399_n 0.0117303f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=2.035
cc_204 VPB N_A_1921_409#_c_1392_n 0.00710574f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1456_n 0.0116916f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.295
cc_206 VPB N_VPWR_c_1457_n 0.0302543f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.665
cc_207 VPB N_VPWR_c_1458_n 0.00856728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1459_n 0.00620939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1460_n 0.0139706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1461_n 0.0203378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1462_n 0.0243365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1463_n 0.0152192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1464_n 0.0163857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1465_n 0.0261554f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1466_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1467_n 0.0638885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1468_n 0.0275707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1469_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1470_n 0.0163062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1471_n 0.0173513f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1472_n 0.0583126f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1473_n 0.0531608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1474_n 0.0209549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1475_n 0.0188539f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1476_n 0.00615076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1477_n 0.00620759f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1478_n 0.00436844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1479_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1480_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1481_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1455_n 0.116787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_30_78#_c_1621_n 0.00206793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_30_78#_c_1615_n 0.00603977f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_234 VPB N_A_30_78#_c_1623_n 0.00983678f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1
cc_235 VPB N_A_30_78#_c_1624_n 0.00170215f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_236 VPB N_A_30_78#_c_1625_n 0.00157227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_30_78#_c_1617_n 0.00724521f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.665
cc_238 VPB N_A_30_78#_c_1627_n 0.00361565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_30_78#_c_1628_n 0.00604038f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB Q 0.00331763f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_241 N_D_M1025_g N_RESET_B_M1009_g 0.0245857f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_242 N_D_c_246_n N_RESET_B_M1009_g 9.4205e-19 $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_243 N_D_c_243_n N_RESET_B_c_604_n 0.0245857f $X=0.402 $Y=1.828 $X2=0 $Y2=0
cc_244 N_D_c_248_n N_RESET_B_c_614_n 0.00630178f $X=0.495 $Y=2.375 $X2=0 $Y2=0
cc_245 N_D_c_249_n N_RESET_B_c_619_n 0.0148339f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_246 N_D_c_245_n N_RESET_B_c_611_n 0.0245857f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_247 N_D_c_251_n N_RESET_B_c_627_n 0.0245857f $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_248 N_D_c_249_n N_VPWR_c_1457_n 0.0113744f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_249 N_D_c_246_n N_VPWR_c_1457_n 0.0172326f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_250 N_D_c_251_n N_VPWR_c_1457_n 9.92489e-19 $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_251 N_D_c_249_n N_VPWR_c_1458_n 3.88309e-19 $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_252 N_D_c_249_n N_VPWR_c_1470_n 0.00413917f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_253 N_D_c_249_n N_VPWR_c_1455_n 0.00855638f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_254 N_D_M1025_g N_A_30_78#_c_1614_n 0.0114706f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_255 N_D_c_246_n N_A_30_78#_c_1614_n 0.00258996f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_256 N_D_c_249_n N_A_30_78#_c_1621_n 0.00129623f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_257 N_D_M1025_g N_A_30_78#_c_1615_n 0.0154787f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_258 N_D_c_246_n N_A_30_78#_c_1615_n 0.088088f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_259 N_D_M1025_g N_A_30_78#_c_1618_n 0.00795006f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_260 N_D_c_245_n N_A_30_78#_c_1618_n 0.00161806f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_261 N_D_c_246_n N_A_30_78#_c_1618_n 0.0286676f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_262 N_D_c_248_n N_A_30_78#_c_1627_n 0.00414406f $X=0.495 $Y=2.375 $X2=0 $Y2=0
cc_263 N_D_c_249_n N_A_30_78#_c_1627_n 0.00223635f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_264 N_D_M1025_g N_VGND_c_1769_n 0.00200176f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_265 N_D_M1025_g N_VGND_c_1777_n 0.00429844f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_266 N_D_M1025_g N_VGND_c_1788_n 0.00539454f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_267 N_CLK_c_278_n N_RESET_B_c_604_n 0.00760467f $X=1.905 $Y=1.775 $X2=0 $Y2=0
cc_268 N_CLK_M1027_g N_RESET_B_c_604_n 0.00576443f $X=1.905 $Y=2.45 $X2=0 $Y2=0
cc_269 N_CLK_c_279_n N_RESET_B_c_605_n 0.0104164f $X=1.985 $Y=1.435 $X2=0 $Y2=0
cc_270 N_CLK_c_278_n N_RESET_B_c_620_n 0.00178944f $X=1.905 $Y=1.775 $X2=0 $Y2=0
cc_271 N_CLK_M1027_g N_RESET_B_c_620_n 0.00329773f $X=1.905 $Y=2.45 $X2=0 $Y2=0
cc_272 CLK N_RESET_B_c_620_n 0.0124899f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_273 N_CLK_c_279_n N_RESET_B_c_611_n 0.00417243f $X=1.985 $Y=1.435 $X2=0 $Y2=0
cc_274 CLK N_A_309_390#_M1015_s 7.75403e-19 $X=2.075 $Y=1.58 $X2=-0.19
+ $Y2=-0.245
cc_275 N_CLK_c_279_n N_A_309_390#_c_939_n 0.024168f $X=1.985 $Y=1.435 $X2=0
+ $Y2=0
cc_276 CLK N_A_309_390#_c_939_n 3.55187e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_277 N_CLK_c_278_n N_A_309_390#_c_941_n 0.0219382f $X=1.905 $Y=1.775 $X2=0
+ $Y2=0
cc_278 N_CLK_M1027_g N_A_309_390#_c_941_n 0.0412212f $X=1.905 $Y=2.45 $X2=0
+ $Y2=0
cc_279 N_CLK_c_279_n N_A_309_390#_c_941_n 0.00112132f $X=1.985 $Y=1.435 $X2=0
+ $Y2=0
cc_280 CLK N_A_309_390#_c_941_n 0.0032861f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_281 N_CLK_c_279_n N_A_309_390#_c_945_n 0.00655396f $X=1.985 $Y=1.435 $X2=0
+ $Y2=0
cc_282 N_CLK_c_278_n N_A_309_390#_c_946_n 0.00291925f $X=1.905 $Y=1.775 $X2=0
+ $Y2=0
cc_283 N_CLK_M1027_g N_A_309_390#_c_946_n 0.00263835f $X=1.905 $Y=2.45 $X2=0
+ $Y2=0
cc_284 N_CLK_c_279_n N_A_309_390#_c_946_n 0.0037005f $X=1.985 $Y=1.435 $X2=0
+ $Y2=0
cc_285 CLK N_A_309_390#_c_946_n 0.034209f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_286 N_CLK_c_278_n N_A_309_390#_c_975_n 2.42596e-19 $X=1.905 $Y=1.775 $X2=0
+ $Y2=0
cc_287 N_CLK_c_279_n N_A_309_390#_c_975_n 0.0134676f $X=1.985 $Y=1.435 $X2=0
+ $Y2=0
cc_288 CLK N_A_309_390#_c_975_n 0.0234841f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_289 N_CLK_c_278_n N_A_309_390#_c_947_n 2.6382e-19 $X=1.905 $Y=1.775 $X2=0
+ $Y2=0
cc_290 CLK N_A_309_390#_c_947_n 0.0316459f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_291 N_CLK_c_278_n N_A_309_390#_c_948_n 0.00101066f $X=1.905 $Y=1.775 $X2=0
+ $Y2=0
cc_292 CLK N_A_309_390#_c_948_n 0.00504033f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_293 N_CLK_c_278_n N_A_309_390#_c_962_n 0.00146257f $X=1.905 $Y=1.775 $X2=0
+ $Y2=0
cc_294 N_CLK_M1027_g N_A_309_390#_c_962_n 0.0062774f $X=1.905 $Y=2.45 $X2=0
+ $Y2=0
cc_295 CLK N_A_309_390#_c_962_n 0.00496992f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_296 N_CLK_M1027_g N_VPWR_c_1458_n 0.00591251f $X=1.905 $Y=2.45 $X2=0 $Y2=0
cc_297 N_CLK_M1027_g N_VPWR_c_1459_n 0.00956982f $X=1.905 $Y=2.45 $X2=0 $Y2=0
cc_298 N_CLK_M1027_g N_VPWR_c_1471_n 0.00374369f $X=1.905 $Y=2.45 $X2=0 $Y2=0
cc_299 N_CLK_M1027_g N_VPWR_c_1455_n 0.00455844f $X=1.905 $Y=2.45 $X2=0 $Y2=0
cc_300 N_CLK_c_278_n N_A_30_78#_c_1623_n 0.00151595f $X=1.905 $Y=1.775 $X2=0
+ $Y2=0
cc_301 N_CLK_M1027_g N_A_30_78#_c_1623_n 0.0195312f $X=1.905 $Y=2.45 $X2=0 $Y2=0
cc_302 CLK N_A_30_78#_c_1623_n 0.00499685f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_303 CLK N_VGND_M1015_d 0.00186195f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_304 N_CLK_c_279_n N_VGND_c_1771_n 0.00254438f $X=1.985 $Y=1.435 $X2=0 $Y2=0
cc_305 N_CLK_c_279_n N_VGND_c_1788_n 9.39239e-19 $X=1.985 $Y=1.435 $X2=0 $Y2=0
cc_306 N_A_495_390#_c_332_n N_A_839_359#_M1020_d 0.00224297f $X=7.285 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_307 N_A_495_390#_c_323_n N_A_839_359#_c_521_n 0.0019113f $X=3.41 $Y=1.99
+ $X2=0 $Y2=0
cc_308 N_A_495_390#_M1008_g N_A_839_359#_c_521_n 0.00233668f $X=3.41 $Y=2.525
+ $X2=0 $Y2=0
cc_309 N_A_495_390#_c_324_n N_A_839_359#_c_521_n 5.89221e-19 $X=4.04 $Y=1.405
+ $X2=0 $Y2=0
cc_310 N_A_495_390#_c_324_n N_A_839_359#_M1006_g 0.00718049f $X=4.04 $Y=1.405
+ $X2=0 $Y2=0
cc_311 N_A_495_390#_M1014_g N_A_839_359#_M1006_g 0.0501476f $X=4.04 $Y=0.9 $X2=0
+ $Y2=0
cc_312 N_A_495_390#_c_331_n N_A_839_359#_M1006_g 0.00327805f $X=5.515 $Y=0.7
+ $X2=0 $Y2=0
cc_313 N_A_495_390#_c_338_n N_A_839_359#_M1006_g 0.00736621f $X=4.39 $Y=0.415
+ $X2=0 $Y2=0
cc_314 N_A_495_390#_c_324_n N_A_839_359#_c_517_n 6.07387e-19 $X=4.04 $Y=1.405
+ $X2=0 $Y2=0
cc_315 N_A_495_390#_M1014_g N_A_839_359#_c_517_n 0.00230405f $X=4.04 $Y=0.9
+ $X2=0 $Y2=0
cc_316 N_A_495_390#_c_331_n N_A_839_359#_c_518_n 0.0748058f $X=5.515 $Y=0.7
+ $X2=0 $Y2=0
cc_317 N_A_495_390#_c_332_n N_A_839_359#_c_518_n 0.00332639f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_318 N_A_495_390#_c_338_n N_A_839_359#_c_518_n 0.00210258f $X=4.39 $Y=0.415
+ $X2=0 $Y2=0
cc_319 N_A_495_390#_M1014_g N_A_839_359#_c_539_n 0.00105317f $X=4.04 $Y=0.9
+ $X2=0 $Y2=0
cc_320 N_A_495_390#_c_330_n N_A_839_359#_c_539_n 0.00107065f $X=4.305 $Y=0.415
+ $X2=0 $Y2=0
cc_321 N_A_495_390#_c_338_n N_A_839_359#_c_539_n 0.00739265f $X=4.39 $Y=0.415
+ $X2=0 $Y2=0
cc_322 N_A_495_390#_c_332_n N_A_839_359#_c_542_n 0.0176299f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_323 N_A_495_390#_c_328_n N_A_839_359#_c_524_n 0.00325656f $X=6.355 $Y=1.27
+ $X2=0 $Y2=0
cc_324 N_A_495_390#_c_326_n N_A_839_359#_c_519_n 4.62933e-19 $X=6.28 $Y=1.195
+ $X2=0 $Y2=0
cc_325 N_A_495_390#_c_326_n N_A_839_359#_c_520_n 0.00207614f $X=6.28 $Y=1.195
+ $X2=0 $Y2=0
cc_326 N_A_495_390#_M1014_g N_RESET_B_c_605_n 0.00526413f $X=4.04 $Y=0.9 $X2=0
+ $Y2=0
cc_327 N_A_495_390#_c_330_n N_RESET_B_c_605_n 0.0234047f $X=4.305 $Y=0.415 $X2=0
+ $Y2=0
cc_328 N_A_495_390#_c_331_n N_RESET_B_c_605_n 0.00226538f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_329 N_A_495_390#_c_337_n N_RESET_B_c_605_n 0.0109684f $X=2.832 $Y=0.415 $X2=0
+ $Y2=0
cc_330 N_A_495_390#_c_338_n N_RESET_B_c_605_n 0.0022188f $X=4.39 $Y=0.415 $X2=0
+ $Y2=0
cc_331 N_A_495_390#_c_331_n N_RESET_B_M1001_g 0.0133177f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_332 N_A_495_390#_c_375_p N_RESET_B_M1001_g 0.00355258f $X=5.6 $Y=0.615 $X2=0
+ $Y2=0
cc_333 N_A_495_390#_c_338_n N_RESET_B_M1001_g 0.00642047f $X=4.39 $Y=0.415 $X2=0
+ $Y2=0
cc_334 N_A_495_390#_M1004_d N_RESET_B_c_620_n 7.7211e-19 $X=2.475 $Y=1.95 $X2=0
+ $Y2=0
cc_335 N_A_495_390#_c_323_n N_RESET_B_c_620_n 0.00317523f $X=3.41 $Y=1.99 $X2=0
+ $Y2=0
cc_336 N_A_495_390#_M1008_g N_RESET_B_c_620_n 0.00362964f $X=3.41 $Y=2.525 $X2=0
+ $Y2=0
cc_337 N_A_495_390#_c_343_n N_RESET_B_c_620_n 0.00497139f $X=3.825 $Y=1.73 $X2=0
+ $Y2=0
cc_338 N_A_495_390#_c_324_n N_RESET_B_c_620_n 2.66122e-19 $X=4.04 $Y=1.405 $X2=0
+ $Y2=0
cc_339 N_A_495_390#_c_336_n N_RESET_B_c_620_n 0.0501768f $X=2.967 $Y=1.95 $X2=0
+ $Y2=0
cc_340 N_A_495_390#_c_334_n N_RESET_B_c_622_n 0.0218177f $X=7.12 $Y=2.14 $X2=0
+ $Y2=0
cc_341 N_A_495_390#_c_347_n N_RESET_B_c_622_n 0.00331406f $X=7.12 $Y=2.14 $X2=0
+ $Y2=0
cc_342 N_A_495_390#_c_326_n N_A_697_463#_M1020_g 0.0126968f $X=6.28 $Y=1.195
+ $X2=0 $Y2=0
cc_343 N_A_495_390#_c_332_n N_A_697_463#_M1020_g 0.0119914f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_344 N_A_495_390#_c_328_n N_A_697_463#_c_814_n 0.0126968f $X=6.355 $Y=1.27
+ $X2=0 $Y2=0
cc_345 N_A_495_390#_M1008_g N_A_697_463#_c_822_n 4.14464e-19 $X=3.41 $Y=2.525
+ $X2=0 $Y2=0
cc_346 N_A_495_390#_c_343_n N_A_697_463#_c_818_n 0.00144393f $X=3.825 $Y=1.73
+ $X2=0 $Y2=0
cc_347 N_A_495_390#_c_324_n N_A_697_463#_c_818_n 0.00334951f $X=4.04 $Y=1.405
+ $X2=0 $Y2=0
cc_348 N_A_495_390#_M1014_g N_A_697_463#_c_818_n 0.0100409f $X=4.04 $Y=0.9 $X2=0
+ $Y2=0
cc_349 N_A_495_390#_c_330_n N_A_697_463#_c_818_n 0.0333997f $X=4.305 $Y=0.415
+ $X2=0 $Y2=0
cc_350 N_A_495_390#_c_338_n N_A_697_463#_c_818_n 0.00455642f $X=4.39 $Y=0.415
+ $X2=0 $Y2=0
cc_351 N_A_495_390#_M1008_g N_A_697_463#_c_819_n 4.15172e-19 $X=3.41 $Y=2.525
+ $X2=0 $Y2=0
cc_352 N_A_495_390#_c_324_n N_A_697_463#_c_819_n 0.0146355f $X=4.04 $Y=1.405
+ $X2=0 $Y2=0
cc_353 N_A_495_390#_M1014_g N_A_697_463#_c_819_n 0.0094578f $X=4.04 $Y=0.9 $X2=0
+ $Y2=0
cc_354 N_A_495_390#_c_336_n N_A_309_390#_c_949_n 0.00183339f $X=2.967 $Y=1.95
+ $X2=0 $Y2=0
cc_355 N_A_495_390#_c_329_n N_A_309_390#_c_939_n 0.0055904f $X=2.967 $Y=1.625
+ $X2=0 $Y2=0
cc_356 N_A_495_390#_c_337_n N_A_309_390#_c_939_n 0.00644381f $X=2.832 $Y=0.415
+ $X2=0 $Y2=0
cc_357 N_A_495_390#_c_323_n N_A_309_390#_c_950_n 0.0215742f $X=3.41 $Y=1.99
+ $X2=0 $Y2=0
cc_358 N_A_495_390#_c_336_n N_A_309_390#_c_950_n 0.0166616f $X=2.967 $Y=1.95
+ $X2=0 $Y2=0
cc_359 N_A_495_390#_M1008_g N_A_309_390#_c_951_n 0.0103507f $X=3.41 $Y=2.525
+ $X2=0 $Y2=0
cc_360 N_A_495_390#_c_323_n N_A_309_390#_c_940_n 0.0169707f $X=3.41 $Y=1.99
+ $X2=0 $Y2=0
cc_361 N_A_495_390#_c_336_n N_A_309_390#_c_940_n 0.00553489f $X=2.967 $Y=1.95
+ $X2=0 $Y2=0
cc_362 N_A_495_390#_c_323_n N_A_309_390#_c_941_n 0.0212328f $X=3.41 $Y=1.99
+ $X2=0 $Y2=0
cc_363 N_A_495_390#_c_329_n N_A_309_390#_c_941_n 0.023801f $X=2.967 $Y=1.625
+ $X2=0 $Y2=0
cc_364 N_A_495_390#_c_336_n N_A_309_390#_c_941_n 0.0178635f $X=2.967 $Y=1.95
+ $X2=0 $Y2=0
cc_365 N_A_495_390#_c_337_n N_A_309_390#_c_941_n 0.00541317f $X=2.832 $Y=0.415
+ $X2=0 $Y2=0
cc_366 N_A_495_390#_M1014_g N_A_309_390#_c_942_n 0.0189282f $X=4.04 $Y=0.9 $X2=0
+ $Y2=0
cc_367 N_A_495_390#_c_330_n N_A_309_390#_c_942_n 0.00349197f $X=4.305 $Y=0.415
+ $X2=0 $Y2=0
cc_368 N_A_495_390#_c_337_n N_A_309_390#_c_942_n 0.00470909f $X=2.832 $Y=0.415
+ $X2=0 $Y2=0
cc_369 N_A_495_390#_M1008_g N_A_309_390#_M1011_g 0.0118691f $X=3.41 $Y=2.525
+ $X2=0 $Y2=0
cc_370 N_A_495_390#_c_324_n N_A_309_390#_M1011_g 0.0050685f $X=4.04 $Y=1.405
+ $X2=0 $Y2=0
cc_371 N_A_495_390#_c_347_n N_A_309_390#_M1013_g 0.00727778f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_372 N_A_495_390#_c_327_n N_A_309_390#_c_943_n 0.0196921f $X=6.715 $Y=1.27
+ $X2=0 $Y2=0
cc_373 N_A_495_390#_c_334_n N_A_309_390#_c_943_n 0.0166975f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_374 N_A_495_390#_c_347_n N_A_309_390#_c_943_n 0.0260156f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_375 N_A_495_390#_c_340_n N_A_309_390#_c_943_n 0.00239794f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_376 N_A_495_390#_c_328_n N_A_309_390#_c_958_n 0.0196921f $X=6.355 $Y=1.27
+ $X2=0 $Y2=0
cc_377 N_A_495_390#_c_332_n N_A_309_390#_M1031_g 0.00912173f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_378 N_A_495_390#_c_334_n N_A_309_390#_M1031_g 0.00885461f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_379 N_A_495_390#_c_335_n N_A_309_390#_M1031_g 0.0230685f $X=7.37 $Y=1.015
+ $X2=0 $Y2=0
cc_380 N_A_495_390#_c_339_n N_A_309_390#_M1031_g 0.0213806f $X=6.88 $Y=1.18
+ $X2=0 $Y2=0
cc_381 N_A_495_390#_c_340_n N_A_309_390#_M1031_g 0.0123873f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_382 N_A_495_390#_M1012_d N_A_309_390#_c_975_n 0.00218798f $X=2.61 $Y=0.595
+ $X2=0 $Y2=0
cc_383 N_A_495_390#_c_329_n N_A_309_390#_c_975_n 0.0140921f $X=2.967 $Y=1.625
+ $X2=0 $Y2=0
cc_384 N_A_495_390#_c_337_n N_A_309_390#_c_975_n 0.00269441f $X=2.832 $Y=0.415
+ $X2=0 $Y2=0
cc_385 N_A_495_390#_M1012_d N_A_309_390#_c_947_n 0.00173384f $X=2.61 $Y=0.595
+ $X2=0 $Y2=0
cc_386 N_A_495_390#_c_329_n N_A_309_390#_c_947_n 0.0336426f $X=2.967 $Y=1.625
+ $X2=0 $Y2=0
cc_387 N_A_495_390#_c_336_n N_A_309_390#_c_947_n 0.0237964f $X=2.967 $Y=1.95
+ $X2=0 $Y2=0
cc_388 N_A_495_390#_c_336_n N_A_309_390#_c_962_n 0.0021988f $X=2.967 $Y=1.95
+ $X2=0 $Y2=0
cc_389 N_A_495_390#_c_332_n N_A_1525_212#_M1005_g 0.00108131f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_390 N_A_495_390#_c_335_n N_A_1525_212#_M1005_g 0.00485618f $X=7.37 $Y=1.015
+ $X2=0 $Y2=0
cc_391 N_A_495_390#_c_340_n N_A_1525_212#_M1005_g 0.00116217f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_392 N_A_495_390#_c_347_n N_A_1525_212#_c_1126_n 0.0212062f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_393 N_A_495_390#_c_345_n N_A_1525_212#_c_1128_n 0.0268843f $X=7.315 $Y=2.39
+ $X2=0 $Y2=0
cc_394 N_A_495_390#_c_334_n N_A_1525_212#_c_1118_n 9.8351e-19 $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_395 N_A_495_390#_c_334_n N_A_1525_212#_c_1123_n 0.00193736f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_396 N_A_495_390#_c_340_n N_A_1525_212#_c_1123_n 0.0239506f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_397 N_A_495_390#_c_340_n N_A_1525_212#_c_1124_n 0.00177987f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_398 N_A_495_390#_c_332_n N_A_1271_74#_M1003_d 0.00941894f $X=7.285 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_399 N_A_495_390#_c_332_n N_A_1271_74#_c_1259_n 0.00860077f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_400 N_A_495_390#_c_326_n N_A_1271_74#_c_1240_n 0.0041612f $X=6.28 $Y=1.195
+ $X2=0 $Y2=0
cc_401 N_A_495_390#_c_327_n N_A_1271_74#_c_1240_n 0.010955f $X=6.715 $Y=1.27
+ $X2=0 $Y2=0
cc_402 N_A_495_390#_c_334_n N_A_1271_74#_c_1240_n 0.00709969f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_403 N_A_495_390#_c_339_n N_A_1271_74#_c_1240_n 0.00131723f $X=6.88 $Y=1.18
+ $X2=0 $Y2=0
cc_404 N_A_495_390#_c_340_n N_A_1271_74#_c_1240_n 0.022475f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_405 N_A_495_390#_c_345_n N_A_1271_74#_c_1252_n 0.00181181f $X=7.315 $Y=2.39
+ $X2=0 $Y2=0
cc_406 N_A_495_390#_c_334_n N_A_1271_74#_c_1252_n 0.0315385f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_407 N_A_495_390#_c_347_n N_A_1271_74#_c_1252_n 0.00442904f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_408 N_A_495_390#_c_327_n N_A_1271_74#_c_1241_n 0.00400734f $X=6.715 $Y=1.27
+ $X2=0 $Y2=0
cc_409 N_A_495_390#_c_332_n N_A_1271_74#_c_1241_n 0.0414158f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_410 N_A_495_390#_c_335_n N_A_1271_74#_c_1241_n 0.0196081f $X=7.37 $Y=1.015
+ $X2=0 $Y2=0
cc_411 N_A_495_390#_c_339_n N_A_1271_74#_c_1241_n 0.00763158f $X=6.88 $Y=1.18
+ $X2=0 $Y2=0
cc_412 N_A_495_390#_c_340_n N_A_1271_74#_c_1241_n 0.0304853f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_413 N_A_495_390#_c_345_n N_A_1271_74#_c_1273_n 0.0126686f $X=7.315 $Y=2.39
+ $X2=0 $Y2=0
cc_414 N_A_495_390#_c_334_n N_A_1271_74#_c_1273_n 0.0234051f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_415 N_A_495_390#_c_347_n N_A_1271_74#_c_1273_n 0.00188634f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_416 N_A_495_390#_c_345_n N_A_1271_74#_c_1253_n 0.00196844f $X=7.315 $Y=2.39
+ $X2=0 $Y2=0
cc_417 N_A_495_390#_c_334_n N_A_1271_74#_c_1253_n 0.0428804f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_418 N_A_495_390#_c_347_n N_A_1271_74#_c_1253_n 0.00431063f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_419 N_A_495_390#_c_334_n N_A_1271_74#_c_1243_n 0.0142968f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_420 N_A_495_390#_c_327_n N_A_1271_74#_c_1244_n 0.00176995f $X=6.715 $Y=1.27
+ $X2=0 $Y2=0
cc_421 N_A_495_390#_c_334_n N_A_1271_74#_c_1244_n 0.00932939f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_422 N_A_495_390#_c_345_n N_VPWR_c_1463_n 0.00125875f $X=7.315 $Y=2.39 $X2=0
+ $Y2=0
cc_423 N_A_495_390#_c_345_n N_VPWR_c_1473_n 0.00391396f $X=7.315 $Y=2.39 $X2=0
+ $Y2=0
cc_424 N_A_495_390#_M1008_g N_VPWR_c_1455_n 9.39239e-19 $X=3.41 $Y=2.525 $X2=0
+ $Y2=0
cc_425 N_A_495_390#_c_345_n N_VPWR_c_1455_n 0.0052212f $X=7.315 $Y=2.39 $X2=0
+ $Y2=0
cc_426 N_A_495_390#_M1004_d N_A_30_78#_c_1624_n 0.00590153f $X=2.475 $Y=1.95
+ $X2=0 $Y2=0
cc_427 N_A_495_390#_c_336_n N_A_30_78#_c_1624_n 0.0263146f $X=2.967 $Y=1.95
+ $X2=0 $Y2=0
cc_428 N_A_495_390#_c_329_n N_A_30_78#_c_1616_n 0.00993888f $X=2.967 $Y=1.625
+ $X2=0 $Y2=0
cc_429 N_A_495_390#_c_323_n N_A_30_78#_c_1625_n 6.21821e-19 $X=3.41 $Y=1.99
+ $X2=0 $Y2=0
cc_430 N_A_495_390#_M1008_g N_A_30_78#_c_1625_n 0.0101303f $X=3.41 $Y=2.525
+ $X2=0 $Y2=0
cc_431 N_A_495_390#_c_343_n N_A_30_78#_c_1625_n 0.00243864f $X=3.825 $Y=1.73
+ $X2=0 $Y2=0
cc_432 N_A_495_390#_c_336_n N_A_30_78#_c_1625_n 0.00268506f $X=2.967 $Y=1.95
+ $X2=0 $Y2=0
cc_433 N_A_495_390#_c_323_n N_A_30_78#_c_1617_n 0.0022386f $X=3.41 $Y=1.99 $X2=0
+ $Y2=0
cc_434 N_A_495_390#_M1008_g N_A_30_78#_c_1617_n 0.00268539f $X=3.41 $Y=2.525
+ $X2=0 $Y2=0
cc_435 N_A_495_390#_c_343_n N_A_30_78#_c_1617_n 0.0133047f $X=3.825 $Y=1.73
+ $X2=0 $Y2=0
cc_436 N_A_495_390#_c_324_n N_A_30_78#_c_1617_n 0.00591355f $X=4.04 $Y=1.405
+ $X2=0 $Y2=0
cc_437 N_A_495_390#_c_329_n N_A_30_78#_c_1617_n 0.00791036f $X=2.967 $Y=1.625
+ $X2=0 $Y2=0
cc_438 N_A_495_390#_c_336_n N_A_30_78#_c_1617_n 0.0321608f $X=2.967 $Y=1.95
+ $X2=0 $Y2=0
cc_439 N_A_495_390#_c_323_n N_A_30_78#_c_1628_n 0.00119431f $X=3.41 $Y=1.99
+ $X2=0 $Y2=0
cc_440 N_A_495_390#_M1008_g N_A_30_78#_c_1628_n 0.00394881f $X=3.41 $Y=2.525
+ $X2=0 $Y2=0
cc_441 N_A_495_390#_c_336_n N_A_30_78#_c_1628_n 0.0242647f $X=2.967 $Y=1.95
+ $X2=0 $Y2=0
cc_442 N_A_495_390#_c_330_n N_A_30_78#_c_1619_n 0.0192833f $X=4.305 $Y=0.415
+ $X2=0 $Y2=0
cc_443 N_A_495_390#_c_336_n N_A_30_78#_c_1619_n 0.0027055f $X=2.967 $Y=1.95
+ $X2=0 $Y2=0
cc_444 N_A_495_390#_c_337_n N_A_30_78#_c_1619_n 0.0296536f $X=2.832 $Y=0.415
+ $X2=0 $Y2=0
cc_445 N_A_495_390#_c_323_n N_A_30_78#_c_1620_n 0.00361109f $X=3.41 $Y=1.99
+ $X2=0 $Y2=0
cc_446 N_A_495_390#_c_343_n N_A_30_78#_c_1620_n 5.77187e-19 $X=3.825 $Y=1.73
+ $X2=0 $Y2=0
cc_447 N_A_495_390#_M1014_g N_A_30_78#_c_1620_n 7.45465e-19 $X=4.04 $Y=0.9 $X2=0
+ $Y2=0
cc_448 N_A_495_390#_c_329_n N_A_30_78#_c_1620_n 0.00935975f $X=2.967 $Y=1.625
+ $X2=0 $Y2=0
cc_449 N_A_495_390#_c_336_n N_A_30_78#_c_1620_n 0.00633174f $X=2.967 $Y=1.95
+ $X2=0 $Y2=0
cc_450 N_A_495_390#_c_331_n N_VGND_M1001_d 0.0203479f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_451 N_A_495_390#_c_375_p N_VGND_M1001_d 0.00355743f $X=5.6 $Y=0.615 $X2=0
+ $Y2=0
cc_452 N_A_495_390#_c_333_n N_VGND_M1001_d 6.7108e-19 $X=5.685 $Y=0.34 $X2=0
+ $Y2=0
cc_453 N_A_495_390#_c_337_n N_VGND_c_1771_n 0.0302166f $X=2.832 $Y=0.415 $X2=0
+ $Y2=0
cc_454 N_A_495_390#_c_332_n N_VGND_c_1772_n 0.00865667f $X=7.285 $Y=0.34 $X2=0
+ $Y2=0
cc_455 N_A_495_390#_c_330_n N_VGND_c_1778_n 0.0540738f $X=4.305 $Y=0.415 $X2=0
+ $Y2=0
cc_456 N_A_495_390#_c_331_n N_VGND_c_1778_n 0.0402161f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_457 N_A_495_390#_c_375_p N_VGND_c_1778_n 0.00152296f $X=5.6 $Y=0.615 $X2=0
+ $Y2=0
cc_458 N_A_495_390#_c_333_n N_VGND_c_1778_n 0.0151294f $X=5.685 $Y=0.34 $X2=0
+ $Y2=0
cc_459 N_A_495_390#_c_337_n N_VGND_c_1778_n 0.0225906f $X=2.832 $Y=0.415 $X2=0
+ $Y2=0
cc_460 N_A_495_390#_c_338_n N_VGND_c_1778_n 0.0126667f $X=4.39 $Y=0.415 $X2=0
+ $Y2=0
cc_461 N_A_495_390#_c_326_n N_VGND_c_1779_n 0.00278271f $X=6.28 $Y=1.195 $X2=0
+ $Y2=0
cc_462 N_A_495_390#_c_331_n N_VGND_c_1779_n 0.00309688f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_463 N_A_495_390#_c_332_n N_VGND_c_1779_n 0.114324f $X=7.285 $Y=0.34 $X2=0
+ $Y2=0
cc_464 N_A_495_390#_c_333_n N_VGND_c_1779_n 0.0119604f $X=5.685 $Y=0.34 $X2=0
+ $Y2=0
cc_465 N_A_495_390#_c_326_n N_VGND_c_1788_n 0.00358928f $X=6.28 $Y=1.195 $X2=0
+ $Y2=0
cc_466 N_A_495_390#_c_330_n N_VGND_c_1788_n 0.0393214f $X=4.305 $Y=0.415 $X2=0
+ $Y2=0
cc_467 N_A_495_390#_c_331_n N_VGND_c_1788_n 0.0181439f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_468 N_A_495_390#_c_332_n N_VGND_c_1788_n 0.0653925f $X=7.285 $Y=0.34 $X2=0
+ $Y2=0
cc_469 N_A_495_390#_c_333_n N_VGND_c_1788_n 0.00656672f $X=5.685 $Y=0.34 $X2=0
+ $Y2=0
cc_470 N_A_495_390#_c_337_n N_VGND_c_1788_n 0.0156671f $X=2.832 $Y=0.415 $X2=0
+ $Y2=0
cc_471 N_A_495_390#_c_338_n N_VGND_c_1788_n 0.00552563f $X=4.39 $Y=0.415 $X2=0
+ $Y2=0
cc_472 N_A_495_390#_c_331_n A_901_138# 0.00102299f $X=5.515 $Y=0.7 $X2=-0.19
+ $Y2=-0.245
cc_473 N_A_839_359#_M1006_g N_RESET_B_c_605_n 0.00556991f $X=4.43 $Y=0.9 $X2=0
+ $Y2=0
cc_474 N_A_839_359#_M1006_g N_RESET_B_M1001_g 0.0488638f $X=4.43 $Y=0.9 $X2=0
+ $Y2=0
cc_475 N_A_839_359#_c_517_n N_RESET_B_M1001_g 0.00101158f $X=4.36 $Y=1.96 $X2=0
+ $Y2=0
cc_476 N_A_839_359#_c_518_n N_RESET_B_M1001_g 0.0120195f $X=5.855 $Y=1.04 $X2=0
+ $Y2=0
cc_477 N_A_839_359#_M1006_g N_RESET_B_c_608_n 0.0157284f $X=4.43 $Y=0.9 $X2=0
+ $Y2=0
cc_478 N_A_839_359#_c_517_n N_RESET_B_c_608_n 4.40421e-19 $X=4.36 $Y=1.96 $X2=0
+ $Y2=0
cc_479 N_A_839_359#_c_521_n N_RESET_B_c_616_n 0.0324725f $X=4.275 $Y=2.21 $X2=0
+ $Y2=0
cc_480 N_A_839_359#_c_518_n N_RESET_B_c_610_n 0.00269956f $X=5.855 $Y=1.04 $X2=0
+ $Y2=0
cc_481 N_A_839_359#_c_521_n N_RESET_B_c_620_n 0.0115222f $X=4.275 $Y=2.21 $X2=0
+ $Y2=0
cc_482 N_A_839_359#_c_517_n N_RESET_B_c_620_n 0.0162413f $X=4.36 $Y=1.96 $X2=0
+ $Y2=0
cc_483 N_A_839_359#_M1028_d N_RESET_B_c_622_n 0.00226165f $X=5.98 $Y=1.735 $X2=0
+ $Y2=0
cc_484 N_A_839_359#_c_524_n N_RESET_B_c_622_n 0.0386269f $X=6.18 $Y=2.02 $X2=0
+ $Y2=0
cc_485 N_A_839_359#_c_518_n N_A_697_463#_M1020_g 0.0124697f $X=5.855 $Y=1.04
+ $X2=0 $Y2=0
cc_486 N_A_839_359#_c_542_n N_A_697_463#_M1020_g 0.0104935f $X=6.02 $Y=0.86
+ $X2=0 $Y2=0
cc_487 N_A_839_359#_c_519_n N_A_697_463#_M1020_g 0.00268294f $X=6.02 $Y=1.042
+ $X2=0 $Y2=0
cc_488 N_A_839_359#_c_520_n N_A_697_463#_M1020_g 0.00639735f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_489 N_A_839_359#_c_519_n N_A_697_463#_c_814_n 0.00463727f $X=6.02 $Y=1.042
+ $X2=0 $Y2=0
cc_490 N_A_839_359#_c_520_n N_A_697_463#_c_814_n 0.0148463f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_491 N_A_839_359#_c_518_n N_A_697_463#_c_815_n 0.0091182f $X=5.855 $Y=1.04
+ $X2=0 $Y2=0
cc_492 N_A_839_359#_c_521_n N_A_697_463#_c_847_n 0.012984f $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_493 N_A_839_359#_c_517_n N_A_697_463#_c_847_n 0.00669016f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_494 N_A_839_359#_c_521_n N_A_697_463#_c_823_n 0.00402075f $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_495 N_A_839_359#_M1006_g N_A_697_463#_c_823_n 0.00141812f $X=4.43 $Y=0.9
+ $X2=0 $Y2=0
cc_496 N_A_839_359#_c_517_n N_A_697_463#_c_823_n 0.0385446f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_497 N_A_839_359#_M1006_g N_A_697_463#_c_816_n 0.00204128f $X=4.43 $Y=0.9
+ $X2=0 $Y2=0
cc_498 N_A_839_359#_c_517_n N_A_697_463#_c_816_n 0.0225894f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_499 N_A_839_359#_c_518_n N_A_697_463#_c_816_n 0.0137783f $X=5.855 $Y=1.04
+ $X2=0 $Y2=0
cc_500 N_A_839_359#_c_518_n N_A_697_463#_c_817_n 0.0680785f $X=5.855 $Y=1.04
+ $X2=0 $Y2=0
cc_501 N_A_839_359#_c_520_n N_A_697_463#_c_817_n 0.0134746f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_502 N_A_839_359#_M1006_g N_A_697_463#_c_818_n 0.00130595f $X=4.43 $Y=0.9
+ $X2=0 $Y2=0
cc_503 N_A_839_359#_c_539_n N_A_697_463#_c_818_n 0.00796739f $X=4.445 $Y=1.04
+ $X2=0 $Y2=0
cc_504 N_A_839_359#_c_521_n N_A_697_463#_c_826_n 0.0100296f $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_505 N_A_839_359#_c_521_n N_A_697_463#_c_819_n 0.00669879f $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_506 N_A_839_359#_M1006_g N_A_697_463#_c_819_n 0.00122789f $X=4.43 $Y=0.9
+ $X2=0 $Y2=0
cc_507 N_A_839_359#_c_517_n N_A_697_463#_c_819_n 0.071821f $X=4.36 $Y=1.96 $X2=0
+ $Y2=0
cc_508 N_A_839_359#_c_539_n N_A_697_463#_c_819_n 0.0059461f $X=4.445 $Y=1.04
+ $X2=0 $Y2=0
cc_509 N_A_839_359#_c_521_n N_A_697_463#_c_864_n 8.80638e-19 $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_510 N_A_839_359#_c_521_n N_A_309_390#_M1011_g 0.0422109f $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_511 N_A_839_359#_c_521_n N_A_309_390#_c_955_n 0.00987628f $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_512 N_A_839_359#_c_524_n N_A_309_390#_c_955_n 0.00434706f $X=6.18 $Y=2.02
+ $X2=0 $Y2=0
cc_513 N_A_839_359#_c_524_n N_A_309_390#_M1013_g 0.0106383f $X=6.18 $Y=2.02
+ $X2=0 $Y2=0
cc_514 N_A_839_359#_c_520_n N_A_309_390#_M1013_g 8.73808e-19 $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_515 N_A_839_359#_c_520_n N_A_309_390#_c_958_n 0.00135615f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_516 N_A_839_359#_c_519_n N_A_1271_74#_c_1240_n 0.00157956f $X=6.02 $Y=1.042
+ $X2=0 $Y2=0
cc_517 N_A_839_359#_c_520_n N_A_1271_74#_c_1240_n 0.0283811f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_518 N_A_839_359#_c_524_n N_A_1271_74#_c_1252_n 0.0250147f $X=6.18 $Y=2.02
+ $X2=0 $Y2=0
cc_519 N_A_839_359#_c_520_n N_A_1271_74#_c_1252_n 0.00658883f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_520 N_A_839_359#_c_520_n N_A_1271_74#_c_1244_n 0.0129728f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_521 N_A_839_359#_c_521_n N_VPWR_c_1460_n 0.00341322f $X=4.275 $Y=2.21 $X2=0
+ $Y2=0
cc_522 N_A_839_359#_c_518_n N_VPWR_c_1462_n 0.00367066f $X=5.855 $Y=1.04 $X2=0
+ $Y2=0
cc_523 N_A_839_359#_c_524_n N_VPWR_c_1462_n 0.0405057f $X=6.18 $Y=2.02 $X2=0
+ $Y2=0
cc_524 N_A_839_359#_c_524_n N_VPWR_c_1473_n 0.00666388f $X=6.18 $Y=2.02 $X2=0
+ $Y2=0
cc_525 N_A_839_359#_c_521_n N_VPWR_c_1455_n 9.39239e-19 $X=4.275 $Y=2.21 $X2=0
+ $Y2=0
cc_526 N_A_839_359#_c_524_n N_VPWR_c_1455_n 0.00905588f $X=6.18 $Y=2.02 $X2=0
+ $Y2=0
cc_527 N_A_839_359#_c_518_n N_VGND_M1001_d 0.0123032f $X=5.855 $Y=1.04 $X2=0
+ $Y2=0
cc_528 N_A_839_359#_c_539_n A_823_138# 0.00170982f $X=4.445 $Y=1.04 $X2=-0.19
+ $Y2=-0.245
cc_529 N_A_839_359#_c_518_n A_901_138# 0.00102299f $X=5.855 $Y=1.04 $X2=-0.19
+ $Y2=-0.245
cc_530 N_RESET_B_c_622_n N_A_697_463#_c_814_n 0.0121958f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_531 N_RESET_B_c_610_n N_A_697_463#_c_815_n 0.00991362f $X=4.88 $Y=1.26 $X2=0
+ $Y2=0
cc_532 N_RESET_B_c_622_n N_A_697_463#_c_815_n 0.00341453f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_533 N_RESET_B_c_620_n N_A_697_463#_c_822_n 0.00685662f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_534 N_RESET_B_c_620_n N_A_697_463#_c_847_n 0.0084236f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_535 N_RESET_B_c_608_n N_A_697_463#_c_823_n 0.00997697f $X=4.88 $Y=1.795 $X2=0
+ $Y2=0
cc_536 N_RESET_B_c_616_n N_A_697_463#_c_823_n 0.00283001f $X=4.895 $Y=2.21 $X2=0
+ $Y2=0
cc_537 N_RESET_B_c_620_n N_A_697_463#_c_823_n 0.0209922f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_538 N_RESET_B_c_623_n N_A_697_463#_c_823_n 0.00242233f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_539 N_RESET_B_c_624_n N_A_697_463#_c_823_n 0.0245177f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_540 N_RESET_B_c_610_n N_A_697_463#_c_816_n 0.00321182f $X=4.88 $Y=1.26 $X2=0
+ $Y2=0
cc_541 N_RESET_B_c_608_n N_A_697_463#_c_817_n 0.0121716f $X=4.88 $Y=1.795 $X2=0
+ $Y2=0
cc_542 N_RESET_B_c_616_n N_A_697_463#_c_817_n 0.00732939f $X=4.895 $Y=2.21 $X2=0
+ $Y2=0
cc_543 N_RESET_B_c_610_n N_A_697_463#_c_817_n 0.0034188f $X=4.88 $Y=1.26 $X2=0
+ $Y2=0
cc_544 N_RESET_B_c_620_n N_A_697_463#_c_817_n 0.00355574f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_545 N_RESET_B_c_622_n N_A_697_463#_c_817_n 0.0096202f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_546 N_RESET_B_c_623_n N_A_697_463#_c_817_n 0.00343479f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_547 N_RESET_B_c_624_n N_A_697_463#_c_817_n 0.019281f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_548 N_RESET_B_c_616_n N_A_697_463#_c_825_n 0.0147184f $X=4.895 $Y=2.21 $X2=0
+ $Y2=0
cc_549 N_RESET_B_c_620_n N_A_697_463#_c_825_n 0.00430979f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_550 N_RESET_B_c_622_n N_A_697_463#_c_825_n 7.06363e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_551 N_RESET_B_c_623_n N_A_697_463#_c_825_n 0.00875681f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_552 N_RESET_B_c_624_n N_A_697_463#_c_825_n 0.0209558f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_553 N_RESET_B_c_616_n N_A_697_463#_c_826_n 8.7672e-19 $X=4.895 $Y=2.21 $X2=0
+ $Y2=0
cc_554 N_RESET_B_c_620_n N_A_697_463#_c_826_n 0.00585268f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_555 N_RESET_B_c_620_n N_A_697_463#_c_819_n 0.0175355f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_556 N_RESET_B_c_620_n N_A_309_390#_c_949_n 0.00791509f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_557 N_RESET_B_c_605_n N_A_309_390#_c_939_n 0.010267f $X=4.715 $Y=0.18 $X2=0
+ $Y2=0
cc_558 N_RESET_B_c_620_n N_A_309_390#_c_950_n 4.52147e-19 $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_559 N_RESET_B_c_605_n N_A_309_390#_c_942_n 0.00526413f $X=4.715 $Y=0.18 $X2=0
+ $Y2=0
cc_560 N_RESET_B_c_620_n N_A_309_390#_M1011_g 0.00155315f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_561 N_RESET_B_c_616_n N_A_309_390#_c_955_n 0.00995786f $X=4.895 $Y=2.21 $X2=0
+ $Y2=0
cc_562 N_RESET_B_c_622_n N_A_309_390#_M1013_g 0.00854421f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_563 N_RESET_B_c_622_n N_A_309_390#_c_943_n 0.00771224f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_564 N_RESET_B_M1009_g N_A_309_390#_c_945_n 0.00310826f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_565 N_RESET_B_c_605_n N_A_309_390#_c_945_n 0.00989069f $X=4.715 $Y=0.18 $X2=0
+ $Y2=0
cc_566 N_RESET_B_c_620_n N_A_309_390#_c_946_n 0.00152612f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_567 N_RESET_B_c_611_n N_A_309_390#_c_946_n 0.00796614f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_568 N_RESET_B_c_612_n N_A_309_390#_c_946_n 0.0555521f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_569 N_RESET_B_c_620_n N_A_309_390#_c_947_n 0.00371929f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_570 N_RESET_B_M1009_g N_A_309_390#_c_948_n 0.0014141f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_571 N_RESET_B_c_612_n N_A_309_390#_c_948_n 8.33879e-19 $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_572 N_RESET_B_c_620_n N_A_309_390#_c_962_n 0.0253069f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_573 N_RESET_B_c_621_n N_A_309_390#_c_962_n 0.00246f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_574 N_RESET_B_c_612_n N_A_309_390#_c_962_n 0.0172519f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_575 N_RESET_B_c_627_n N_A_309_390#_c_962_n 0.00236342f $X=1.12 $Y=1.985 $X2=0
+ $Y2=0
cc_576 N_RESET_B_M1017_g N_A_1525_212#_M1005_g 0.0164487f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_577 N_RESET_B_c_617_n N_A_1525_212#_c_1126_n 0.0164306f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_578 N_RESET_B_c_622_n N_A_1525_212#_c_1126_n 4.99514e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_579 N_RESET_B_c_628_n N_A_1525_212#_c_1126_n 0.00182389f $X=8.23 $Y=2.11
+ $X2=0 $Y2=0
cc_580 N_RESET_B_c_617_n N_A_1525_212#_c_1127_n 0.00475599f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_581 N_RESET_B_c_622_n N_A_1525_212#_c_1127_n 0.0054475f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_582 N_RESET_B_c_625_n N_A_1525_212#_c_1127_n 0.00136519f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_583 N_RESET_B_c_628_n N_A_1525_212#_c_1127_n 0.00431246f $X=8.23 $Y=2.11
+ $X2=0 $Y2=0
cc_584 N_RESET_B_c_617_n N_A_1525_212#_c_1128_n 0.0121565f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_585 N_RESET_B_c_617_n N_A_1525_212#_c_1118_n 0.00147213f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_586 N_RESET_B_M1017_g N_A_1525_212#_c_1118_n 0.0193933f $X=8.24 $Y=0.615
+ $X2=0 $Y2=0
cc_587 N_RESET_B_c_622_n N_A_1525_212#_c_1118_n 0.00138661f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_588 N_RESET_B_c_625_n N_A_1525_212#_c_1118_n 8.33981e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_589 N_RESET_B_c_628_n N_A_1525_212#_c_1118_n 4.18149e-19 $X=8.23 $Y=2.11
+ $X2=0 $Y2=0
cc_590 N_RESET_B_M1017_g N_A_1525_212#_c_1119_n 0.013811f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_591 N_RESET_B_c_617_n N_A_1525_212#_c_1130_n 0.0117959f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_592 N_RESET_B_c_628_n N_A_1525_212#_c_1130_n 0.00789453f $X=8.23 $Y=2.11
+ $X2=0 $Y2=0
cc_593 N_RESET_B_M1017_g N_A_1525_212#_c_1120_n 0.00343438f $X=8.24 $Y=0.615
+ $X2=0 $Y2=0
cc_594 N_RESET_B_c_617_n N_A_1525_212#_c_1131_n 0.00297602f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_595 N_RESET_B_c_617_n N_A_1525_212#_c_1133_n 8.22326e-19 $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_596 N_RESET_B_c_628_n N_A_1525_212#_c_1133_n 0.0092621f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_597 N_RESET_B_M1017_g N_A_1525_212#_c_1123_n 0.00118187f $X=8.24 $Y=0.615
+ $X2=0 $Y2=0
cc_598 N_RESET_B_M1017_g N_A_1525_212#_c_1124_n 0.021263f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_599 N_RESET_B_c_622_n N_A_1271_74#_M1013_d 0.00308066f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_600 N_RESET_B_M1017_g N_A_1271_74#_M1018_g 0.0755988f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_601 N_RESET_B_c_617_n N_A_1271_74#_c_1245_n 0.00922978f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_602 N_RESET_B_M1017_g N_A_1271_74#_c_1245_n 0.00125436f $X=8.24 $Y=0.615
+ $X2=0 $Y2=0
cc_603 N_RESET_B_c_628_n N_A_1271_74#_c_1245_n 0.00157069f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_604 N_RESET_B_c_617_n N_A_1271_74#_c_1246_n 0.0124349f $X=8.235 $Y=2.39 $X2=0
+ $Y2=0
cc_605 N_RESET_B_M1017_g N_A_1271_74#_c_1237_n 0.0061479f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_606 N_RESET_B_c_622_n N_A_1271_74#_c_1252_n 0.0172254f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_607 N_RESET_B_c_622_n N_A_1271_74#_c_1273_n 0.0184591f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_608 N_RESET_B_c_622_n N_A_1271_74#_c_1253_n 0.0225824f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_609 N_RESET_B_c_625_n N_A_1271_74#_c_1253_n 0.00231685f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_610 N_RESET_B_c_628_n N_A_1271_74#_c_1253_n 0.023913f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_611 N_RESET_B_c_617_n N_A_1271_74#_c_1242_n 0.00115984f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_612 N_RESET_B_M1017_g N_A_1271_74#_c_1242_n 0.0108634f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_613 N_RESET_B_c_622_n N_A_1271_74#_c_1242_n 0.00539223f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_614 N_RESET_B_c_625_n N_A_1271_74#_c_1242_n 0.00832147f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_615 N_RESET_B_c_628_n N_A_1271_74#_c_1242_n 0.0386217f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_616 N_RESET_B_c_622_n N_A_1271_74#_c_1244_n 0.00603357f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_617 N_RESET_B_M1017_g N_A_1271_74#_c_1257_n 0.00100578f $X=8.24 $Y=0.615
+ $X2=0 $Y2=0
cc_618 N_RESET_B_c_620_n N_VPWR_M1027_d 0.00719239f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_619 N_RESET_B_c_619_n N_VPWR_c_1457_n 4.75294e-19 $X=0.962 $Y=2.465 $X2=0
+ $Y2=0
cc_620 N_RESET_B_c_619_n N_VPWR_c_1458_n 0.00674875f $X=0.962 $Y=2.465 $X2=0
+ $Y2=0
cc_621 N_RESET_B_c_616_n N_VPWR_c_1460_n 0.00360709f $X=4.895 $Y=2.21 $X2=0
+ $Y2=0
cc_622 N_RESET_B_c_608_n N_VPWR_c_1462_n 0.001224f $X=4.88 $Y=1.795 $X2=0 $Y2=0
cc_623 N_RESET_B_c_616_n N_VPWR_c_1462_n 0.0119495f $X=4.895 $Y=2.21 $X2=0 $Y2=0
cc_624 N_RESET_B_c_622_n N_VPWR_c_1462_n 0.0323618f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_625 N_RESET_B_c_623_n N_VPWR_c_1462_n 5.54746e-19 $X=5.185 $Y=2.035 $X2=0
+ $Y2=0
cc_626 N_RESET_B_c_624_n N_VPWR_c_1462_n 0.0200056f $X=5.04 $Y=2.035 $X2=0 $Y2=0
cc_627 N_RESET_B_c_617_n N_VPWR_c_1463_n 0.0075111f $X=8.235 $Y=2.39 $X2=0 $Y2=0
cc_628 N_RESET_B_c_625_n N_VPWR_c_1463_n 0.00200394f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_629 N_RESET_B_c_628_n N_VPWR_c_1463_n 0.0263442f $X=8.23 $Y=2.11 $X2=0 $Y2=0
cc_630 N_RESET_B_c_617_n N_VPWR_c_1468_n 0.00511025f $X=8.235 $Y=2.39 $X2=0
+ $Y2=0
cc_631 N_RESET_B_c_619_n N_VPWR_c_1470_n 0.00427882f $X=0.962 $Y=2.465 $X2=0
+ $Y2=0
cc_632 N_RESET_B_c_616_n N_VPWR_c_1455_n 9.39239e-19 $X=4.895 $Y=2.21 $X2=0
+ $Y2=0
cc_633 N_RESET_B_c_617_n N_VPWR_c_1455_n 0.0052212f $X=8.235 $Y=2.39 $X2=0 $Y2=0
cc_634 N_RESET_B_c_619_n N_VPWR_c_1455_n 0.00426366f $X=0.962 $Y=2.465 $X2=0
+ $Y2=0
cc_635 N_RESET_B_M1009_g N_A_30_78#_c_1614_n 0.00360662f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_636 N_RESET_B_c_619_n N_A_30_78#_c_1621_n 2.2337e-19 $X=0.962 $Y=2.465 $X2=0
+ $Y2=0
cc_637 N_RESET_B_M1009_g N_A_30_78#_c_1615_n 0.00906064f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_638 N_RESET_B_c_604_n N_A_30_78#_c_1615_n 0.0101328f $X=1.09 $Y=1.885 $X2=0
+ $Y2=0
cc_639 N_RESET_B_c_614_n N_A_30_78#_c_1615_n 0.00440557f $X=0.962 $Y=2.358 $X2=0
+ $Y2=0
cc_640 N_RESET_B_c_621_n N_A_30_78#_c_1615_n 0.00138196f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_641 N_RESET_B_c_611_n N_A_30_78#_c_1615_n 0.00561754f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_642 N_RESET_B_c_612_n N_A_30_78#_c_1615_n 0.0697209f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_643 N_RESET_B_c_627_n N_A_30_78#_c_1615_n 0.00573231f $X=1.12 $Y=1.985 $X2=0
+ $Y2=0
cc_644 N_RESET_B_c_614_n N_A_30_78#_c_1623_n 0.00724168f $X=0.962 $Y=2.358 $X2=0
+ $Y2=0
cc_645 N_RESET_B_c_619_n N_A_30_78#_c_1623_n 0.0115485f $X=0.962 $Y=2.465 $X2=0
+ $Y2=0
cc_646 N_RESET_B_c_620_n N_A_30_78#_c_1623_n 0.0267402f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_647 N_RESET_B_c_621_n N_A_30_78#_c_1623_n 0.00450272f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_648 N_RESET_B_c_612_n N_A_30_78#_c_1623_n 0.0176357f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_649 N_RESET_B_c_627_n N_A_30_78#_c_1623_n 0.00402806f $X=1.12 $Y=1.985 $X2=0
+ $Y2=0
cc_650 N_RESET_B_c_620_n N_A_30_78#_c_1624_n 0.00348055f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_651 N_RESET_B_c_620_n N_A_30_78#_c_1625_n 0.00930953f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_652 N_RESET_B_c_620_n N_A_30_78#_c_1617_n 0.0132413f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_653 N_RESET_B_M1009_g N_A_30_78#_c_1618_n 9.19771e-19 $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_654 N_RESET_B_c_614_n N_A_30_78#_c_1627_n 0.00195298f $X=0.962 $Y=2.358 $X2=0
+ $Y2=0
cc_655 N_RESET_B_c_619_n N_A_30_78#_c_1627_n 0.00460939f $X=0.962 $Y=2.465 $X2=0
+ $Y2=0
cc_656 N_RESET_B_c_627_n N_A_30_78#_c_1627_n 8.70663e-19 $X=1.12 $Y=1.985 $X2=0
+ $Y2=0
cc_657 N_RESET_B_c_620_n N_A_30_78#_c_1628_n 0.0114706f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_658 N_RESET_B_c_620_n N_A_30_78#_c_1620_n 0.00579057f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_659 N_RESET_B_M1009_g N_VGND_c_1769_n 0.00266841f $X=0.9 $Y=0.6 $X2=0 $Y2=0
cc_660 N_RESET_B_c_605_n N_VGND_c_1769_n 0.0210995f $X=4.715 $Y=0.18 $X2=0 $Y2=0
cc_661 N_RESET_B_c_611_n N_VGND_c_1769_n 0.00202483f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_662 N_RESET_B_c_612_n N_VGND_c_1769_n 0.0157941f $X=1.12 $Y=1.305 $X2=0 $Y2=0
cc_663 N_RESET_B_c_605_n N_VGND_c_1770_n 0.0227427f $X=4.715 $Y=0.18 $X2=0 $Y2=0
cc_664 N_RESET_B_c_605_n N_VGND_c_1771_n 0.0257653f $X=4.715 $Y=0.18 $X2=0 $Y2=0
cc_665 N_RESET_B_M1017_g N_VGND_c_1772_n 0.0104625f $X=8.24 $Y=0.615 $X2=0 $Y2=0
cc_666 N_RESET_B_c_606_n N_VGND_c_1777_n 0.00688107f $X=0.975 $Y=0.18 $X2=0
+ $Y2=0
cc_667 N_RESET_B_c_605_n N_VGND_c_1778_n 0.068465f $X=4.715 $Y=0.18 $X2=0 $Y2=0
cc_668 N_RESET_B_M1017_g N_VGND_c_1780_n 0.0045897f $X=8.24 $Y=0.615 $X2=0 $Y2=0
cc_669 N_RESET_B_c_605_n N_VGND_c_1788_n 0.0925422f $X=4.715 $Y=0.18 $X2=0 $Y2=0
cc_670 N_RESET_B_c_606_n N_VGND_c_1788_n 0.0110889f $X=0.975 $Y=0.18 $X2=0 $Y2=0
cc_671 N_RESET_B_M1017_g N_VGND_c_1788_n 0.0044912f $X=8.24 $Y=0.615 $X2=0 $Y2=0
cc_672 N_A_697_463#_c_822_n N_A_309_390#_c_951_n 0.00480341f $X=3.935 $Y=2.637
+ $X2=0 $Y2=0
cc_673 N_A_697_463#_c_819_n N_A_309_390#_c_940_n 2.98612e-19 $X=4.092 $Y=2.4
+ $X2=0 $Y2=0
cc_674 N_A_697_463#_c_818_n N_A_309_390#_c_942_n 0.00203816f $X=4.02 $Y=0.86
+ $X2=0 $Y2=0
cc_675 N_A_697_463#_c_819_n N_A_309_390#_c_942_n 9.89095e-19 $X=4.092 $Y=2.4
+ $X2=0 $Y2=0
cc_676 N_A_697_463#_c_822_n N_A_309_390#_M1011_g 0.00661964f $X=3.935 $Y=2.637
+ $X2=0 $Y2=0
cc_677 N_A_697_463#_c_826_n N_A_309_390#_M1011_g 0.0087208f $X=4.092 $Y=2.485
+ $X2=0 $Y2=0
cc_678 N_A_697_463#_c_819_n N_A_309_390#_M1011_g 0.00488974f $X=4.092 $Y=2.4
+ $X2=0 $Y2=0
cc_679 N_A_697_463#_c_814_n N_A_309_390#_c_955_n 0.0103562f $X=5.905 $Y=1.66
+ $X2=0 $Y2=0
cc_680 N_A_697_463#_c_847_n N_A_309_390#_c_955_n 0.00179819f $X=4.615 $Y=2.485
+ $X2=0 $Y2=0
cc_681 N_A_697_463#_c_825_n N_A_309_390#_c_955_n 0.00520468f $X=5.12 $Y=2.475
+ $X2=0 $Y2=0
cc_682 N_A_697_463#_c_826_n N_A_309_390#_c_955_n 0.00248246f $X=4.092 $Y=2.485
+ $X2=0 $Y2=0
cc_683 N_A_697_463#_c_864_n N_A_309_390#_c_955_n 0.00104522f $X=4.7 $Y=2.445
+ $X2=0 $Y2=0
cc_684 N_A_697_463#_c_814_n N_A_309_390#_M1013_g 0.0208385f $X=5.905 $Y=1.66
+ $X2=0 $Y2=0
cc_685 N_A_697_463#_c_814_n N_A_309_390#_c_958_n 0.0046962f $X=5.905 $Y=1.66
+ $X2=0 $Y2=0
cc_686 N_A_697_463#_c_847_n N_VPWR_M1010_d 0.00456062f $X=4.615 $Y=2.485 $X2=0
+ $Y2=0
cc_687 N_A_697_463#_c_864_n N_VPWR_M1010_d 0.00285796f $X=4.7 $Y=2.445 $X2=0
+ $Y2=0
cc_688 N_A_697_463#_c_847_n N_VPWR_c_1460_n 0.0153067f $X=4.615 $Y=2.485 $X2=0
+ $Y2=0
cc_689 N_A_697_463#_c_826_n N_VPWR_c_1460_n 7.88629e-19 $X=4.092 $Y=2.485 $X2=0
+ $Y2=0
cc_690 N_A_697_463#_c_864_n N_VPWR_c_1460_n 0.0116728f $X=4.7 $Y=2.445 $X2=0
+ $Y2=0
cc_691 N_A_697_463#_c_825_n N_VPWR_c_1461_n 0.00614556f $X=5.12 $Y=2.475 $X2=0
+ $Y2=0
cc_692 N_A_697_463#_c_864_n N_VPWR_c_1461_n 3.43985e-19 $X=4.7 $Y=2.445 $X2=0
+ $Y2=0
cc_693 N_A_697_463#_c_814_n N_VPWR_c_1462_n 0.0144085f $X=5.905 $Y=1.66 $X2=0
+ $Y2=0
cc_694 N_A_697_463#_c_815_n N_VPWR_c_1462_n 0.00770753f $X=5.73 $Y=1.41 $X2=0
+ $Y2=0
cc_695 N_A_697_463#_c_817_n N_VPWR_c_1462_n 0.0131953f $X=5.52 $Y=1.41 $X2=0
+ $Y2=0
cc_696 N_A_697_463#_c_825_n N_VPWR_c_1462_n 0.0177351f $X=5.12 $Y=2.475 $X2=0
+ $Y2=0
cc_697 N_A_697_463#_c_822_n N_VPWR_c_1472_n 0.00903319f $X=3.935 $Y=2.637 $X2=0
+ $Y2=0
cc_698 N_A_697_463#_c_847_n N_VPWR_c_1472_n 0.00181305f $X=4.615 $Y=2.485 $X2=0
+ $Y2=0
cc_699 N_A_697_463#_c_826_n N_VPWR_c_1472_n 0.00674063f $X=4.092 $Y=2.485 $X2=0
+ $Y2=0
cc_700 N_A_697_463#_c_814_n N_VPWR_c_1455_n 8.51577e-19 $X=5.905 $Y=1.66 $X2=0
+ $Y2=0
cc_701 N_A_697_463#_c_822_n N_VPWR_c_1455_n 0.0113949f $X=3.935 $Y=2.637 $X2=0
+ $Y2=0
cc_702 N_A_697_463#_c_847_n N_VPWR_c_1455_n 0.00437505f $X=4.615 $Y=2.485 $X2=0
+ $Y2=0
cc_703 N_A_697_463#_c_825_n N_VPWR_c_1455_n 0.011063f $X=5.12 $Y=2.475 $X2=0
+ $Y2=0
cc_704 N_A_697_463#_c_826_n N_VPWR_c_1455_n 0.00838337f $X=4.092 $Y=2.485 $X2=0
+ $Y2=0
cc_705 N_A_697_463#_c_864_n N_VPWR_c_1455_n 0.00141382f $X=4.7 $Y=2.445 $X2=0
+ $Y2=0
cc_706 N_A_697_463#_c_819_n N_A_30_78#_c_1616_n 0.00473328f $X=4.092 $Y=2.4
+ $X2=0 $Y2=0
cc_707 N_A_697_463#_M1008_d N_A_30_78#_c_1625_n 0.00293566f $X=3.485 $Y=2.315
+ $X2=0 $Y2=0
cc_708 N_A_697_463#_c_822_n N_A_30_78#_c_1625_n 0.0172064f $X=3.935 $Y=2.637
+ $X2=0 $Y2=0
cc_709 N_A_697_463#_c_819_n N_A_30_78#_c_1625_n 0.0135548f $X=4.092 $Y=2.4 $X2=0
+ $Y2=0
cc_710 N_A_697_463#_c_819_n N_A_30_78#_c_1617_n 0.057085f $X=4.092 $Y=2.4 $X2=0
+ $Y2=0
cc_711 N_A_697_463#_c_819_n N_A_30_78#_c_1628_n 0.00118944f $X=4.092 $Y=2.4
+ $X2=0 $Y2=0
cc_712 N_A_697_463#_c_818_n N_A_30_78#_c_1619_n 0.0144022f $X=4.02 $Y=0.86 $X2=0
+ $Y2=0
cc_713 N_A_697_463#_c_818_n N_A_30_78#_c_1620_n 0.0077624f $X=4.02 $Y=0.86 $X2=0
+ $Y2=0
cc_714 N_A_697_463#_c_819_n N_A_30_78#_c_1620_n 0.0137021f $X=4.092 $Y=2.4 $X2=0
+ $Y2=0
cc_715 N_A_697_463#_c_826_n A_798_463# 6.1426e-19 $X=4.092 $Y=2.485 $X2=-0.19
+ $Y2=-0.245
cc_716 N_A_697_463#_c_819_n A_798_463# 0.00100253f $X=4.092 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_717 N_A_697_463#_M1020_g N_VGND_c_1778_n 0.0012551f $X=5.805 $Y=0.74 $X2=0
+ $Y2=0
cc_718 N_A_697_463#_M1020_g N_VGND_c_1779_n 0.00278271f $X=5.805 $Y=0.74 $X2=0
+ $Y2=0
cc_719 N_A_697_463#_M1020_g N_VGND_c_1788_n 0.00358928f $X=5.805 $Y=0.74 $X2=0
+ $Y2=0
cc_720 N_A_309_390#_M1031_g N_A_1525_212#_M1005_g 0.0390746f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_721 N_A_309_390#_M1031_g N_A_1525_212#_c_1118_n 0.0184343f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_722 N_A_309_390#_M1031_g N_A_1525_212#_c_1123_n 4.84439e-19 $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_723 N_A_309_390#_M1031_g N_A_1525_212#_c_1124_n 0.0192269f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_724 N_A_309_390#_c_958_n N_A_1271_74#_c_1240_n 2.49182e-19 $X=6.485 $Y=1.66
+ $X2=0 $Y2=0
cc_725 N_A_309_390#_M1013_g N_A_1271_74#_c_1252_n 0.0101572f $X=6.41 $Y=2.31
+ $X2=0 $Y2=0
cc_726 N_A_309_390#_c_943_n N_A_1271_74#_c_1252_n 0.00688758f $X=7.255 $Y=1.66
+ $X2=0 $Y2=0
cc_727 N_A_309_390#_M1031_g N_A_1271_74#_c_1241_n 0.00513624f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_728 N_A_309_390#_M1031_g N_A_1271_74#_c_1243_n 0.00152295f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_729 N_A_309_390#_c_943_n N_A_1271_74#_c_1244_n 0.00544498f $X=7.255 $Y=1.66
+ $X2=0 $Y2=0
cc_730 N_A_309_390#_c_958_n N_A_1271_74#_c_1244_n 0.00457177f $X=6.485 $Y=1.66
+ $X2=0 $Y2=0
cc_731 N_A_309_390#_M1031_g N_A_1271_74#_c_1244_n 2.71569e-19 $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_732 N_A_309_390#_c_949_n N_VPWR_c_1459_n 0.00477194f $X=2.4 $Y=1.875 $X2=0
+ $Y2=0
cc_733 N_A_309_390#_c_950_n N_VPWR_c_1459_n 0.00317361f $X=2.89 $Y=3.075 $X2=0
+ $Y2=0
cc_734 N_A_309_390#_M1011_g N_VPWR_c_1460_n 0.00608962f $X=3.915 $Y=2.525 $X2=0
+ $Y2=0
cc_735 N_A_309_390#_c_955_n N_VPWR_c_1460_n 0.0250293f $X=6.32 $Y=3.15 $X2=0
+ $Y2=0
cc_736 N_A_309_390#_c_955_n N_VPWR_c_1461_n 0.0218823f $X=6.32 $Y=3.15 $X2=0
+ $Y2=0
cc_737 N_A_309_390#_c_955_n N_VPWR_c_1462_n 0.025868f $X=6.32 $Y=3.15 $X2=0
+ $Y2=0
cc_738 N_A_309_390#_M1013_g N_VPWR_c_1462_n 0.00120875f $X=6.41 $Y=2.31 $X2=0
+ $Y2=0
cc_739 N_A_309_390#_c_960_n N_VPWR_c_1462_n 0.00521396f $X=6.41 $Y=3.15 $X2=0
+ $Y2=0
cc_740 N_A_309_390#_c_949_n N_VPWR_c_1472_n 0.00446964f $X=2.4 $Y=1.875 $X2=0
+ $Y2=0
cc_741 N_A_309_390#_c_952_n N_VPWR_c_1472_n 0.0432568f $X=2.965 $Y=3.15 $X2=0
+ $Y2=0
cc_742 N_A_309_390#_c_955_n N_VPWR_c_1473_n 0.020324f $X=6.32 $Y=3.15 $X2=0
+ $Y2=0
cc_743 N_A_309_390#_c_949_n N_VPWR_c_1455_n 0.00542671f $X=2.4 $Y=1.875 $X2=0
+ $Y2=0
cc_744 N_A_309_390#_c_951_n N_VPWR_c_1455_n 0.0248529f $X=3.84 $Y=3.15 $X2=0
+ $Y2=0
cc_745 N_A_309_390#_c_952_n N_VPWR_c_1455_n 0.00684408f $X=2.965 $Y=3.15 $X2=0
+ $Y2=0
cc_746 N_A_309_390#_c_955_n N_VPWR_c_1455_n 0.0528687f $X=6.32 $Y=3.15 $X2=0
+ $Y2=0
cc_747 N_A_309_390#_c_959_n N_VPWR_c_1455_n 0.00416815f $X=3.915 $Y=3.15 $X2=0
+ $Y2=0
cc_748 N_A_309_390#_c_960_n N_VPWR_c_1455_n 0.0125228f $X=6.41 $Y=3.15 $X2=0
+ $Y2=0
cc_749 N_A_309_390#_c_945_n N_A_30_78#_c_1615_n 0.00404291f $X=1.71 $Y=0.625
+ $X2=0 $Y2=0
cc_750 N_A_309_390#_c_948_n N_A_30_78#_c_1615_n 0.00516976f $X=1.665 $Y=1.06
+ $X2=0 $Y2=0
cc_751 N_A_309_390#_c_962_n N_A_30_78#_c_1615_n 2.92206e-19 $X=1.69 $Y=2.075
+ $X2=0 $Y2=0
cc_752 N_A_309_390#_M1027_s N_A_30_78#_c_1623_n 0.00736088f $X=1.545 $Y=1.95
+ $X2=0 $Y2=0
cc_753 N_A_309_390#_c_949_n N_A_30_78#_c_1623_n 0.0174587f $X=2.4 $Y=1.875 $X2=0
+ $Y2=0
cc_754 N_A_309_390#_c_950_n N_A_30_78#_c_1623_n 4.31583e-19 $X=2.89 $Y=3.075
+ $X2=0 $Y2=0
cc_755 N_A_309_390#_c_962_n N_A_30_78#_c_1623_n 0.0250396f $X=1.69 $Y=2.075
+ $X2=0 $Y2=0
cc_756 N_A_309_390#_c_950_n N_A_30_78#_c_1624_n 0.00962873f $X=2.89 $Y=3.075
+ $X2=0 $Y2=0
cc_757 N_A_309_390#_c_940_n N_A_30_78#_c_1616_n 0.00469531f $X=3.465 $Y=1.275
+ $X2=0 $Y2=0
cc_758 N_A_309_390#_c_942_n N_A_30_78#_c_1616_n 0.00457746f $X=3.54 $Y=1.2 $X2=0
+ $Y2=0
cc_759 N_A_309_390#_M1011_g N_A_30_78#_c_1625_n 0.00145586f $X=3.915 $Y=2.525
+ $X2=0 $Y2=0
cc_760 N_A_309_390#_c_941_n N_A_30_78#_c_1617_n 0.00232594f $X=3.085 $Y=1.275
+ $X2=0 $Y2=0
cc_761 N_A_309_390#_c_950_n N_A_30_78#_c_1628_n 0.0121708f $X=2.89 $Y=3.075
+ $X2=0 $Y2=0
cc_762 N_A_309_390#_c_951_n N_A_30_78#_c_1628_n 0.00505717f $X=3.84 $Y=3.15
+ $X2=0 $Y2=0
cc_763 N_A_309_390#_c_940_n N_A_30_78#_c_1619_n 0.00197897f $X=3.465 $Y=1.275
+ $X2=0 $Y2=0
cc_764 N_A_309_390#_c_942_n N_A_30_78#_c_1619_n 0.00435411f $X=3.54 $Y=1.2 $X2=0
+ $Y2=0
cc_765 N_A_309_390#_c_940_n N_A_30_78#_c_1620_n 0.0143746f $X=3.465 $Y=1.275
+ $X2=0 $Y2=0
cc_766 N_A_309_390#_c_941_n N_A_30_78#_c_1620_n 7.53147e-19 $X=3.085 $Y=1.275
+ $X2=0 $Y2=0
cc_767 N_A_309_390#_c_975_n N_VGND_M1015_d 0.00805699f $X=2.445 $Y=1.06 $X2=0
+ $Y2=0
cc_768 N_A_309_390#_c_945_n N_VGND_c_1769_n 0.0395992f $X=1.71 $Y=0.625 $X2=0
+ $Y2=0
cc_769 N_A_309_390#_c_945_n N_VGND_c_1770_n 0.0186352f $X=1.71 $Y=0.625 $X2=0
+ $Y2=0
cc_770 N_A_309_390#_c_939_n N_VGND_c_1771_n 0.00242994f $X=2.535 $Y=1.41 $X2=0
+ $Y2=0
cc_771 N_A_309_390#_c_945_n N_VGND_c_1771_n 0.0172677f $X=1.71 $Y=0.625 $X2=0
+ $Y2=0
cc_772 N_A_309_390#_c_975_n N_VGND_c_1771_n 0.0233584f $X=2.445 $Y=1.06 $X2=0
+ $Y2=0
cc_773 N_A_309_390#_M1031_g N_VGND_c_1772_n 4.38128e-19 $X=7.33 $Y=0.615 $X2=0
+ $Y2=0
cc_774 N_A_309_390#_M1031_g N_VGND_c_1779_n 9.34015e-19 $X=7.33 $Y=0.615 $X2=0
+ $Y2=0
cc_775 N_A_309_390#_c_939_n N_VGND_c_1788_n 8.51577e-19 $X=2.535 $Y=1.41 $X2=0
+ $Y2=0
cc_776 N_A_309_390#_c_945_n N_VGND_c_1788_n 0.0137621f $X=1.71 $Y=0.625 $X2=0
+ $Y2=0
cc_777 N_A_1525_212#_c_1119_n N_A_1271_74#_M1018_g 0.0108536f $X=8.68 $Y=1.305
+ $X2=0 $Y2=0
cc_778 N_A_1525_212#_c_1120_n N_A_1271_74#_M1018_g 0.0236543f $X=8.845 $Y=0.615
+ $X2=0 $Y2=0
cc_779 N_A_1525_212#_c_1122_n N_A_1271_74#_M1018_g 0.00397247f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_780 N_A_1525_212#_c_1125_n N_A_1271_74#_M1018_g 0.00478437f $X=8.845 $Y=1.305
+ $X2=0 $Y2=0
cc_781 N_A_1525_212#_c_1131_n N_A_1271_74#_c_1245_n 7.30818e-19 $X=8.8 $Y=2.445
+ $X2=0 $Y2=0
cc_782 N_A_1525_212#_c_1132_n N_A_1271_74#_c_1245_n 0.0134689f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_783 N_A_1525_212#_c_1133_n N_A_1271_74#_c_1245_n 0.00277746f $X=8.885 $Y=2.19
+ $X2=0 $Y2=0
cc_784 N_A_1525_212#_c_1130_n N_A_1271_74#_c_1246_n 0.00989487f $X=8.715 $Y=2.61
+ $X2=0 $Y2=0
cc_785 N_A_1525_212#_c_1131_n N_A_1271_74#_c_1246_n 0.00482538f $X=8.8 $Y=2.445
+ $X2=0 $Y2=0
cc_786 N_A_1525_212#_c_1132_n N_A_1271_74#_c_1236_n 0.00213341f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_787 N_A_1525_212#_c_1122_n N_A_1271_74#_c_1236_n 0.0139731f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_788 N_A_1525_212#_c_1133_n N_A_1271_74#_c_1237_n 0.0010617f $X=8.885 $Y=2.19
+ $X2=0 $Y2=0
cc_789 N_A_1525_212#_c_1121_n N_A_1271_74#_c_1237_n 0.00714341f $X=9.205
+ $Y=1.305 $X2=0 $Y2=0
cc_790 N_A_1525_212#_c_1122_n N_A_1271_74#_c_1237_n 0.00618579f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_791 N_A_1525_212#_c_1125_n N_A_1271_74#_c_1237_n 0.00565398f $X=8.845
+ $Y=1.305 $X2=0 $Y2=0
cc_792 N_A_1525_212#_c_1122_n N_A_1271_74#_c_1249_n 0.00269774f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_793 N_A_1525_212#_c_1131_n N_A_1271_74#_c_1250_n 7.46191e-19 $X=8.8 $Y=2.445
+ $X2=0 $Y2=0
cc_794 N_A_1525_212#_c_1132_n N_A_1271_74#_c_1250_n 0.00172099f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_795 N_A_1525_212#_c_1122_n N_A_1271_74#_c_1250_n 0.00125184f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_796 N_A_1525_212#_c_1120_n N_A_1271_74#_M1019_g 0.00350395f $X=8.845 $Y=0.615
+ $X2=0 $Y2=0
cc_797 N_A_1525_212#_c_1121_n N_A_1271_74#_M1019_g 0.00377053f $X=9.205 $Y=1.305
+ $X2=0 $Y2=0
cc_798 N_A_1525_212#_c_1122_n N_A_1271_74#_M1019_g 0.00338537f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_799 N_A_1525_212#_c_1128_n N_A_1271_74#_c_1253_n 0.00151725f $X=7.735 $Y=2.39
+ $X2=0 $Y2=0
cc_800 N_A_1525_212#_c_1118_n N_A_1271_74#_c_1253_n 0.0136876f $X=7.735 $Y=1.975
+ $X2=0 $Y2=0
cc_801 N_A_1525_212#_c_1126_n N_A_1271_74#_c_1242_n 2.78684e-19 $X=7.735
+ $Y=2.065 $X2=0 $Y2=0
cc_802 N_A_1525_212#_c_1118_n N_A_1271_74#_c_1242_n 0.0105727f $X=7.735 $Y=1.975
+ $X2=0 $Y2=0
cc_803 N_A_1525_212#_c_1119_n N_A_1271_74#_c_1242_n 0.0522284f $X=8.68 $Y=1.305
+ $X2=0 $Y2=0
cc_804 N_A_1525_212#_c_1123_n N_A_1271_74#_c_1242_n 0.023491f $X=7.79 $Y=1.225
+ $X2=0 $Y2=0
cc_805 N_A_1525_212#_c_1124_n N_A_1271_74#_c_1242_n 0.00116263f $X=7.79 $Y=1.225
+ $X2=0 $Y2=0
cc_806 N_A_1525_212#_c_1125_n N_A_1271_74#_c_1242_n 0.00190438f $X=8.845
+ $Y=1.305 $X2=0 $Y2=0
cc_807 N_A_1525_212#_c_1130_n N_A_1271_74#_c_1257_n 2.74753e-19 $X=8.715 $Y=2.61
+ $X2=0 $Y2=0
cc_808 N_A_1525_212#_c_1132_n N_A_1271_74#_c_1257_n 0.00882758f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_809 N_A_1525_212#_c_1133_n N_A_1271_74#_c_1257_n 0.0119175f $X=8.885 $Y=2.19
+ $X2=0 $Y2=0
cc_810 N_A_1525_212#_c_1121_n N_A_1271_74#_c_1257_n 0.00177485f $X=9.205
+ $Y=1.305 $X2=0 $Y2=0
cc_811 N_A_1525_212#_c_1122_n N_A_1271_74#_c_1257_n 0.0242588f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_812 N_A_1525_212#_c_1125_n N_A_1271_74#_c_1257_n 0.0257641f $X=8.845 $Y=1.305
+ $X2=0 $Y2=0
cc_813 N_A_1525_212#_c_1132_n N_A_1921_409#_c_1399_n 0.011653f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_814 N_A_1525_212#_c_1122_n N_A_1921_409#_c_1399_n 0.00461168f $X=9.29
+ $Y=2.105 $X2=0 $Y2=0
cc_815 N_A_1525_212#_c_1120_n N_A_1921_409#_c_1391_n 0.00484112f $X=8.845
+ $Y=0.615 $X2=0 $Y2=0
cc_816 N_A_1525_212#_c_1121_n N_A_1921_409#_c_1391_n 0.00459026f $X=9.205
+ $Y=1.305 $X2=0 $Y2=0
cc_817 N_A_1525_212#_c_1122_n N_A_1921_409#_c_1392_n 0.0210733f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_818 N_A_1525_212#_c_1121_n N_A_1921_409#_c_1393_n 0.00528833f $X=9.205
+ $Y=1.305 $X2=0 $Y2=0
cc_819 N_A_1525_212#_c_1122_n N_A_1921_409#_c_1393_n 0.0123556f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_820 N_A_1525_212#_c_1132_n N_VPWR_M1033_d 0.00763182f $X=9.205 $Y=2.19 $X2=0
+ $Y2=0
cc_821 N_A_1525_212#_c_1122_n N_VPWR_M1033_d 0.00173132f $X=9.29 $Y=2.105 $X2=0
+ $Y2=0
cc_822 N_A_1525_212#_c_1128_n N_VPWR_c_1463_n 0.0101713f $X=7.735 $Y=2.39 $X2=0
+ $Y2=0
cc_823 N_A_1525_212#_c_1130_n N_VPWR_c_1463_n 0.0142734f $X=8.715 $Y=2.61 $X2=0
+ $Y2=0
cc_824 N_A_1525_212#_c_1130_n N_VPWR_c_1464_n 0.0232957f $X=8.715 $Y=2.61 $X2=0
+ $Y2=0
cc_825 N_A_1525_212#_c_1132_n N_VPWR_c_1464_n 0.0245347f $X=9.205 $Y=2.19 $X2=0
+ $Y2=0
cc_826 N_A_1525_212#_c_1130_n N_VPWR_c_1468_n 0.01191f $X=8.715 $Y=2.61 $X2=0
+ $Y2=0
cc_827 N_A_1525_212#_c_1128_n N_VPWR_c_1473_n 0.00470366f $X=7.735 $Y=2.39 $X2=0
+ $Y2=0
cc_828 N_A_1525_212#_c_1128_n N_VPWR_c_1455_n 0.00473388f $X=7.735 $Y=2.39 $X2=0
+ $Y2=0
cc_829 N_A_1525_212#_c_1130_n N_VPWR_c_1455_n 0.0185129f $X=8.715 $Y=2.61 $X2=0
+ $Y2=0
cc_830 N_A_1525_212#_M1005_g N_VGND_c_1772_n 0.00870177f $X=7.72 $Y=0.615 $X2=0
+ $Y2=0
cc_831 N_A_1525_212#_c_1119_n N_VGND_c_1772_n 0.00751614f $X=8.68 $Y=1.305 $X2=0
+ $Y2=0
cc_832 N_A_1525_212#_c_1120_n N_VGND_c_1772_n 0.0106511f $X=8.845 $Y=0.615 $X2=0
+ $Y2=0
cc_833 N_A_1525_212#_c_1123_n N_VGND_c_1772_n 0.00718492f $X=7.79 $Y=1.225 $X2=0
+ $Y2=0
cc_834 N_A_1525_212#_c_1124_n N_VGND_c_1772_n 9.12984e-19 $X=7.79 $Y=1.225 $X2=0
+ $Y2=0
cc_835 N_A_1525_212#_c_1120_n N_VGND_c_1773_n 0.045283f $X=8.845 $Y=0.615 $X2=0
+ $Y2=0
cc_836 N_A_1525_212#_c_1121_n N_VGND_c_1773_n 0.0132803f $X=9.205 $Y=1.305 $X2=0
+ $Y2=0
cc_837 N_A_1525_212#_M1005_g N_VGND_c_1779_n 0.0045897f $X=7.72 $Y=0.615 $X2=0
+ $Y2=0
cc_838 N_A_1525_212#_c_1120_n N_VGND_c_1780_n 0.0127604f $X=8.845 $Y=0.615 $X2=0
+ $Y2=0
cc_839 N_A_1525_212#_M1005_g N_VGND_c_1788_n 0.0044912f $X=7.72 $Y=0.615 $X2=0
+ $Y2=0
cc_840 N_A_1525_212#_c_1120_n N_VGND_c_1788_n 0.011834f $X=8.845 $Y=0.615 $X2=0
+ $Y2=0
cc_841 N_A_1271_74#_c_1245_n N_A_1921_409#_c_1399_n 5.28212e-19 $X=8.945 $Y=2.3
+ $X2=0 $Y2=0
cc_842 N_A_1271_74#_c_1246_n N_A_1921_409#_c_1399_n 3.28834e-19 $X=8.945 $Y=2.39
+ $X2=0 $Y2=0
cc_843 N_A_1271_74#_c_1250_n N_A_1921_409#_c_1399_n 0.0159253f $X=9.53 $Y=1.97
+ $X2=0 $Y2=0
cc_844 N_A_1271_74#_c_1239_n N_A_1921_409#_c_1399_n 0.0016406f $X=9.562 $Y=1.63
+ $X2=0 $Y2=0
cc_845 N_A_1271_74#_M1019_g N_A_1921_409#_c_1391_n 0.0181066f $X=9.61 $Y=0.74
+ $X2=0 $Y2=0
cc_846 N_A_1271_74#_c_1249_n N_A_1921_409#_c_1392_n 0.00666991f $X=9.53 $Y=1.88
+ $X2=0 $Y2=0
cc_847 N_A_1271_74#_c_1250_n N_A_1921_409#_c_1392_n 0.00141733f $X=9.53 $Y=1.97
+ $X2=0 $Y2=0
cc_848 N_A_1271_74#_c_1239_n N_A_1921_409#_c_1392_n 0.00365747f $X=9.562 $Y=1.63
+ $X2=0 $Y2=0
cc_849 N_A_1271_74#_M1019_g N_A_1921_409#_c_1393_n 0.00613547f $X=9.61 $Y=0.74
+ $X2=0 $Y2=0
cc_850 N_A_1271_74#_c_1239_n N_A_1921_409#_c_1393_n 0.00242696f $X=9.562 $Y=1.63
+ $X2=0 $Y2=0
cc_851 N_A_1271_74#_M1019_g N_A_1921_409#_c_1394_n 0.0181431f $X=9.61 $Y=0.74
+ $X2=0 $Y2=0
cc_852 N_A_1271_74#_c_1253_n N_VPWR_c_1463_n 0.00184051f $X=7.54 $Y=2.475 $X2=0
+ $Y2=0
cc_853 N_A_1271_74#_c_1246_n N_VPWR_c_1464_n 0.0100164f $X=8.945 $Y=2.39 $X2=0
+ $Y2=0
cc_854 N_A_1271_74#_c_1250_n N_VPWR_c_1464_n 0.00627469f $X=9.53 $Y=1.97 $X2=0
+ $Y2=0
cc_855 N_A_1271_74#_c_1250_n N_VPWR_c_1465_n 0.00466121f $X=9.53 $Y=1.97 $X2=0
+ $Y2=0
cc_856 N_A_1271_74#_c_1246_n N_VPWR_c_1468_n 0.00511015f $X=8.945 $Y=2.39 $X2=0
+ $Y2=0
cc_857 N_A_1271_74#_c_1273_n N_VPWR_c_1473_n 0.0207747f $X=7.455 $Y=2.64 $X2=0
+ $Y2=0
cc_858 N_A_1271_74#_c_1367_p N_VPWR_c_1473_n 0.00391127f $X=6.685 $Y=2.64 $X2=0
+ $Y2=0
cc_859 N_A_1271_74#_c_1250_n N_VPWR_c_1474_n 0.00510653f $X=9.53 $Y=1.97 $X2=0
+ $Y2=0
cc_860 N_A_1271_74#_c_1246_n N_VPWR_c_1455_n 0.0052212f $X=8.945 $Y=2.39 $X2=0
+ $Y2=0
cc_861 N_A_1271_74#_c_1250_n N_VPWR_c_1455_n 0.0052212f $X=9.53 $Y=1.97 $X2=0
+ $Y2=0
cc_862 N_A_1271_74#_c_1273_n N_VPWR_c_1455_n 0.029938f $X=7.455 $Y=2.64 $X2=0
+ $Y2=0
cc_863 N_A_1271_74#_c_1367_p N_VPWR_c_1455_n 0.00557315f $X=6.685 $Y=2.64 $X2=0
+ $Y2=0
cc_864 N_A_1271_74#_c_1273_n A_1478_493# 0.00315877f $X=7.455 $Y=2.64 $X2=-0.19
+ $Y2=-0.245
cc_865 N_A_1271_74#_M1018_g N_VGND_c_1772_n 0.00147575f $X=8.63 $Y=0.615 $X2=0
+ $Y2=0
cc_866 N_A_1271_74#_M1018_g N_VGND_c_1773_n 0.00438924f $X=8.63 $Y=0.615 $X2=0
+ $Y2=0
cc_867 N_A_1271_74#_c_1236_n N_VGND_c_1773_n 0.00293701f $X=9.44 $Y=1.63 $X2=0
+ $Y2=0
cc_868 N_A_1271_74#_M1019_g N_VGND_c_1773_n 0.00488092f $X=9.61 $Y=0.74 $X2=0
+ $Y2=0
cc_869 N_A_1271_74#_M1019_g N_VGND_c_1774_n 0.00412165f $X=9.61 $Y=0.74 $X2=0
+ $Y2=0
cc_870 N_A_1271_74#_M1018_g N_VGND_c_1780_n 0.00527282f $X=8.63 $Y=0.615 $X2=0
+ $Y2=0
cc_871 N_A_1271_74#_M1019_g N_VGND_c_1781_n 0.00434272f $X=9.61 $Y=0.74 $X2=0
+ $Y2=0
cc_872 N_A_1271_74#_M1018_g N_VGND_c_1788_n 0.00534666f $X=8.63 $Y=0.615 $X2=0
+ $Y2=0
cc_873 N_A_1271_74#_M1019_g N_VGND_c_1788_n 0.00830282f $X=9.61 $Y=0.74 $X2=0
+ $Y2=0
cc_874 N_A_1921_409#_c_1399_n N_VPWR_c_1464_n 0.0180508f $X=9.755 $Y=2.195 $X2=0
+ $Y2=0
cc_875 N_A_1921_409#_c_1383_n N_VPWR_c_1465_n 0.00728605f $X=10.475 $Y=1.375
+ $X2=0 $Y2=0
cc_876 N_A_1921_409#_c_1396_n N_VPWR_c_1465_n 0.0053787f $X=10.565 $Y=1.765
+ $X2=0 $Y2=0
cc_877 N_A_1921_409#_c_1392_n N_VPWR_c_1465_n 0.0728323f $X=9.755 $Y=2.03 $X2=0
+ $Y2=0
cc_878 N_A_1921_409#_c_1393_n N_VPWR_c_1465_n 0.00302521f $X=10.09 $Y=1.465
+ $X2=0 $Y2=0
cc_879 N_A_1921_409#_c_1394_n N_VPWR_c_1465_n 0.00372647f $X=10.09 $Y=1.375
+ $X2=0 $Y2=0
cc_880 N_A_1921_409#_c_1398_n N_VPWR_c_1467_n 0.00835395f $X=11.015 $Y=1.765
+ $X2=0 $Y2=0
cc_881 N_A_1921_409#_c_1399_n N_VPWR_c_1474_n 0.0111926f $X=9.755 $Y=2.195 $X2=0
+ $Y2=0
cc_882 N_A_1921_409#_c_1396_n N_VPWR_c_1475_n 0.00461464f $X=10.565 $Y=1.765
+ $X2=0 $Y2=0
cc_883 N_A_1921_409#_c_1398_n N_VPWR_c_1475_n 0.00417277f $X=11.015 $Y=1.765
+ $X2=0 $Y2=0
cc_884 N_A_1921_409#_c_1396_n N_VPWR_c_1455_n 0.00912521f $X=10.565 $Y=1.765
+ $X2=0 $Y2=0
cc_885 N_A_1921_409#_c_1398_n N_VPWR_c_1455_n 0.00769367f $X=11.015 $Y=1.765
+ $X2=0 $Y2=0
cc_886 N_A_1921_409#_c_1399_n N_VPWR_c_1455_n 0.0115381f $X=9.755 $Y=2.195 $X2=0
+ $Y2=0
cc_887 N_A_1921_409#_c_1384_n Q 0.00718159f $X=10.565 $Y=1.675 $X2=0 $Y2=0
cc_888 N_A_1921_409#_c_1396_n Q 0.00700399f $X=10.565 $Y=1.765 $X2=0 $Y2=0
cc_889 N_A_1921_409#_M1029_g Q 0.0157053f $X=10.6 $Y=0.74 $X2=0 $Y2=0
cc_890 N_A_1921_409#_c_1386_n Q 0.00813241f $X=10.925 $Y=1.375 $X2=0 $Y2=0
cc_891 N_A_1921_409#_c_1387_n Q 0.0128965f $X=11.015 $Y=1.675 $X2=0 $Y2=0
cc_892 N_A_1921_409#_c_1398_n Q 0.0235958f $X=11.015 $Y=1.765 $X2=0 $Y2=0
cc_893 N_A_1921_409#_M1032_g Q 0.0192861f $X=11.03 $Y=0.74 $X2=0 $Y2=0
cc_894 N_A_1921_409#_c_1389_n Q 0.00396751f $X=10.575 $Y=1.375 $X2=0 $Y2=0
cc_895 N_A_1921_409#_c_1390_n Q 0.00693891f $X=11.015 $Y=1.375 $X2=0 $Y2=0
cc_896 N_A_1921_409#_c_1391_n Q 0.00478422f $X=9.825 $Y=0.515 $X2=0 $Y2=0
cc_897 N_A_1921_409#_c_1393_n Q 0.0113958f $X=10.09 $Y=1.465 $X2=0 $Y2=0
cc_898 N_A_1921_409#_c_1394_n Q 5.0889e-19 $X=10.09 $Y=1.375 $X2=0 $Y2=0
cc_899 N_A_1921_409#_c_1391_n N_VGND_c_1773_n 0.0258169f $X=9.825 $Y=0.515 $X2=0
+ $Y2=0
cc_900 N_A_1921_409#_M1029_g N_VGND_c_1774_n 0.00647412f $X=10.6 $Y=0.74 $X2=0
+ $Y2=0
cc_901 N_A_1921_409#_c_1391_n N_VGND_c_1774_n 0.051504f $X=9.825 $Y=0.515 $X2=0
+ $Y2=0
cc_902 N_A_1921_409#_c_1394_n N_VGND_c_1774_n 0.0102912f $X=10.09 $Y=1.375 $X2=0
+ $Y2=0
cc_903 N_A_1921_409#_M1032_g N_VGND_c_1776_n 0.00647412f $X=11.03 $Y=0.74 $X2=0
+ $Y2=0
cc_904 N_A_1921_409#_c_1391_n N_VGND_c_1781_n 0.0145639f $X=9.825 $Y=0.515 $X2=0
+ $Y2=0
cc_905 N_A_1921_409#_M1029_g N_VGND_c_1782_n 0.00434272f $X=10.6 $Y=0.74 $X2=0
+ $Y2=0
cc_906 N_A_1921_409#_M1032_g N_VGND_c_1782_n 0.00434272f $X=11.03 $Y=0.74 $X2=0
+ $Y2=0
cc_907 N_A_1921_409#_M1029_g N_VGND_c_1788_n 0.00825283f $X=10.6 $Y=0.74 $X2=0
+ $Y2=0
cc_908 N_A_1921_409#_M1032_g N_VGND_c_1788_n 0.00823925f $X=11.03 $Y=0.74 $X2=0
+ $Y2=0
cc_909 N_A_1921_409#_c_1391_n N_VGND_c_1788_n 0.0119984f $X=9.825 $Y=0.515 $X2=0
+ $Y2=0
cc_910 N_VPWR_c_1457_n N_A_30_78#_c_1621_n 0.0230711f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_911 N_VPWR_c_1458_n N_A_30_78#_c_1621_n 0.00966405f $X=1.18 $Y=2.815 $X2=0
+ $Y2=0
cc_912 N_VPWR_c_1470_n N_A_30_78#_c_1621_n 0.00879902f $X=1.015 $Y=3.33 $X2=0
+ $Y2=0
cc_913 N_VPWR_c_1455_n N_A_30_78#_c_1621_n 0.007299f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_914 N_VPWR_M1023_d N_A_30_78#_c_1623_n 0.00245596f $X=1.02 $Y=2.54 $X2=0
+ $Y2=0
cc_915 N_VPWR_M1027_d N_A_30_78#_c_1623_n 0.00602617f $X=1.98 $Y=1.95 $X2=0
+ $Y2=0
cc_916 N_VPWR_c_1458_n N_A_30_78#_c_1623_n 0.0212934f $X=1.18 $Y=2.815 $X2=0
+ $Y2=0
cc_917 N_VPWR_c_1459_n N_A_30_78#_c_1623_n 0.0205269f $X=2.12 $Y=2.825 $X2=0
+ $Y2=0
cc_918 N_VPWR_c_1471_n N_A_30_78#_c_1623_n 0.00722345f $X=1.955 $Y=3.33 $X2=0
+ $Y2=0
cc_919 N_VPWR_c_1472_n N_A_30_78#_c_1623_n 0.00237421f $X=4.42 $Y=3.33 $X2=0
+ $Y2=0
cc_920 N_VPWR_c_1455_n N_A_30_78#_c_1623_n 0.028103f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_921 N_VPWR_c_1472_n N_A_30_78#_c_1624_n 0.00637223f $X=4.42 $Y=3.33 $X2=0
+ $Y2=0
cc_922 N_VPWR_c_1455_n N_A_30_78#_c_1624_n 0.0116928f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_923 N_VPWR_c_1457_n N_A_30_78#_c_1627_n 0.00766055f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_924 N_VPWR_c_1470_n N_A_30_78#_c_1627_n 2.70505e-19 $X=1.015 $Y=3.33 $X2=0
+ $Y2=0
cc_925 N_VPWR_c_1455_n N_A_30_78#_c_1627_n 0.00140703f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_926 N_VPWR_c_1472_n N_A_30_78#_c_1628_n 0.00674442f $X=4.42 $Y=3.33 $X2=0
+ $Y2=0
cc_927 N_VPWR_c_1455_n N_A_30_78#_c_1628_n 0.00974055f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_928 N_VPWR_c_1465_n Q 0.00316191f $X=10.315 $Y=1.985 $X2=0 $Y2=0
cc_929 N_VPWR_c_1467_n Q 0.0862588f $X=11.24 $Y=1.985 $X2=0 $Y2=0
cc_930 N_VPWR_c_1475_n Q 0.0145191f $X=11.155 $Y=3.33 $X2=0 $Y2=0
cc_931 N_VPWR_c_1455_n Q 0.011926f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_932 N_A_30_78#_c_1614_n A_117_78# 0.00232882f $X=0.665 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_933 N_A_30_78#_c_1614_n N_VGND_c_1769_n 0.00732263f $X=0.665 $Y=0.745 $X2=0
+ $Y2=0
cc_934 N_A_30_78#_c_1618_n N_VGND_c_1769_n 0.00454959f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_935 N_A_30_78#_c_1614_n N_VGND_c_1777_n 0.00539861f $X=0.665 $Y=0.745 $X2=0
+ $Y2=0
cc_936 N_A_30_78#_c_1618_n N_VGND_c_1777_n 0.0131067f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_937 N_A_30_78#_c_1614_n N_VGND_c_1788_n 0.0106165f $X=0.665 $Y=0.745 $X2=0
+ $Y2=0
cc_938 N_A_30_78#_c_1618_n N_VGND_c_1788_n 0.0117869f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_939 Q N_VGND_c_1774_n 0.0294122f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_940 Q N_VGND_c_1776_n 0.0294122f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_941 Q N_VGND_c_1782_n 0.0144922f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_942 Q N_VGND_c_1788_n 0.0118826f $X=10.715 $Y=0.47 $X2=0 $Y2=0
