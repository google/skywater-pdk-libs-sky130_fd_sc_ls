* NGSPICE file created from sky130_fd_sc_ls__o21a_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_116_387# A2 a_216_387# VPB phighvt w=1e+06u l=150000u
+  ad=7e+11p pd=5.4e+06u as=6.192e+11p ps=5.04e+06u
M1001 VPWR a_216_387# X VPB phighvt w=1.12e+06u l=150000u
+  ad=2.0608e+12p pd=1.474e+07u as=6.72e+11p ps=5.68e+06u
M1002 VPWR B1 a_216_387# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_125# A2 VGND VNB nshort w=640000u l=150000u
+  ad=7.744e+11p pd=7.54e+06u as=1.1573e+12p ps=1.034e+07u
M1004 VGND A2 a_27_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A1 a_116_387# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_216_387# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_216_387# VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1008 VGND a_216_387# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_216_387# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_125# B1 a_216_387# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1011 VGND A1 a_27_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_216_387# B1 VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_125# A1 VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_216_387# B1 a_27_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_216_387# A2 a_116_387# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_116_387# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_216_387# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_216_387# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_216_387# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

