* NGSPICE file created from sky130_fd_sc_ls__nand4_1.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nand4_1 A B C D VGND VNB VPB VPWR Y
M1000 a_181_74# D VGND VNB nshort w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.923e+11p ps=2.72e+06u
M1001 a_259_74# C a_181_74# VNB nshort w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1002 a_373_74# B a_259_74# VNB nshort w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1003 Y D VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=7.28e+11p pd=5.78e+06u as=1.232e+12p ps=8.92e+06u
M1004 Y B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR C Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A a_373_74# VNB nshort w=740000u l=150000u
+  ad=2.085e+11p pd=2.05e+06u as=0p ps=0u
.ends

