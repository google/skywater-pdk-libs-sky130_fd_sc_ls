* File: sky130_fd_sc_ls__and4_4.pxi.spice
* Created: Wed Sep  2 10:55:37 2020
* 
x_PM_SKY130_FD_SC_LS__AND4_4%A N_A_M1001_g N_A_c_136_n N_A_M1000_g N_A_M1003_g
+ N_A_c_137_n N_A_M1015_g A N_A_c_135_n PM_SKY130_FD_SC_LS__AND4_4%A
x_PM_SKY130_FD_SC_LS__AND4_4%B N_B_c_183_n N_B_M1017_g N_B_M1002_g N_B_c_185_n
+ N_B_c_186_n N_B_M1016_g N_B_c_192_n N_B_M1023_g N_B_c_188_n N_B_c_189_n B
+ N_B_c_190_n PM_SKY130_FD_SC_LS__AND4_4%B
x_PM_SKY130_FD_SC_LS__AND4_4%D N_D_c_247_n N_D_M1012_g N_D_c_252_n N_D_M1004_g
+ N_D_c_248_n N_D_M1018_g N_D_c_249_n N_D_c_250_n N_D_c_255_n N_D_M1010_g
+ N_D_c_251_n D PM_SKY130_FD_SC_LS__AND4_4%D
x_PM_SKY130_FD_SC_LS__AND4_4%C N_C_M1019_g N_C_M1006_g N_C_c_309_n N_C_c_310_n
+ N_C_M1020_g N_C_c_312_n N_C_c_313_n N_C_c_314_n N_C_M1009_g N_C_c_315_n
+ N_C_c_316_n N_C_c_321_n N_C_c_317_n C N_C_c_318_n PM_SKY130_FD_SC_LS__AND4_4%C
x_PM_SKY130_FD_SC_LS__AND4_4%A_116_392# N_A_116_392#_M1001_d
+ N_A_116_392#_M1017_d N_A_116_392#_M1015_d N_A_116_392#_M1006_d
+ N_A_116_392#_M1010_d N_A_116_392#_M1007_g N_A_116_392#_c_410_n
+ N_A_116_392#_M1005_g N_A_116_392#_M1013_g N_A_116_392#_c_411_n
+ N_A_116_392#_M1008_g N_A_116_392#_M1021_g N_A_116_392#_c_412_n
+ N_A_116_392#_M1011_g N_A_116_392#_M1022_g N_A_116_392#_c_413_n
+ N_A_116_392#_M1014_g N_A_116_392#_c_404_n N_A_116_392#_c_431_n
+ N_A_116_392#_c_405_n N_A_116_392#_c_415_n N_A_116_392#_c_416_n
+ N_A_116_392#_c_417_n N_A_116_392#_c_406_n N_A_116_392#_c_407_n
+ N_A_116_392#_c_456_n N_A_116_392#_c_420_n N_A_116_392#_c_465_n
+ N_A_116_392#_c_421_n N_A_116_392#_c_422_n N_A_116_392#_c_423_n
+ N_A_116_392#_c_408_n N_A_116_392#_c_538_p N_A_116_392#_c_458_n
+ N_A_116_392#_c_470_n N_A_116_392#_c_424_n N_A_116_392#_c_409_n
+ PM_SKY130_FD_SC_LS__AND4_4%A_116_392#
x_PM_SKY130_FD_SC_LS__AND4_4%VPWR N_VPWR_M1017_s N_VPWR_M1000_s N_VPWR_M1023_s
+ N_VPWR_M1004_s N_VPWR_M1009_s N_VPWR_M1008_s N_VPWR_M1014_s N_VPWR_c_594_n
+ N_VPWR_c_595_n N_VPWR_c_596_n N_VPWR_c_597_n N_VPWR_c_598_n N_VPWR_c_599_n
+ N_VPWR_c_600_n N_VPWR_c_601_n N_VPWR_c_602_n VPWR N_VPWR_c_603_n
+ N_VPWR_c_604_n N_VPWR_c_605_n N_VPWR_c_606_n N_VPWR_c_607_n N_VPWR_c_608_n
+ N_VPWR_c_609_n N_VPWR_c_610_n N_VPWR_c_611_n N_VPWR_c_612_n N_VPWR_c_613_n
+ N_VPWR_c_593_n PM_SKY130_FD_SC_LS__AND4_4%VPWR
x_PM_SKY130_FD_SC_LS__AND4_4%X N_X_M1007_s N_X_M1021_s N_X_M1005_d N_X_M1011_d
+ N_X_c_693_n N_X_c_702_n N_X_c_694_n N_X_c_695_n N_X_c_703_n N_X_c_704_n
+ N_X_c_696_n N_X_c_705_n N_X_c_706_n N_X_c_697_n N_X_c_698_n N_X_c_699_n
+ N_X_c_700_n N_X_c_743_n X PM_SKY130_FD_SC_LS__AND4_4%X
x_PM_SKY130_FD_SC_LS__AND4_4%A_32_119# N_A_32_119#_M1002_s N_A_32_119#_M1016_s
+ N_A_32_119#_M1020_s N_A_32_119#_c_771_n N_A_32_119#_c_772_n
+ N_A_32_119#_c_773_n N_A_32_119#_c_774_n N_A_32_119#_c_775_n
+ N_A_32_119#_c_776_n PM_SKY130_FD_SC_LS__AND4_4%A_32_119#
x_PM_SKY130_FD_SC_LS__AND4_4%A_119_119# N_A_119_119#_M1002_d
+ N_A_119_119#_M1003_s N_A_119_119#_c_820_n
+ PM_SKY130_FD_SC_LS__AND4_4%A_119_119#
x_PM_SKY130_FD_SC_LS__AND4_4%A_463_119# N_A_463_119#_M1019_d
+ N_A_463_119#_M1018_s N_A_463_119#_c_832_n N_A_463_119#_c_830_n
+ N_A_463_119#_c_831_n PM_SKY130_FD_SC_LS__AND4_4%A_463_119#
x_PM_SKY130_FD_SC_LS__AND4_4%VGND N_VGND_M1012_d N_VGND_M1007_d N_VGND_M1013_d
+ N_VGND_M1022_d N_VGND_c_859_n N_VGND_c_860_n N_VGND_c_861_n N_VGND_c_862_n
+ N_VGND_c_863_n N_VGND_c_864_n N_VGND_c_865_n VGND N_VGND_c_866_n
+ N_VGND_c_867_n N_VGND_c_868_n N_VGND_c_869_n N_VGND_c_870_n N_VGND_c_871_n
+ PM_SKY130_FD_SC_LS__AND4_4%VGND
cc_1 VNB N_A_M1001_g 0.0180096f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=0.915
cc_2 VNB N_A_M1003_g 0.0192586f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.915
cc_3 VNB A 9.7276e-19 $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_4 VNB N_A_c_135_n 0.025056f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.667
cc_5 VNB N_B_c_183_n 0.0254848f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.45
cc_6 VNB N_B_M1002_g 0.0418516f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.46
cc_7 VNB N_B_c_185_n 0.0851374f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.45
cc_8 VNB N_B_c_186_n 0.012806f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.915
cc_9 VNB N_B_M1016_g 0.0243266f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.46
cc_10 VNB N_B_c_188_n 0.0122598f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.615
cc_11 VNB N_B_c_189_n 0.010328f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.615
cc_12 VNB N_B_c_190_n 0.0094034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_D_c_247_n 0.0154852f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.45
cc_14 VNB N_D_c_248_n 0.0155847f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.46
cc_15 VNB N_D_c_249_n 0.00732157f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.915
cc_16 VNB N_D_c_250_n 0.047667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_D_c_251_n 0.00422422f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_18 VNB N_C_M1019_g 0.0232199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_C_c_309_n 0.0897065f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.915
cc_20 VNB N_C_c_310_n 0.00962308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_C_M1020_g 0.0300619f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.46
cc_22 VNB N_C_c_312_n 0.0387235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C_c_313_n 0.06444f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.667
cc_24 VNB N_C_c_314_n 0.0297301f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.615
cc_25 VNB N_C_c_315_n 0.0121624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_C_c_316_n 0.0105983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C_c_317_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_C_c_318_n 0.0103457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_116_392#_M1007_g 0.0234337f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.667
cc_30 VNB N_A_116_392#_M1013_g 0.0216149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_116_392#_M1021_g 0.0217861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_116_392#_M1022_g 0.0225815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_116_392#_c_404_n 0.00305189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_116_392#_c_405_n 0.00332779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_116_392#_c_406_n 0.00724257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_116_392#_c_407_n 0.00734814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_116_392#_c_408_n 0.00411229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_116_392#_c_409_n 0.109607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VPWR_c_593_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_X_c_693_n 0.00253173f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_41 VNB N_X_c_694_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.667
cc_42 VNB N_X_c_695_n 0.00208383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_X_c_696_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_X_c_697_n 0.0121765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_X_c_698_n 0.0127074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_X_c_699_n 2.15025e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_X_c_700_n 0.00279164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB X 0.0180896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_32_119#_c_771_n 0.0318742f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.885
cc_50 VNB N_A_32_119#_c_772_n 0.0219024f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.46
cc_51 VNB N_A_32_119#_c_773_n 0.00972966f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_52 VNB N_A_32_119#_c_774_n 0.00207833f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.667
cc_53 VNB N_A_32_119#_c_775_n 0.0143797f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.615
cc_54 VNB N_A_32_119#_c_776_n 0.0026989f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.615
cc_55 VNB N_A_463_119#_c_830_n 0.00261392f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.915
cc_56 VNB N_A_463_119#_c_831_n 0.00259991f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_57 VNB N_VGND_c_859_n 0.00881902f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_58 VNB N_VGND_c_860_n 0.0252934f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.667
cc_59 VNB N_VGND_c_861_n 0.00508214f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.667
cc_60 VNB N_VGND_c_862_n 0.0135817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_863_n 0.0232481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_864_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_865_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_866_n 0.0720971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_867_n 0.0353709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_868_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_869_n 0.0043699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_870_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_871_n 0.352482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VPB N_A_c_136_n 0.0148981f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.885
cc_71 VPB N_A_c_137_n 0.0153402f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.885
cc_72 VPB A 0.00235587f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_73 VPB N_A_c_135_n 0.0316581f $X=-0.19 $Y=1.66 $X2=1.38 $Y2=1.667
cc_74 VPB N_B_c_183_n 0.0443003f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.45
cc_75 VPB N_B_c_192_n 0.0276468f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_B_c_189_n 0.00170971f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=1.615
cc_77 VPB N_B_c_190_n 0.0054581f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_D_c_252_n 0.018112f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_D_c_249_n 0.0103289f $X=-0.19 $Y=1.66 $X2=1.38 $Y2=0.915
cc_80 VPB N_D_c_250_n 0.0290192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_D_c_255_n 0.0198f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.885
cc_82 VPB N_D_c_251_n 0.0123035f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_83 VPB D 0.00304223f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.667
cc_84 VPB N_C_c_314_n 0.0350822f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=1.615
cc_85 VPB N_C_c_316_n 0.00336987f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_C_c_321_n 0.0294232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_C_c_318_n 0.00386538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_116_392#_c_410_n 0.0166603f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=1.615
cc_89 VPB N_A_116_392#_c_411_n 0.0156114f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_116_392#_c_412_n 0.0147069f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_116_392#_c_413_n 0.0173993f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_116_392#_c_404_n 0.00702866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_116_392#_c_415_n 0.00442853f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_116_392#_c_416_n 0.00310079f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_116_392#_c_417_n 0.00181251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_116_392#_c_406_n 0.00420469f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_116_392#_c_407_n 7.78204e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_116_392#_c_420_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_116_392#_c_421_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_116_392#_c_422_n 0.00261914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_116_392#_c_423_n 0.00135055f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_116_392#_c_424_n 0.00796949f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_116_392#_c_409_n 0.0294634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_594_n 0.0112292f $X=-0.19 $Y=1.66 $X2=1.38 $Y2=1.667
cc_105 VPB N_VPWR_c_595_n 0.051952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_596_n 0.00270216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_597_n 0.00799067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_598_n 0.00931414f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_599_n 0.00907555f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_600_n 0.00510801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_601_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_602_n 0.059413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_603_n 0.019508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_604_n 0.016911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_605_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_606_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_607_n 0.0215588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_608_n 0.0175706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_609_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_610_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_611_n 0.0135466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_612_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_613_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_593_n 0.0903849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_X_c_702_n 0.002914f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=1.667
cc_126 VPB N_X_c_703_n 0.0023626f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_X_c_704_n 0.00230344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_X_c_705_n 0.00132334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_X_c_706_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 N_A_c_136_n N_B_c_183_n 0.0328919f $X=0.955 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_131 N_A_c_135_n N_B_c_183_n 0.0227344f $X=1.38 $Y=1.667 $X2=-0.19 $Y2=-0.245
cc_132 N_A_M1001_g N_B_M1002_g 0.0227344f $X=0.95 $Y=0.915 $X2=0 $Y2=0
cc_133 N_A_M1001_g N_B_c_185_n 0.00880809f $X=0.95 $Y=0.915 $X2=0 $Y2=0
cc_134 N_A_M1003_g N_B_c_185_n 0.00880809f $X=1.38 $Y=0.915 $X2=0 $Y2=0
cc_135 N_A_M1003_g N_B_M1016_g 0.0291179f $X=1.38 $Y=0.915 $X2=0 $Y2=0
cc_136 N_A_c_137_n N_B_c_192_n 0.00675566f $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_137 N_A_c_135_n N_B_c_188_n 6.11939e-19 $X=1.38 $Y=1.667 $X2=0 $Y2=0
cc_138 A N_B_c_189_n 8.36911e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A_c_135_n N_B_c_189_n 0.0184422f $X=1.38 $Y=1.667 $X2=0 $Y2=0
cc_140 N_A_c_135_n N_B_c_190_n 2.96224e-19 $X=1.38 $Y=1.667 $X2=0 $Y2=0
cc_141 N_A_M1001_g N_A_116_392#_c_404_n 0.00461704f $X=0.95 $Y=0.915 $X2=0 $Y2=0
cc_142 N_A_c_136_n N_A_116_392#_c_404_n 0.0024644f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_143 N_A_M1003_g N_A_116_392#_c_404_n 9.34592e-19 $X=1.38 $Y=0.915 $X2=0 $Y2=0
cc_144 A N_A_116_392#_c_404_n 0.0235661f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_145 N_A_c_135_n N_A_116_392#_c_404_n 0.0106678f $X=1.38 $Y=1.667 $X2=0 $Y2=0
cc_146 N_A_M1001_g N_A_116_392#_c_431_n 0.00245644f $X=0.95 $Y=0.915 $X2=0 $Y2=0
cc_147 N_A_M1001_g N_A_116_392#_c_405_n 0.0113714f $X=0.95 $Y=0.915 $X2=0 $Y2=0
cc_148 N_A_M1003_g N_A_116_392#_c_405_n 0.00556676f $X=1.38 $Y=0.915 $X2=0 $Y2=0
cc_149 A N_A_116_392#_c_405_n 0.0187733f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A_c_135_n N_A_116_392#_c_405_n 7.06359e-19 $X=1.38 $Y=1.667 $X2=0 $Y2=0
cc_151 N_A_c_136_n N_A_116_392#_c_415_n 0.0199437f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_152 N_A_c_137_n N_A_116_392#_c_415_n 0.0193547f $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_153 A N_A_116_392#_c_415_n 0.025582f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_154 N_A_c_135_n N_A_116_392#_c_415_n 0.00442963f $X=1.38 $Y=1.667 $X2=0 $Y2=0
cc_155 N_A_c_137_n N_A_116_392#_c_416_n 8.2201e-19 $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_156 A N_A_116_392#_c_416_n 7.13846e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A_c_135_n N_A_116_392#_c_416_n 0.00144931f $X=1.38 $Y=1.667 $X2=0 $Y2=0
cc_158 N_A_c_137_n N_A_116_392#_c_417_n 0.00518098f $X=1.405 $Y=1.885 $X2=0
+ $Y2=0
cc_159 A N_A_116_392#_c_407_n 0.0143347f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_160 N_A_c_135_n N_A_116_392#_c_407_n 0.00162846f $X=1.38 $Y=1.667 $X2=0 $Y2=0
cc_161 N_A_c_136_n N_VPWR_c_596_n 0.0145292f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_162 N_A_c_137_n N_VPWR_c_596_n 0.0100586f $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_163 N_A_c_137_n N_VPWR_c_597_n 6.39103e-19 $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_164 N_A_c_136_n N_VPWR_c_603_n 0.00413917f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_165 N_A_c_137_n N_VPWR_c_604_n 0.00413917f $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_166 N_A_c_136_n N_VPWR_c_593_n 0.0081781f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_167 N_A_c_137_n N_VPWR_c_593_n 0.00817943f $X=1.405 $Y=1.885 $X2=0 $Y2=0
cc_168 N_A_M1001_g N_A_32_119#_c_772_n 0.00361508f $X=0.95 $Y=0.915 $X2=0 $Y2=0
cc_169 N_A_M1003_g N_A_32_119#_c_772_n 0.00361508f $X=1.38 $Y=0.915 $X2=0 $Y2=0
cc_170 N_A_M1001_g N_A_119_119#_c_820_n 0.00855819f $X=0.95 $Y=0.915 $X2=0 $Y2=0
cc_171 N_A_M1003_g N_A_119_119#_c_820_n 0.0113852f $X=1.38 $Y=0.915 $X2=0 $Y2=0
cc_172 A N_A_119_119#_c_820_n 0.00146023f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_173 N_B_M1016_g N_C_M1019_g 0.0123703f $X=1.81 $Y=0.915 $X2=0 $Y2=0
cc_174 N_B_c_185_n N_C_c_310_n 0.0123703f $X=1.735 $Y=0.18 $X2=0 $Y2=0
cc_175 N_B_c_188_n N_C_c_315_n 0.00937754f $X=1.832 $Y=1.46 $X2=0 $Y2=0
cc_176 N_B_c_192_n N_C_c_316_n 0.00837718f $X=1.87 $Y=1.885 $X2=0 $Y2=0
cc_177 N_B_c_189_n N_C_c_316_n 0.010557f $X=1.87 $Y=1.7 $X2=0 $Y2=0
cc_178 N_B_c_192_n N_C_c_321_n 0.0187009f $X=1.87 $Y=1.885 $X2=0 $Y2=0
cc_179 N_B_c_183_n N_A_116_392#_c_404_n 0.00650457f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_180 N_B_M1002_g N_A_116_392#_c_404_n 0.00885625f $X=0.52 $Y=0.915 $X2=0 $Y2=0
cc_181 N_B_c_190_n N_A_116_392#_c_404_n 0.0252572f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_182 N_B_M1002_g N_A_116_392#_c_431_n 0.0023738f $X=0.52 $Y=0.915 $X2=0 $Y2=0
cc_183 N_B_M1016_g N_A_116_392#_c_405_n 7.51685e-19 $X=1.81 $Y=0.915 $X2=0 $Y2=0
cc_184 N_B_c_192_n N_A_116_392#_c_416_n 0.00416122f $X=1.87 $Y=1.885 $X2=0 $Y2=0
cc_185 N_B_c_192_n N_A_116_392#_c_417_n 0.0024225f $X=1.87 $Y=1.885 $X2=0 $Y2=0
cc_186 N_B_c_192_n N_A_116_392#_c_406_n 0.00997747f $X=1.87 $Y=1.885 $X2=0 $Y2=0
cc_187 N_B_c_188_n N_A_116_392#_c_406_n 0.00192947f $X=1.832 $Y=1.46 $X2=0 $Y2=0
cc_188 N_B_c_189_n N_A_116_392#_c_406_n 0.00994393f $X=1.87 $Y=1.7 $X2=0 $Y2=0
cc_189 N_B_c_192_n N_A_116_392#_c_456_n 7.68141e-19 $X=1.87 $Y=1.885 $X2=0 $Y2=0
cc_190 N_B_c_192_n N_A_116_392#_c_420_n 2.02005e-19 $X=1.87 $Y=1.885 $X2=0 $Y2=0
cc_191 N_B_c_192_n N_A_116_392#_c_458_n 0.00131763f $X=1.87 $Y=1.885 $X2=0 $Y2=0
cc_192 N_B_c_183_n N_VPWR_c_595_n 0.0080553f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_193 N_B_c_190_n N_VPWR_c_595_n 0.0230778f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_194 N_B_c_183_n N_VPWR_c_596_n 0.0020477f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_195 N_B_c_192_n N_VPWR_c_596_n 5.07366e-19 $X=1.87 $Y=1.885 $X2=0 $Y2=0
cc_196 N_B_c_192_n N_VPWR_c_597_n 0.0151602f $X=1.87 $Y=1.885 $X2=0 $Y2=0
cc_197 N_B_c_183_n N_VPWR_c_603_n 0.00461464f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_198 N_B_c_192_n N_VPWR_c_604_n 0.00413917f $X=1.87 $Y=1.885 $X2=0 $Y2=0
cc_199 N_B_c_183_n N_VPWR_c_593_n 0.00911857f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_200 N_B_c_192_n N_VPWR_c_593_n 0.00817943f $X=1.87 $Y=1.885 $X2=0 $Y2=0
cc_201 N_B_c_183_n N_A_32_119#_c_771_n 0.00388745f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_202 N_B_M1002_g N_A_32_119#_c_771_n 0.00491408f $X=0.52 $Y=0.915 $X2=0 $Y2=0
cc_203 N_B_c_190_n N_A_32_119#_c_771_n 0.0191995f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_204 N_B_M1002_g N_A_32_119#_c_772_n 0.0171399f $X=0.52 $Y=0.915 $X2=0 $Y2=0
cc_205 N_B_c_185_n N_A_32_119#_c_772_n 0.0170084f $X=1.735 $Y=0.18 $X2=0 $Y2=0
cc_206 N_B_M1016_g N_A_32_119#_c_772_n 0.0152701f $X=1.81 $Y=0.915 $X2=0 $Y2=0
cc_207 N_B_M1016_g N_A_32_119#_c_774_n 0.00258587f $X=1.81 $Y=0.915 $X2=0 $Y2=0
cc_208 N_B_M1016_g N_A_32_119#_c_776_n 0.00174203f $X=1.81 $Y=0.915 $X2=0 $Y2=0
cc_209 N_B_M1002_g N_A_119_119#_c_820_n 0.00334426f $X=0.52 $Y=0.915 $X2=0 $Y2=0
cc_210 N_B_M1016_g N_A_119_119#_c_820_n 0.00320291f $X=1.81 $Y=0.915 $X2=0 $Y2=0
cc_211 N_B_c_186_n N_VGND_c_866_n 0.0319108f $X=0.595 $Y=0.18 $X2=0 $Y2=0
cc_212 N_B_c_185_n N_VGND_c_871_n 0.0315727f $X=1.735 $Y=0.18 $X2=0 $Y2=0
cc_213 N_B_c_186_n N_VGND_c_871_n 0.00563808f $X=0.595 $Y=0.18 $X2=0 $Y2=0
cc_214 N_D_c_247_n N_C_M1019_g 0.0214926f $X=2.67 $Y=1.345 $X2=0 $Y2=0
cc_215 N_D_c_247_n N_C_c_309_n 0.00994861f $X=2.67 $Y=1.345 $X2=0 $Y2=0
cc_216 N_D_c_248_n N_C_c_309_n 0.00992356f $X=3.26 $Y=1.345 $X2=0 $Y2=0
cc_217 N_D_c_248_n N_C_M1020_g 0.0258115f $X=3.26 $Y=1.345 $X2=0 $Y2=0
cc_218 N_D_c_251_n N_C_M1020_g 0.00768122f $X=3.705 $Y=1.725 $X2=0 $Y2=0
cc_219 N_D_c_250_n N_C_c_314_n 0.00356952f $X=3.335 $Y=1.725 $X2=0 $Y2=0
cc_220 N_D_c_255_n N_C_c_314_n 0.0203274f $X=3.705 $Y=1.885 $X2=0 $Y2=0
cc_221 N_D_c_251_n N_C_c_314_n 0.0103605f $X=3.705 $Y=1.725 $X2=0 $Y2=0
cc_222 N_D_c_247_n N_C_c_315_n 0.00684318f $X=2.67 $Y=1.345 $X2=0 $Y2=0
cc_223 N_D_c_250_n N_C_c_316_n 0.0159302f $X=3.335 $Y=1.725 $X2=0 $Y2=0
cc_224 D N_C_c_316_n 6.03167e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_225 N_D_c_252_n N_C_c_321_n 0.00813438f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_226 N_D_c_250_n N_C_c_321_n 0.00712163f $X=3.335 $Y=1.725 $X2=0 $Y2=0
cc_227 N_D_c_250_n N_C_c_318_n 0.00498553f $X=3.335 $Y=1.725 $X2=0 $Y2=0
cc_228 N_D_c_251_n N_C_c_318_n 0.00332603f $X=3.705 $Y=1.725 $X2=0 $Y2=0
cc_229 N_D_c_250_n N_A_116_392#_c_406_n 0.0101364f $X=3.335 $Y=1.725 $X2=0 $Y2=0
cc_230 D N_A_116_392#_c_406_n 0.0135702f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_231 N_D_c_252_n N_A_116_392#_c_456_n 0.00443864f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_232 N_D_c_250_n N_A_116_392#_c_456_n 0.00592418f $X=3.335 $Y=1.725 $X2=0
+ $Y2=0
cc_233 D N_A_116_392#_c_456_n 0.00221382f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_234 N_D_c_252_n N_A_116_392#_c_420_n 0.0142372f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_235 N_D_c_252_n N_A_116_392#_c_465_n 0.0158416f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_236 N_D_c_250_n N_A_116_392#_c_465_n 0.0110137f $X=3.335 $Y=1.725 $X2=0 $Y2=0
cc_237 N_D_c_255_n N_A_116_392#_c_465_n 0.0182672f $X=3.705 $Y=1.885 $X2=0 $Y2=0
cc_238 D N_A_116_392#_c_465_n 0.0235751f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_239 N_D_c_255_n N_A_116_392#_c_421_n 0.00453404f $X=3.705 $Y=1.885 $X2=0
+ $Y2=0
cc_240 N_D_c_252_n N_A_116_392#_c_470_n 2.24111e-19 $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_241 N_D_c_255_n N_A_116_392#_c_424_n 3.58983e-19 $X=3.705 $Y=1.885 $X2=0
+ $Y2=0
cc_242 N_D_c_252_n N_VPWR_c_598_n 0.00399486f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_243 N_D_c_255_n N_VPWR_c_598_n 0.0120401f $X=3.705 $Y=1.885 $X2=0 $Y2=0
cc_244 N_D_c_252_n N_VPWR_c_605_n 0.00445602f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_245 N_D_c_255_n N_VPWR_c_606_n 0.00413917f $X=3.705 $Y=1.885 $X2=0 $Y2=0
cc_246 N_D_c_252_n N_VPWR_c_593_n 0.00861803f $X=2.82 $Y=1.885 $X2=0 $Y2=0
cc_247 N_D_c_255_n N_VPWR_c_593_n 0.00818241f $X=3.705 $Y=1.885 $X2=0 $Y2=0
cc_248 N_D_c_247_n N_A_32_119#_c_775_n 0.011277f $X=2.67 $Y=1.345 $X2=0 $Y2=0
cc_249 N_D_c_248_n N_A_32_119#_c_775_n 0.0129724f $X=3.26 $Y=1.345 $X2=0 $Y2=0
cc_250 N_D_c_249_n N_A_32_119#_c_775_n 0.00533033f $X=3.615 $Y=1.725 $X2=0 $Y2=0
cc_251 N_D_c_250_n N_A_32_119#_c_775_n 0.00799205f $X=3.335 $Y=1.725 $X2=0 $Y2=0
cc_252 N_D_c_251_n N_A_32_119#_c_775_n 0.00138333f $X=3.705 $Y=1.725 $X2=0 $Y2=0
cc_253 D N_A_32_119#_c_775_n 0.0244958f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_254 N_D_c_247_n N_A_463_119#_c_832_n 0.00814407f $X=2.67 $Y=1.345 $X2=0 $Y2=0
cc_255 N_D_c_248_n N_A_463_119#_c_832_n 0.00722037f $X=3.26 $Y=1.345 $X2=0 $Y2=0
cc_256 N_D_c_247_n N_A_463_119#_c_830_n 0.00575669f $X=2.67 $Y=1.345 $X2=0 $Y2=0
cc_257 N_D_c_248_n N_A_463_119#_c_830_n 8.58549e-19 $X=3.26 $Y=1.345 $X2=0 $Y2=0
cc_258 N_D_c_247_n N_A_463_119#_c_831_n 7.89916e-19 $X=2.67 $Y=1.345 $X2=0 $Y2=0
cc_259 N_D_c_248_n N_A_463_119#_c_831_n 0.00606088f $X=3.26 $Y=1.345 $X2=0 $Y2=0
cc_260 N_D_c_247_n N_VGND_c_859_n 0.00354211f $X=2.67 $Y=1.345 $X2=0 $Y2=0
cc_261 N_D_c_248_n N_VGND_c_859_n 0.00353848f $X=3.26 $Y=1.345 $X2=0 $Y2=0
cc_262 N_D_c_247_n N_VGND_c_871_n 9.39239e-19 $X=2.67 $Y=1.345 $X2=0 $Y2=0
cc_263 N_D_c_248_n N_VGND_c_871_n 9.39239e-19 $X=3.26 $Y=1.345 $X2=0 $Y2=0
cc_264 N_C_c_312_n N_A_116_392#_M1007_g 0.00925508f $X=4.125 $Y=0.18 $X2=0 $Y2=0
cc_265 N_C_c_314_n N_A_116_392#_c_410_n 0.0294753f $X=4.205 $Y=1.885 $X2=0 $Y2=0
cc_266 N_C_c_315_n N_A_116_392#_c_406_n 0.00201969f $X=2.275 $Y=1.46 $X2=0 $Y2=0
cc_267 N_C_c_316_n N_A_116_392#_c_406_n 0.00790199f $X=2.347 $Y=1.735 $X2=0
+ $Y2=0
cc_268 N_C_c_321_n N_A_116_392#_c_406_n 0.0102621f $X=2.347 $Y=1.885 $X2=0 $Y2=0
cc_269 N_C_c_321_n N_A_116_392#_c_456_n 0.00614378f $X=2.347 $Y=1.885 $X2=0
+ $Y2=0
cc_270 N_C_c_321_n N_A_116_392#_c_420_n 0.0083713f $X=2.347 $Y=1.885 $X2=0 $Y2=0
cc_271 N_C_M1020_g N_A_116_392#_c_465_n 3.83636e-19 $X=3.69 $Y=0.915 $X2=0 $Y2=0
cc_272 N_C_c_314_n N_A_116_392#_c_421_n 0.00990613f $X=4.205 $Y=1.885 $X2=0
+ $Y2=0
cc_273 N_C_c_314_n N_A_116_392#_c_422_n 0.0132811f $X=4.205 $Y=1.885 $X2=0 $Y2=0
cc_274 N_C_c_318_n N_A_116_392#_c_422_n 0.0166511f $X=4.2 $Y=1.51 $X2=0 $Y2=0
cc_275 N_C_c_314_n N_A_116_392#_c_423_n 0.00398618f $X=4.205 $Y=1.885 $X2=0
+ $Y2=0
cc_276 N_C_c_318_n N_A_116_392#_c_423_n 0.0118112f $X=4.2 $Y=1.51 $X2=0 $Y2=0
cc_277 N_C_c_313_n N_A_116_392#_c_408_n 0.00115834f $X=4.2 $Y=1.345 $X2=0 $Y2=0
cc_278 N_C_c_314_n N_A_116_392#_c_408_n 0.00211809f $X=4.205 $Y=1.885 $X2=0
+ $Y2=0
cc_279 N_C_c_318_n N_A_116_392#_c_408_n 0.0242915f $X=4.2 $Y=1.51 $X2=0 $Y2=0
cc_280 N_C_c_321_n N_A_116_392#_c_470_n 0.00162804f $X=2.347 $Y=1.885 $X2=0
+ $Y2=0
cc_281 N_C_c_314_n N_A_116_392#_c_424_n 0.00190723f $X=4.205 $Y=1.885 $X2=0
+ $Y2=0
cc_282 N_C_c_318_n N_A_116_392#_c_424_n 0.0146704f $X=4.2 $Y=1.51 $X2=0 $Y2=0
cc_283 N_C_c_313_n N_A_116_392#_c_409_n 0.00925508f $X=4.2 $Y=1.345 $X2=0 $Y2=0
cc_284 N_C_c_314_n N_A_116_392#_c_409_n 0.0151065f $X=4.205 $Y=1.885 $X2=0 $Y2=0
cc_285 N_C_c_318_n N_A_116_392#_c_409_n 5.84105e-19 $X=4.2 $Y=1.51 $X2=0 $Y2=0
cc_286 N_C_c_321_n N_VPWR_c_597_n 0.00815893f $X=2.347 $Y=1.885 $X2=0 $Y2=0
cc_287 N_C_c_314_n N_VPWR_c_598_n 4.9921e-19 $X=4.205 $Y=1.885 $X2=0 $Y2=0
cc_288 N_C_c_314_n N_VPWR_c_599_n 0.00608458f $X=4.205 $Y=1.885 $X2=0 $Y2=0
cc_289 N_C_c_321_n N_VPWR_c_605_n 0.00445602f $X=2.347 $Y=1.885 $X2=0 $Y2=0
cc_290 N_C_c_314_n N_VPWR_c_606_n 0.00445602f $X=4.205 $Y=1.885 $X2=0 $Y2=0
cc_291 N_C_c_314_n N_VPWR_c_593_n 0.00858414f $X=4.205 $Y=1.885 $X2=0 $Y2=0
cc_292 N_C_c_321_n N_VPWR_c_593_n 0.00857515f $X=2.347 $Y=1.885 $X2=0 $Y2=0
cc_293 N_C_M1019_g N_A_32_119#_c_772_n 0.0053794f $X=2.24 $Y=0.915 $X2=0 $Y2=0
cc_294 N_C_M1019_g N_A_32_119#_c_774_n 0.00226802f $X=2.24 $Y=0.915 $X2=0 $Y2=0
cc_295 N_C_M1019_g N_A_32_119#_c_775_n 0.0131304f $X=2.24 $Y=0.915 $X2=0 $Y2=0
cc_296 N_C_M1020_g N_A_32_119#_c_775_n 0.0169435f $X=3.69 $Y=0.915 $X2=0 $Y2=0
cc_297 N_C_c_313_n N_A_32_119#_c_775_n 0.00458254f $X=4.2 $Y=1.345 $X2=0 $Y2=0
cc_298 N_C_c_314_n N_A_32_119#_c_775_n 2.4826e-19 $X=4.205 $Y=1.885 $X2=0 $Y2=0
cc_299 N_C_c_315_n N_A_32_119#_c_775_n 0.00237026f $X=2.275 $Y=1.46 $X2=0 $Y2=0
cc_300 N_C_c_321_n N_A_32_119#_c_775_n 3.74671e-19 $X=2.347 $Y=1.885 $X2=0 $Y2=0
cc_301 N_C_c_318_n N_A_32_119#_c_775_n 0.00707047f $X=4.2 $Y=1.51 $X2=0 $Y2=0
cc_302 N_C_c_309_n N_A_463_119#_c_832_n 0.00192114f $X=3.615 $Y=0.18 $X2=0 $Y2=0
cc_303 N_C_M1019_g N_A_463_119#_c_830_n 0.0050314f $X=2.24 $Y=0.915 $X2=0 $Y2=0
cc_304 N_C_c_309_n N_A_463_119#_c_830_n 0.00377905f $X=3.615 $Y=0.18 $X2=0 $Y2=0
cc_305 N_C_c_309_n N_A_463_119#_c_831_n 0.00378414f $X=3.615 $Y=0.18 $X2=0 $Y2=0
cc_306 N_C_M1020_g N_A_463_119#_c_831_n 0.0096002f $X=3.69 $Y=0.915 $X2=0 $Y2=0
cc_307 N_C_c_313_n N_A_463_119#_c_831_n 0.00117577f $X=4.2 $Y=1.345 $X2=0 $Y2=0
cc_308 N_C_M1019_g N_VGND_c_859_n 0.00579091f $X=2.24 $Y=0.915 $X2=0 $Y2=0
cc_309 N_C_c_309_n N_VGND_c_859_n 0.025075f $X=3.615 $Y=0.18 $X2=0 $Y2=0
cc_310 N_C_M1020_g N_VGND_c_859_n 0.00579091f $X=3.69 $Y=0.915 $X2=0 $Y2=0
cc_311 N_C_c_312_n N_VGND_c_860_n 0.0281566f $X=4.125 $Y=0.18 $X2=0 $Y2=0
cc_312 N_C_c_314_n N_VGND_c_860_n 2.53681e-19 $X=4.205 $Y=1.885 $X2=0 $Y2=0
cc_313 N_C_c_318_n N_VGND_c_860_n 0.00238772f $X=4.2 $Y=1.51 $X2=0 $Y2=0
cc_314 N_C_c_310_n N_VGND_c_866_n 0.0195624f $X=2.315 $Y=0.18 $X2=0 $Y2=0
cc_315 N_C_c_309_n N_VGND_c_867_n 0.0386165f $X=3.615 $Y=0.18 $X2=0 $Y2=0
cc_316 N_C_c_309_n N_VGND_c_871_n 0.0259073f $X=3.615 $Y=0.18 $X2=0 $Y2=0
cc_317 N_C_c_310_n N_VGND_c_871_n 0.00935062f $X=2.315 $Y=0.18 $X2=0 $Y2=0
cc_318 N_C_c_312_n N_VGND_c_871_n 0.0322624f $X=4.125 $Y=0.18 $X2=0 $Y2=0
cc_319 N_C_c_317_n N_VGND_c_871_n 0.00841737f $X=3.69 $Y=0.18 $X2=0 $Y2=0
cc_320 N_A_116_392#_c_415_n N_VPWR_M1000_s 0.00201f $X=1.56 $Y=2.095 $X2=0 $Y2=0
cc_321 N_A_116_392#_c_465_n N_VPWR_M1004_s 0.0171089f $X=3.815 $Y=2.055 $X2=0
+ $Y2=0
cc_322 N_A_116_392#_c_422_n N_VPWR_M1009_s 0.007784f $X=4.535 $Y=2.035 $X2=0
+ $Y2=0
cc_323 N_A_116_392#_c_423_n N_VPWR_M1009_s 0.00134158f $X=4.62 $Y=1.95 $X2=0
+ $Y2=0
cc_324 N_A_116_392#_c_404_n N_VPWR_c_595_n 0.0125828f $X=0.805 $Y=1.95 $X2=0
+ $Y2=0
cc_325 N_A_116_392#_c_415_n N_VPWR_c_596_n 0.0178275f $X=1.56 $Y=2.095 $X2=0
+ $Y2=0
cc_326 N_A_116_392#_c_417_n N_VPWR_c_596_n 0.0351505f $X=1.645 $Y=2.46 $X2=0
+ $Y2=0
cc_327 N_A_116_392#_c_416_n N_VPWR_c_597_n 6.31475e-19 $X=1.645 $Y=1.95 $X2=0
+ $Y2=0
cc_328 N_A_116_392#_c_417_n N_VPWR_c_597_n 0.0481964f $X=1.645 $Y=2.46 $X2=0
+ $Y2=0
cc_329 N_A_116_392#_c_406_n N_VPWR_c_597_n 0.0274392f $X=2.43 $Y=1.685 $X2=0
+ $Y2=0
cc_330 N_A_116_392#_c_456_n N_VPWR_c_597_n 0.00187864f $X=2.595 $Y=1.97 $X2=0
+ $Y2=0
cc_331 N_A_116_392#_c_420_n N_VPWR_c_597_n 0.0322718f $X=2.595 $Y=2.815 $X2=0
+ $Y2=0
cc_332 N_A_116_392#_c_458_n N_VPWR_c_597_n 0.0211398f $X=1.645 $Y=2.105 $X2=0
+ $Y2=0
cc_333 N_A_116_392#_c_420_n N_VPWR_c_598_n 0.0260284f $X=2.595 $Y=2.815 $X2=0
+ $Y2=0
cc_334 N_A_116_392#_c_465_n N_VPWR_c_598_n 0.051548f $X=3.815 $Y=2.055 $X2=0
+ $Y2=0
cc_335 N_A_116_392#_c_421_n N_VPWR_c_598_n 0.0290836f $X=3.98 $Y=2.815 $X2=0
+ $Y2=0
cc_336 N_A_116_392#_c_410_n N_VPWR_c_599_n 0.00736481f $X=4.765 $Y=1.765 $X2=0
+ $Y2=0
cc_337 N_A_116_392#_c_421_n N_VPWR_c_599_n 0.0266809f $X=3.98 $Y=2.815 $X2=0
+ $Y2=0
cc_338 N_A_116_392#_c_422_n N_VPWR_c_599_n 0.0248633f $X=4.535 $Y=2.035 $X2=0
+ $Y2=0
cc_339 N_A_116_392#_c_411_n N_VPWR_c_600_n 0.00630489f $X=5.265 $Y=1.765 $X2=0
+ $Y2=0
cc_340 N_A_116_392#_c_412_n N_VPWR_c_600_n 0.0134288f $X=5.715 $Y=1.765 $X2=0
+ $Y2=0
cc_341 N_A_116_392#_c_413_n N_VPWR_c_600_n 6.21454e-19 $X=6.165 $Y=1.765 $X2=0
+ $Y2=0
cc_342 N_A_116_392#_c_413_n N_VPWR_c_602_n 0.0260839f $X=6.165 $Y=1.765 $X2=0
+ $Y2=0
cc_343 N_A_116_392#_c_417_n N_VPWR_c_604_n 0.00749631f $X=1.645 $Y=2.46 $X2=0
+ $Y2=0
cc_344 N_A_116_392#_c_420_n N_VPWR_c_605_n 0.014552f $X=2.595 $Y=2.815 $X2=0
+ $Y2=0
cc_345 N_A_116_392#_c_421_n N_VPWR_c_606_n 0.0145938f $X=3.98 $Y=2.815 $X2=0
+ $Y2=0
cc_346 N_A_116_392#_c_410_n N_VPWR_c_607_n 0.00461464f $X=4.765 $Y=1.765 $X2=0
+ $Y2=0
cc_347 N_A_116_392#_c_411_n N_VPWR_c_607_n 0.00445602f $X=5.265 $Y=1.765 $X2=0
+ $Y2=0
cc_348 N_A_116_392#_c_412_n N_VPWR_c_608_n 0.00413917f $X=5.715 $Y=1.765 $X2=0
+ $Y2=0
cc_349 N_A_116_392#_c_413_n N_VPWR_c_608_n 0.00445602f $X=6.165 $Y=1.765 $X2=0
+ $Y2=0
cc_350 N_A_116_392#_c_410_n N_VPWR_c_593_n 0.00909946f $X=4.765 $Y=1.765 $X2=0
+ $Y2=0
cc_351 N_A_116_392#_c_411_n N_VPWR_c_593_n 0.0085805f $X=5.265 $Y=1.765 $X2=0
+ $Y2=0
cc_352 N_A_116_392#_c_412_n N_VPWR_c_593_n 0.00817726f $X=5.715 $Y=1.765 $X2=0
+ $Y2=0
cc_353 N_A_116_392#_c_413_n N_VPWR_c_593_n 0.00860566f $X=6.165 $Y=1.765 $X2=0
+ $Y2=0
cc_354 N_A_116_392#_c_417_n N_VPWR_c_593_n 0.0062048f $X=1.645 $Y=2.46 $X2=0
+ $Y2=0
cc_355 N_A_116_392#_c_420_n N_VPWR_c_593_n 0.0119791f $X=2.595 $Y=2.815 $X2=0
+ $Y2=0
cc_356 N_A_116_392#_c_421_n N_VPWR_c_593_n 0.0120466f $X=3.98 $Y=2.815 $X2=0
+ $Y2=0
cc_357 N_A_116_392#_M1007_g N_X_c_693_n 4.72738e-19 $X=4.75 $Y=0.74 $X2=0 $Y2=0
cc_358 N_A_116_392#_M1013_g N_X_c_693_n 4.28846e-19 $X=5.21 $Y=0.74 $X2=0 $Y2=0
cc_359 N_A_116_392#_c_410_n N_X_c_702_n 0.00545879f $X=4.765 $Y=1.765 $X2=0
+ $Y2=0
cc_360 N_A_116_392#_c_411_n N_X_c_702_n 0.0126706f $X=5.265 $Y=1.765 $X2=0 $Y2=0
cc_361 N_A_116_392#_c_412_n N_X_c_702_n 7.68526e-19 $X=5.715 $Y=1.765 $X2=0
+ $Y2=0
cc_362 N_A_116_392#_M1013_g N_X_c_694_n 0.0128692f $X=5.21 $Y=0.74 $X2=0 $Y2=0
cc_363 N_A_116_392#_M1021_g N_X_c_694_n 0.0126341f $X=5.71 $Y=0.74 $X2=0 $Y2=0
cc_364 N_A_116_392#_c_538_p N_X_c_694_n 0.0446871f $X=5.52 $Y=1.465 $X2=0 $Y2=0
cc_365 N_A_116_392#_c_409_n N_X_c_694_n 0.00381149f $X=6.14 $Y=1.532 $X2=0 $Y2=0
cc_366 N_A_116_392#_c_538_p N_X_c_695_n 0.0210857f $X=5.52 $Y=1.465 $X2=0 $Y2=0
cc_367 N_A_116_392#_c_409_n N_X_c_695_n 0.00302844f $X=6.14 $Y=1.532 $X2=0 $Y2=0
cc_368 N_A_116_392#_c_411_n N_X_c_703_n 0.0120074f $X=5.265 $Y=1.765 $X2=0 $Y2=0
cc_369 N_A_116_392#_c_412_n N_X_c_703_n 0.0147308f $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_370 N_A_116_392#_c_538_p N_X_c_703_n 0.035367f $X=5.52 $Y=1.465 $X2=0 $Y2=0
cc_371 N_A_116_392#_c_409_n N_X_c_703_n 0.00948886f $X=6.14 $Y=1.532 $X2=0 $Y2=0
cc_372 N_A_116_392#_c_410_n N_X_c_704_n 0.00106358f $X=4.765 $Y=1.765 $X2=0
+ $Y2=0
cc_373 N_A_116_392#_c_411_n N_X_c_704_n 9.20137e-19 $X=5.265 $Y=1.765 $X2=0
+ $Y2=0
cc_374 N_A_116_392#_c_423_n N_X_c_704_n 0.00689176f $X=4.62 $Y=1.95 $X2=0 $Y2=0
cc_375 N_A_116_392#_c_538_p N_X_c_704_n 0.0277622f $X=5.52 $Y=1.465 $X2=0 $Y2=0
cc_376 N_A_116_392#_c_409_n N_X_c_704_n 0.00814019f $X=6.14 $Y=1.532 $X2=0 $Y2=0
cc_377 N_A_116_392#_M1013_g N_X_c_696_n 8.71574e-19 $X=5.21 $Y=0.74 $X2=0 $Y2=0
cc_378 N_A_116_392#_M1021_g N_X_c_696_n 0.0089455f $X=5.71 $Y=0.74 $X2=0 $Y2=0
cc_379 N_A_116_392#_M1022_g N_X_c_696_n 0.0167949f $X=6.14 $Y=0.74 $X2=0 $Y2=0
cc_380 N_A_116_392#_c_412_n N_X_c_705_n 8.7136e-19 $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_381 N_A_116_392#_c_413_n N_X_c_705_n 0.00168349f $X=6.165 $Y=1.765 $X2=0
+ $Y2=0
cc_382 N_A_116_392#_c_409_n N_X_c_705_n 0.00921806f $X=6.14 $Y=1.532 $X2=0 $Y2=0
cc_383 N_A_116_392#_c_412_n N_X_c_706_n 0.00476552f $X=5.715 $Y=1.765 $X2=0
+ $Y2=0
cc_384 N_A_116_392#_c_413_n N_X_c_706_n 0.0108676f $X=6.165 $Y=1.765 $X2=0 $Y2=0
cc_385 N_A_116_392#_M1022_g N_X_c_697_n 0.0133814f $X=6.14 $Y=0.74 $X2=0 $Y2=0
cc_386 N_A_116_392#_c_409_n N_X_c_697_n 0.00109998f $X=6.14 $Y=1.532 $X2=0 $Y2=0
cc_387 N_A_116_392#_c_409_n N_X_c_698_n 0.0149907f $X=6.14 $Y=1.532 $X2=0 $Y2=0
cc_388 N_A_116_392#_c_538_p N_X_c_699_n 0.012613f $X=5.52 $Y=1.465 $X2=0 $Y2=0
cc_389 N_A_116_392#_c_409_n N_X_c_699_n 0.0163181f $X=6.14 $Y=1.532 $X2=0 $Y2=0
cc_390 N_A_116_392#_M1021_g N_X_c_700_n 0.00132316f $X=5.71 $Y=0.74 $X2=0 $Y2=0
cc_391 N_A_116_392#_M1022_g N_X_c_700_n 0.00108831f $X=6.14 $Y=0.74 $X2=0 $Y2=0
cc_392 N_A_116_392#_c_409_n N_X_c_700_n 0.0026075f $X=6.14 $Y=1.532 $X2=0 $Y2=0
cc_393 N_A_116_392#_c_413_n N_X_c_743_n 0.00292387f $X=6.165 $Y=1.765 $X2=0
+ $Y2=0
cc_394 N_A_116_392#_M1022_g X 0.00612865f $X=6.14 $Y=0.74 $X2=0 $Y2=0
cc_395 N_A_116_392#_c_409_n X 0.00819458f $X=6.14 $Y=1.532 $X2=0 $Y2=0
cc_396 N_A_116_392#_c_431_n N_A_32_119#_c_771_n 0.00727685f $X=0.89 $Y=1.13
+ $X2=0 $Y2=0
cc_397 N_A_116_392#_c_406_n N_A_32_119#_c_775_n 0.0330606f $X=2.43 $Y=1.685
+ $X2=0 $Y2=0
cc_398 N_A_116_392#_c_465_n N_A_32_119#_c_775_n 0.0167929f $X=3.815 $Y=2.055
+ $X2=0 $Y2=0
cc_399 N_A_116_392#_c_405_n N_A_32_119#_c_776_n 0.00211728f $X=1.165 $Y=1.09
+ $X2=0 $Y2=0
cc_400 N_A_116_392#_c_406_n N_A_32_119#_c_776_n 0.00966614f $X=2.43 $Y=1.685
+ $X2=0 $Y2=0
cc_401 N_A_116_392#_c_431_n N_A_119_119#_M1002_d 0.00366647f $X=0.89 $Y=1.13
+ $X2=-0.19 $Y2=-0.245
cc_402 N_A_116_392#_M1001_d N_A_119_119#_c_820_n 0.00315171f $X=1.025 $Y=0.595
+ $X2=0 $Y2=0
cc_403 N_A_116_392#_c_431_n N_A_119_119#_c_820_n 0.00911672f $X=0.89 $Y=1.13
+ $X2=0 $Y2=0
cc_404 N_A_116_392#_c_405_n N_A_119_119#_c_820_n 0.0235835f $X=1.165 $Y=1.09
+ $X2=0 $Y2=0
cc_405 N_A_116_392#_M1007_g N_VGND_c_860_n 0.00254859f $X=4.75 $Y=0.74 $X2=0
+ $Y2=0
cc_406 N_A_116_392#_c_408_n N_VGND_c_860_n 0.0116185f $X=4.705 $Y=1.465 $X2=0
+ $Y2=0
cc_407 N_A_116_392#_M1007_g N_VGND_c_861_n 4.58515e-19 $X=4.75 $Y=0.74 $X2=0
+ $Y2=0
cc_408 N_A_116_392#_M1013_g N_VGND_c_861_n 0.00973022f $X=5.21 $Y=0.74 $X2=0
+ $Y2=0
cc_409 N_A_116_392#_M1021_g N_VGND_c_861_n 0.00406778f $X=5.71 $Y=0.74 $X2=0
+ $Y2=0
cc_410 N_A_116_392#_M1022_g N_VGND_c_863_n 0.00364571f $X=6.14 $Y=0.74 $X2=0
+ $Y2=0
cc_411 N_A_116_392#_M1007_g N_VGND_c_864_n 0.00461464f $X=4.75 $Y=0.74 $X2=0
+ $Y2=0
cc_412 N_A_116_392#_M1013_g N_VGND_c_864_n 0.00383152f $X=5.21 $Y=0.74 $X2=0
+ $Y2=0
cc_413 N_A_116_392#_M1021_g N_VGND_c_868_n 0.00434272f $X=5.71 $Y=0.74 $X2=0
+ $Y2=0
cc_414 N_A_116_392#_M1022_g N_VGND_c_868_n 0.00434272f $X=6.14 $Y=0.74 $X2=0
+ $Y2=0
cc_415 N_A_116_392#_M1007_g N_VGND_c_871_n 0.00908834f $X=4.75 $Y=0.74 $X2=0
+ $Y2=0
cc_416 N_A_116_392#_M1013_g N_VGND_c_871_n 0.00757833f $X=5.21 $Y=0.74 $X2=0
+ $Y2=0
cc_417 N_A_116_392#_M1021_g N_VGND_c_871_n 0.00820718f $X=5.71 $Y=0.74 $X2=0
+ $Y2=0
cc_418 N_A_116_392#_M1022_g N_VGND_c_871_n 0.00823975f $X=6.14 $Y=0.74 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_599_n N_X_c_702_n 0.00127913f $X=4.48 $Y=2.455 $X2=0 $Y2=0
cc_420 N_VPWR_c_600_n N_X_c_702_n 0.0563525f $X=5.49 $Y=2.305 $X2=0 $Y2=0
cc_421 N_VPWR_c_607_n N_X_c_702_n 0.0145938f $X=5.405 $Y=3.33 $X2=0 $Y2=0
cc_422 N_VPWR_c_593_n N_X_c_702_n 0.0120466f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_423 N_VPWR_M1008_s N_X_c_703_n 0.00222494f $X=5.34 $Y=1.84 $X2=0 $Y2=0
cc_424 N_VPWR_c_600_n N_X_c_703_n 0.0154248f $X=5.49 $Y=2.305 $X2=0 $Y2=0
cc_425 N_VPWR_c_600_n N_X_c_706_n 0.0551997f $X=5.49 $Y=2.305 $X2=0 $Y2=0
cc_426 N_VPWR_c_602_n N_X_c_706_n 0.0370736f $X=6.44 $Y=1.985 $X2=0 $Y2=0
cc_427 N_VPWR_c_608_n N_X_c_706_n 0.0110241f $X=6.275 $Y=3.33 $X2=0 $Y2=0
cc_428 N_VPWR_c_593_n N_X_c_706_n 0.00909194f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_429 N_VPWR_c_602_n N_X_c_698_n 0.0290533f $X=6.44 $Y=1.985 $X2=0 $Y2=0
cc_430 N_VPWR_c_602_n N_X_c_743_n 0.00711242f $X=6.44 $Y=1.985 $X2=0 $Y2=0
cc_431 N_X_c_694_n N_VGND_M1013_d 0.00250873f $X=5.76 $Y=1.045 $X2=0 $Y2=0
cc_432 N_X_c_697_n N_VGND_M1022_d 0.00409179f $X=6.365 $Y=1.045 $X2=0 $Y2=0
cc_433 N_X_c_693_n N_VGND_c_860_n 0.00154841f $X=4.995 $Y=0.515 $X2=0 $Y2=0
cc_434 N_X_c_695_n N_VGND_c_860_n 0.00167954f $X=5.08 $Y=1.045 $X2=0 $Y2=0
cc_435 N_X_c_693_n N_VGND_c_861_n 0.0164981f $X=4.995 $Y=0.515 $X2=0 $Y2=0
cc_436 N_X_c_694_n N_VGND_c_861_n 0.0209867f $X=5.76 $Y=1.045 $X2=0 $Y2=0
cc_437 N_X_c_696_n N_VGND_c_861_n 0.0173003f $X=5.925 $Y=0.515 $X2=0 $Y2=0
cc_438 N_X_c_696_n N_VGND_c_863_n 0.0131449f $X=5.925 $Y=0.515 $X2=0 $Y2=0
cc_439 N_X_c_697_n N_VGND_c_863_n 0.0148546f $X=6.365 $Y=1.045 $X2=0 $Y2=0
cc_440 N_X_c_693_n N_VGND_c_864_n 0.011066f $X=4.995 $Y=0.515 $X2=0 $Y2=0
cc_441 N_X_c_696_n N_VGND_c_868_n 0.0144922f $X=5.925 $Y=0.515 $X2=0 $Y2=0
cc_442 N_X_c_693_n N_VGND_c_871_n 0.00915947f $X=4.995 $Y=0.515 $X2=0 $Y2=0
cc_443 N_X_c_696_n N_VGND_c_871_n 0.0118826f $X=5.925 $Y=0.515 $X2=0 $Y2=0
cc_444 N_A_32_119#_c_772_n N_A_119_119#_c_820_n 0.0706419f $X=1.94 $Y=0.4 $X2=0
+ $Y2=0
cc_445 N_A_32_119#_c_775_n N_A_463_119#_M1019_d 0.00176461f $X=3.64 $Y=1.215
+ $X2=-0.19 $Y2=-0.245
cc_446 N_A_32_119#_c_775_n N_A_463_119#_M1018_s 0.00205484f $X=3.64 $Y=1.215
+ $X2=0 $Y2=0
cc_447 N_A_32_119#_c_775_n N_A_463_119#_c_832_n 0.0399118f $X=3.64 $Y=1.215
+ $X2=0 $Y2=0
cc_448 N_A_32_119#_c_774_n N_A_463_119#_c_830_n 0.0144855f $X=2.025 $Y=0.74
+ $X2=0 $Y2=0
cc_449 N_A_32_119#_c_775_n N_A_463_119#_c_830_n 0.0163142f $X=3.64 $Y=1.215
+ $X2=0 $Y2=0
cc_450 N_A_32_119#_c_775_n N_A_463_119#_c_831_n 0.0139562f $X=3.64 $Y=1.215
+ $X2=0 $Y2=0
cc_451 N_A_32_119#_c_775_n N_VGND_M1012_d 0.00393441f $X=3.64 $Y=1.215 $X2=-0.19
+ $Y2=-0.245
cc_452 N_A_32_119#_c_775_n N_VGND_c_860_n 0.00854438f $X=3.64 $Y=1.215 $X2=0
+ $Y2=0
cc_453 N_A_32_119#_c_772_n N_VGND_c_866_n 0.0805444f $X=1.94 $Y=0.4 $X2=0 $Y2=0
cc_454 N_A_32_119#_c_773_n N_VGND_c_866_n 0.0129707f $X=0.39 $Y=0.4 $X2=0 $Y2=0
cc_455 N_A_32_119#_c_772_n N_VGND_c_871_n 0.0564887f $X=1.94 $Y=0.4 $X2=0 $Y2=0
cc_456 N_A_32_119#_c_773_n N_VGND_c_871_n 0.00942301f $X=0.39 $Y=0.4 $X2=0 $Y2=0
cc_457 N_A_463_119#_c_832_n N_VGND_M1012_d 0.00687044f $X=3.3 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_458 N_A_463_119#_c_832_n N_VGND_c_859_n 0.0258995f $X=3.3 $Y=0.875 $X2=0
+ $Y2=0
cc_459 N_A_463_119#_c_830_n N_VGND_c_859_n 0.00237208f $X=2.455 $Y=0.765 $X2=0
+ $Y2=0
cc_460 N_A_463_119#_c_831_n N_VGND_c_859_n 0.00249965f $X=3.475 $Y=0.74 $X2=0
+ $Y2=0
cc_461 N_A_463_119#_c_830_n N_VGND_c_866_n 0.00714062f $X=2.455 $Y=0.765 $X2=0
+ $Y2=0
cc_462 N_A_463_119#_c_831_n N_VGND_c_867_n 0.00726962f $X=3.475 $Y=0.74 $X2=0
+ $Y2=0
cc_463 N_A_463_119#_c_832_n N_VGND_c_871_n 0.0116638f $X=3.3 $Y=0.875 $X2=0
+ $Y2=0
cc_464 N_A_463_119#_c_830_n N_VGND_c_871_n 0.00877363f $X=2.455 $Y=0.765 $X2=0
+ $Y2=0
cc_465 N_A_463_119#_c_831_n N_VGND_c_871_n 0.00899467f $X=3.475 $Y=0.74 $X2=0
+ $Y2=0
