* File: sky130_fd_sc_ls__o21ai_4.spice
* Created: Wed Sep  2 11:18:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o21ai_4.pex.spice"
.subckt sky130_fd_sc_ls__o21ai_4  VNB VPB A1 B1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* B1	B1
* A1	A1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A1_M1008_g N_A_27_74#_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75005 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1008_d N_A1_M1016_g N_A_27_74#_M1016_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75004.5 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A1_M1017_g N_A_27_74#_M1016_s VNB NSHORT L=0.15 W=0.74
+ AD=0.10915 AS=0.1036 PD=1.035 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75004.1 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1017_d N_A1_M1019_g N_A_27_74#_M1019_s VNB NSHORT L=0.15 W=0.74
+ AD=0.10915 AS=0.1036 PD=1.035 PS=1.02 NRD=2.424 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75003.7 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g N_A_27_74#_M1019_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1003_d N_B1_M1004_g N_A_27_74#_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1009_d N_B1_M1009_g N_A_27_74#_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1018 N_Y_M1009_d N_B1_M1018_g N_A_27_74#_M1018_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.11285 PD=1.02 PS=1.045 NRD=0 NRS=4.044 M=1 R=4.93333 SA=75003.2
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_27_74#_M1018_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.11285 PD=1.02 PS=1.045 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.7
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1000_d N_A2_M1007_g N_A_27_74#_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.1
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_A2_M1014_g N_A_27_74#_M1007_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.5
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1014_d N_A2_M1021_g N_A_27_74#_M1021_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75005
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g N_A_116_368#_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1012 N_VPWR_M1012_d N_A1_M1012_g N_A_116_368#_M1001_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1012_d N_A1_M1013_g N_A_116_368#_M1013_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1015 N_VPWR_M1015_d N_A1_M1015_g N_A_116_368#_M1013_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1005 N_Y_M1005_d N_B1_M1005_g N_VPWR_M1015_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75000.8 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1005_d N_B1_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.4256 PD=1.42 PS=3 NRD=1.7533 NRS=16.7056 M=1 R=7.46667
+ SA=75002.5 SB=75000.3 A=0.168 P=2.54 MULT=1
MM1002 N_A_116_368#_M1002_d N_A2_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1006 N_A_116_368#_M1006_d N_A2_M1006_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1010 N_A_116_368#_M1006_d N_A2_M1010_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1020 N_A_116_368#_M1020_d N_A2_M1020_g N_Y_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX22_noxref VNB VPB NWDIODE A=11.4204 P=16
c_51 VNB 0 1.07857e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ls__o21ai_4.pxi.spice"
*
.ends
*
*
