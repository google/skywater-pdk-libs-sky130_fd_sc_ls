* NGSPICE file created from sky130_fd_sc_ls__a41o_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 VPWR a_113_98# X VPB phighvt w=1.12e+06u l=150000u
+  ad=2.6382e+12p pd=1.979e+07u as=6.72e+11p ps=5.68e+06u
M1001 VGND a_113_98# X VNB nshort w=740000u l=150000u
+  ad=1.5409e+12p pd=1.26e+07u as=4.144e+11p ps=4.08e+06u
M1002 a_1205_74# A4 VGND VNB nshort w=740000u l=150000u
+  ad=6.216e+11p pd=6.12e+06u as=0p ps=0u
M1003 a_1205_74# A3 a_1010_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1004 VPWR A3 a_27_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.035e+12p ps=1.607e+07u
M1005 X a_113_98# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_113_98# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_751_74# A2 a_1010_74# VNB nshort w=740000u l=150000u
+  ad=6.216e+11p pd=6.12e+06u as=0p ps=0u
M1008 a_113_98# B1 VGND VNB nshort w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1009 a_27_392# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_392# A4 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_113_98# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_113_98# A1 a_751_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_751_74# A1 a_113_98# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A4 a_1205_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_113_98# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_392# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND B1 a_113_98# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1010_74# A3 a_1205_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A1 a_27_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A4 a_27_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_113_98# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_392# B1 a_113_98# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=3.5e+11p ps=2.7e+06u
M1023 a_113_98# B1 a_27_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A2 a_27_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 X a_113_98# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1010_74# A2 a_751_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_27_392# A3 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

