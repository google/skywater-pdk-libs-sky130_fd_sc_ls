* File: sky130_fd_sc_ls__decaphe_6.pxi.spice
* Created: Fri Aug 28 13:12:42 2020
* 
x_PM_SKY130_FD_SC_LS__DECAPHE_6%VGND N_VGND_M1000_s N_VGND_c_13_n N_VGND_c_14_n
+ VGND N_VGND_c_15_n N_VGND_M1001_g N_VGND_c_16_n N_VGND_c_17_n
+ PM_SKY130_FD_SC_LS__DECAPHE_6%VGND
x_PM_SKY130_FD_SC_LS__DECAPHE_6%VPWR N_VPWR_M1001_s N_VPWR_M1000_g VPWR
+ N_VPWR_c_31_n N_VPWR_c_32_n N_VPWR_c_33_n VPWR
+ PM_SKY130_FD_SC_LS__DECAPHE_6%VPWR
cc_1 VNB N_VGND_c_13_n 0.0130276f $X=-0.19 $Y=-0.245 $X2=2.178 $Y2=0.497
cc_2 VNB N_VGND_c_14_n 0.0883521f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=0.497
cc_3 VNB N_VGND_c_15_n 0.0470015f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.515
cc_4 VNB N_VGND_c_16_n 0.0542007f $X=-0.19 $Y=-0.245 $X2=2.62 $Y2=0.38
cc_5 VNB N_VGND_c_17_n 0.169234f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0
cc_6 VNB VPWR 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_VPWR_c_31_n 0.0839869f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=2.467
cc_8 VNB N_VPWR_c_32_n 0.137489f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0
cc_9 VNB N_VPWR_c_33_n 0.0245969f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0
cc_10 VPB N_VGND_c_15_n 0.161761f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=1.515
cc_11 VPB VPWR 0.0453372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_12 VPB N_VPWR_c_33_n 0.1706f $X=-0.19 $Y=1.66 $X2=2.64 $Y2=0
cc_13 N_VGND_c_13_n N_VPWR_c_31_n 0.0330165f $X=2.178 $Y=0.497 $X2=0 $Y2=0
cc_14 N_VGND_c_14_n N_VPWR_c_31_n 0.110835f $X=1.195 $Y=0.497 $X2=0 $Y2=0
cc_15 N_VGND_c_15_n N_VPWR_c_31_n 0.0515862f $X=0.915 $Y=1.515 $X2=0 $Y2=0
cc_16 N_VGND_c_13_n N_VPWR_c_32_n 0.0888789f $X=2.178 $Y=0.497 $X2=0 $Y2=0
cc_17 N_VGND_c_14_n N_VPWR_c_32_n 0.00593011f $X=1.195 $Y=0.497 $X2=0 $Y2=0
cc_18 N_VGND_c_15_n N_VPWR_c_32_n 0.0715919f $X=0.915 $Y=1.515 $X2=0 $Y2=0
cc_19 N_VGND_c_16_n N_VPWR_c_32_n 0.0437934f $X=2.62 $Y=0.38 $X2=0 $Y2=0
cc_20 N_VGND_c_13_n N_VPWR_c_33_n 0.0688373f $X=2.178 $Y=0.497 $X2=0 $Y2=0
cc_21 N_VGND_c_14_n N_VPWR_c_33_n 0.126794f $X=1.195 $Y=0.497 $X2=0 $Y2=0
cc_22 N_VGND_c_15_n N_VPWR_c_33_n 0.380599f $X=0.915 $Y=1.515 $X2=0 $Y2=0
cc_23 N_VGND_c_16_n N_VPWR_c_33_n 0.0517547f $X=2.62 $Y=0.38 $X2=0 $Y2=0
