* File: sky130_fd_sc_ls__or2_4.spice
* Created: Fri Aug 28 13:57:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__or2_4.pex.spice"
.subckt sky130_fd_sc_ls__or2_4  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_X_M1005_d N_A_83_260#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1006 N_X_M1005_d N_A_83_260#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1012 N_X_M1012_d N_A_83_260#_M1012_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.74
+ AD=0.13505 AS=0.1036 PD=1.105 PS=1.02 NRD=3.24 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1012_d N_A_83_260#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.13505 AS=0.1295 PD=1.105 PS=1.09 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_83_260#_M1004_d N_A_M1004_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.12395 AS=0.1295 PD=1.075 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.1
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_B_M1002_g N_A_83_260#_M1004_d VNB NSHORT L=0.15 W=0.74
+ AD=0.9287 AS=0.12395 PD=3.99 PS=1.075 NRD=0 NRS=8.916 M=1 R=4.93333 SA=75002.6
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_A_83_260#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.3 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1008_d N_A_83_260#_M1008_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75002.9 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1008_d N_A_83_260#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_83_260#_M1011_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.222098 AS=0.168 PD=1.59019 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75002 A=0.168 P=2.54 MULT=1
MM1000 N_A_493_388#_M1000_d N_A_M1000_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.198302 PD=1.3 PS=1.41981 NRD=1.9503 NRS=18.715 M=1 R=6.66667
+ SA=75002.1 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1003 N_A_83_260#_M1003_d N_B_M1003_g N_A_493_388#_M1000_d VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75002.6 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1007 N_A_83_260#_M1003_d N_B_M1007_g N_A_493_388#_M1007_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75003 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1010 N_A_493_388#_M1007_s N_A_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.32 PD=1.35 PS=2.64 NRD=1.9503 NRS=3.9203 M=1 R=6.66667
+ SA=75003.5 SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ls__or2_4.pxi.spice"
*
.ends
*
*
