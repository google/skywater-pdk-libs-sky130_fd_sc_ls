* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 VPWR B1 a_1215_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VPWR A2_N a_114_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 VPWR B1 a_1215_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 Y a_114_368# a_857_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 VPWR A1_N a_114_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X5 a_857_74# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 Y B2 a_1215_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 VGND A1_N a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X8 a_27_74# A2_N a_114_368# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 a_114_368# A2_N a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X10 VPWR a_114_368# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X11 Y B2 a_1215_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X12 VPWR A1_N a_114_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X13 a_114_368# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 Y a_114_368# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X15 a_857_74# a_114_368# Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 a_114_368# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X17 a_1215_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X18 a_114_368# A2_N a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X19 VGND B2 a_857_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X20 a_857_74# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 VGND B1 a_857_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 a_114_368# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X23 a_1215_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X24 a_114_368# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X25 a_1215_368# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X26 a_1215_368# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X27 a_27_74# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X28 Y a_114_368# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X29 a_857_74# a_114_368# Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X30 VGND B2 a_857_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X31 a_27_74# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X32 a_857_74# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X33 VGND B1 a_857_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X34 VPWR a_114_368# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X35 VGND A1_N a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X36 Y a_114_368# a_857_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X37 a_857_74# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X38 a_27_74# A2_N a_114_368# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X39 VPWR A2_N a_114_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
.ends
