* File: sky130_fd_sc_ls__a21bo_2.pxi.spice
* Created: Fri Aug 28 12:50:17 2020
* 
x_PM_SKY130_FD_SC_LS__A21BO_2%B1_N N_B1_N_c_72_n N_B1_N_M1005_g N_B1_N_c_73_n
+ N_B1_N_M1009_g B1_N N_B1_N_c_74_n PM_SKY130_FD_SC_LS__A21BO_2%B1_N
x_PM_SKY130_FD_SC_LS__A21BO_2%A_187_244# N_A_187_244#_M1002_d
+ N_A_187_244#_M1007_s N_A_187_244#_c_99_n N_A_187_244#_c_107_n
+ N_A_187_244#_M1001_g N_A_187_244#_c_100_n N_A_187_244#_M1004_g
+ N_A_187_244#_c_108_n N_A_187_244#_M1003_g N_A_187_244#_c_101_n
+ N_A_187_244#_M1011_g N_A_187_244#_c_117_p N_A_187_244#_c_102_n
+ N_A_187_244#_c_103_n N_A_187_244#_c_104_n N_A_187_244#_c_105_n
+ N_A_187_244#_c_111_n N_A_187_244#_c_121_p
+ PM_SKY130_FD_SC_LS__A21BO_2%A_187_244#
x_PM_SKY130_FD_SC_LS__A21BO_2%A_32_368# N_A_32_368#_M1009_s N_A_32_368#_M1005_s
+ N_A_32_368#_M1002_g N_A_32_368#_c_206_n N_A_32_368#_M1007_g
+ N_A_32_368#_c_200_n N_A_32_368#_c_201_n N_A_32_368#_c_202_n
+ N_A_32_368#_c_208_n N_A_32_368#_c_214_n N_A_32_368#_c_209_n
+ N_A_32_368#_c_203_n N_A_32_368#_c_240_n N_A_32_368#_c_204_n
+ N_A_32_368#_c_249_n N_A_32_368#_c_205_n N_A_32_368#_c_261_p
+ PM_SKY130_FD_SC_LS__A21BO_2%A_32_368#
x_PM_SKY130_FD_SC_LS__A21BO_2%A1 N_A1_M1010_g N_A1_c_294_n N_A1_c_298_n
+ N_A1_M1008_g A1 N_A1_c_295_n N_A1_c_296_n PM_SKY130_FD_SC_LS__A21BO_2%A1
x_PM_SKY130_FD_SC_LS__A21BO_2%A2 N_A2_M1006_g N_A2_c_339_n N_A2_M1000_g A2
+ PM_SKY130_FD_SC_LS__A21BO_2%A2
x_PM_SKY130_FD_SC_LS__A21BO_2%VPWR N_VPWR_M1005_d N_VPWR_M1003_s N_VPWR_M1008_d
+ N_VPWR_c_364_n N_VPWR_c_365_n N_VPWR_c_366_n VPWR N_VPWR_c_367_n
+ N_VPWR_c_368_n N_VPWR_c_369_n N_VPWR_c_370_n N_VPWR_c_363_n N_VPWR_c_372_n
+ N_VPWR_c_373_n N_VPWR_c_374_n PM_SKY130_FD_SC_LS__A21BO_2%VPWR
x_PM_SKY130_FD_SC_LS__A21BO_2%X N_X_M1004_d N_X_M1001_d N_X_c_421_n N_X_c_422_n
+ N_X_c_424_n X PM_SKY130_FD_SC_LS__A21BO_2%X
x_PM_SKY130_FD_SC_LS__A21BO_2%A_504_392# N_A_504_392#_M1007_d
+ N_A_504_392#_M1000_d N_A_504_392#_c_462_n N_A_504_392#_c_457_n
+ N_A_504_392#_c_458_n N_A_504_392#_c_459_n
+ PM_SKY130_FD_SC_LS__A21BO_2%A_504_392#
x_PM_SKY130_FD_SC_LS__A21BO_2%VGND N_VGND_M1009_d N_VGND_M1011_s N_VGND_M1006_d
+ N_VGND_c_482_n N_VGND_c_483_n N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n
+ N_VGND_c_487_n VGND N_VGND_c_488_n N_VGND_c_489_n N_VGND_c_490_n
+ N_VGND_c_491_n PM_SKY130_FD_SC_LS__A21BO_2%VGND
cc_1 VNB N_B1_N_c_72_n 0.0631144f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.765
cc_2 VNB N_B1_N_c_73_n 0.0228559f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.22
cc_3 VNB N_B1_N_c_74_n 0.0225328f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.385
cc_4 VNB N_A_187_244#_c_99_n 0.0142239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_A_187_244#_c_100_n 0.0176121f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_6 VNB N_A_187_244#_c_101_n 0.019167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_187_244#_c_102_n 0.00881618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_187_244#_c_103_n 0.00390742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_187_244#_c_104_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_187_244#_c_105_n 0.0535198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_32_368#_M1002_g 0.0221011f $X=-0.19 $Y=-0.245 $X2=0.452 $Y2=1.385
cc_12 VNB N_A_32_368#_c_200_n 0.0465265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_32_368#_c_201_n 0.00860503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_32_368#_c_202_n 0.00372942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_32_368#_c_203_n 0.00426191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_32_368#_c_204_n 0.00620465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_32_368#_c_205_n 0.0225067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_M1010_g 0.0204236f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.26
cc_19 VNB N_A1_c_294_n 0.00318739f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.835
cc_20 VNB N_A1_c_295_n 0.0297901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_296_n 0.0159715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_M1006_g 0.0408671f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.26
cc_23 VNB N_A2_c_339_n 0.0348821f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.835
cc_24 VNB A2 0.00472574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_363_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_421_n 0.00239017f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_27 VNB N_X_c_422_n 0.00285947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_482_n 0.0157102f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_29 VNB N_VGND_c_483_n 0.0124379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_484_n 0.0125057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_485_n 0.037498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_486_n 0.0259864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_487_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_488_n 0.0189193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_489_n 0.0312656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_490_n 0.01106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_491_n 0.243653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_B1_N_c_72_n 0.0312809f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_39 VPB N_A_187_244#_c_99_n 7.39253e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_187_244#_c_107_n 0.0225482f $X=-0.19 $Y=1.66 $X2=0.452 $Y2=1.385
cc_41 VPB N_A_187_244#_c_108_n 0.0170807f $X=-0.19 $Y=1.66 $X2=0.345 $Y2=1.365
cc_42 VPB N_A_187_244#_c_103_n 6.19153e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_187_244#_c_105_n 0.00713204f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_187_244#_c_111_n 0.0186717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_32_368#_c_206_n 0.0287527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_32_368#_c_202_n 0.00372942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_32_368#_c_208_n 0.0188199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_32_368#_c_209_n 0.022634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_32_368#_c_203_n 0.00325623f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_32_368#_c_204_n 0.017765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A1_c_294_n 0.00627606f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=0.835
cc_52 VPB N_A1_c_298_n 0.0214598f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_53 VPB N_A1_c_296_n 0.00540584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A2_c_339_n 0.0543628f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=0.835
cc_55 VPB A2 0.00276779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_364_n 0.016612f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_57 VPB N_VPWR_c_365_n 0.0113776f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_366_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_367_n 0.0208665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_368_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_369_n 0.0303553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_370_n 0.0197879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_363_n 0.087454f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_372_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_373_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_374_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_X_c_422_n 0.00167527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_X_c_424_n 0.00267794f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_69 VPB N_A_504_392#_c_457_n 0.0148981f $X=-0.19 $Y=1.66 $X2=0.345 $Y2=1.385
cc_70 VPB N_A_504_392#_c_458_n 0.03021f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_504_392#_c_459_n 0.00179738f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 N_B1_N_c_72_n N_A_187_244#_c_99_n 0.00596292f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_73 N_B1_N_c_72_n N_A_187_244#_c_107_n 0.0248953f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_74 N_B1_N_c_73_n N_A_187_244#_c_100_n 0.0180021f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_75 N_B1_N_c_72_n N_A_187_244#_c_105_n 0.0205347f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_76 N_B1_N_c_72_n N_A_32_368#_c_208_n 0.0122036f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_77 N_B1_N_c_74_n N_A_32_368#_c_208_n 0.0196805f $X=0.345 $Y=1.385 $X2=0 $Y2=0
cc_78 N_B1_N_c_72_n N_A_32_368#_c_214_n 0.0174568f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_79 N_B1_N_c_72_n N_A_32_368#_c_209_n 0.00730766f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_80 N_B1_N_c_72_n N_A_32_368#_c_203_n 0.0185309f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_81 N_B1_N_c_73_n N_A_32_368#_c_203_n 0.00946285f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_82 N_B1_N_c_74_n N_A_32_368#_c_203_n 0.0268756f $X=0.345 $Y=1.385 $X2=0 $Y2=0
cc_83 N_B1_N_c_72_n N_A_32_368#_c_205_n 0.00331257f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_84 N_B1_N_c_73_n N_A_32_368#_c_205_n 0.018243f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_85 N_B1_N_c_74_n N_A_32_368#_c_205_n 0.0204716f $X=0.345 $Y=1.385 $X2=0 $Y2=0
cc_86 N_B1_N_c_72_n N_VPWR_c_364_n 0.00382931f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_87 N_B1_N_c_72_n N_VPWR_c_367_n 0.00393265f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_88 N_B1_N_c_72_n N_VPWR_c_363_n 0.00462577f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_89 N_B1_N_c_73_n N_X_c_421_n 0.00117035f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_90 N_B1_N_c_72_n N_X_c_422_n 2.83559e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_91 N_B1_N_c_73_n N_X_c_422_n 4.56618e-19 $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_92 N_B1_N_c_73_n N_VGND_c_482_n 0.00400491f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_93 N_B1_N_c_73_n N_VGND_c_486_n 0.00432822f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_94 N_B1_N_c_73_n N_VGND_c_491_n 0.00487769f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_95 N_A_187_244#_c_101_n N_A_32_368#_M1002_g 0.0084396f $X=1.615 $Y=1.22 $X2=0
+ $Y2=0
cc_96 N_A_187_244#_c_117_p N_A_32_368#_M1002_g 0.00596357f $X=2.385 $Y=1.005
+ $X2=0 $Y2=0
cc_97 N_A_187_244#_c_102_n N_A_32_368#_M1002_g 0.0010596f $X=1.735 $Y=1.005
+ $X2=0 $Y2=0
cc_98 N_A_187_244#_c_103_n N_A_32_368#_M1002_g 0.00527003f $X=2.47 $Y=1.76 $X2=0
+ $Y2=0
cc_99 N_A_187_244#_c_104_n N_A_32_368#_M1002_g 0.0122808f $X=2.645 $Y=0.515
+ $X2=0 $Y2=0
cc_100 N_A_187_244#_c_121_p N_A_32_368#_M1002_g 0.0068369f $X=2.597 $Y=1.005
+ $X2=0 $Y2=0
cc_101 N_A_187_244#_c_103_n N_A_32_368#_c_206_n 0.00151302f $X=2.47 $Y=1.76
+ $X2=0 $Y2=0
cc_102 N_A_187_244#_c_111_n N_A_32_368#_c_206_n 0.0329581f $X=2.22 $Y=2.225
+ $X2=0 $Y2=0
cc_103 N_A_187_244#_c_117_p N_A_32_368#_c_200_n 0.00602892f $X=2.385 $Y=1.005
+ $X2=0 $Y2=0
cc_104 N_A_187_244#_c_102_n N_A_32_368#_c_200_n 0.00180262f $X=1.735 $Y=1.005
+ $X2=0 $Y2=0
cc_105 N_A_187_244#_c_105_n N_A_32_368#_c_200_n 0.0206727f $X=1.525 $Y=1.385
+ $X2=0 $Y2=0
cc_106 N_A_187_244#_c_111_n N_A_32_368#_c_200_n 0.00530616f $X=2.22 $Y=2.225
+ $X2=0 $Y2=0
cc_107 N_A_187_244#_c_103_n N_A_32_368#_c_201_n 0.00903297f $X=2.47 $Y=1.76
+ $X2=0 $Y2=0
cc_108 N_A_187_244#_c_103_n N_A_32_368#_c_202_n 0.00353279f $X=2.47 $Y=1.76
+ $X2=0 $Y2=0
cc_109 N_A_187_244#_c_107_n N_A_32_368#_c_209_n 7.15205e-19 $X=1.025 $Y=1.765
+ $X2=0 $Y2=0
cc_110 N_A_187_244#_c_107_n N_A_32_368#_c_203_n 0.00625411f $X=1.025 $Y=1.765
+ $X2=0 $Y2=0
cc_111 N_A_187_244#_c_100_n N_A_32_368#_c_203_n 5.80921e-19 $X=1.185 $Y=1.22
+ $X2=0 $Y2=0
cc_112 N_A_187_244#_c_105_n N_A_32_368#_c_203_n 0.00367991f $X=1.525 $Y=1.385
+ $X2=0 $Y2=0
cc_113 N_A_187_244#_c_107_n N_A_32_368#_c_240_n 0.0172439f $X=1.025 $Y=1.765
+ $X2=0 $Y2=0
cc_114 N_A_187_244#_c_108_n N_A_32_368#_c_240_n 0.0201541f $X=1.475 $Y=1.765
+ $X2=0 $Y2=0
cc_115 N_A_187_244#_c_111_n N_A_32_368#_c_240_n 0.011361f $X=2.22 $Y=2.225 $X2=0
+ $Y2=0
cc_116 N_A_187_244#_c_108_n N_A_32_368#_c_204_n 0.00289451f $X=1.475 $Y=1.765
+ $X2=0 $Y2=0
cc_117 N_A_187_244#_c_117_p N_A_32_368#_c_204_n 0.0286626f $X=2.385 $Y=1.005
+ $X2=0 $Y2=0
cc_118 N_A_187_244#_c_102_n N_A_32_368#_c_204_n 0.0350515f $X=1.735 $Y=1.005
+ $X2=0 $Y2=0
cc_119 N_A_187_244#_c_103_n N_A_32_368#_c_204_n 0.0314791f $X=2.47 $Y=1.76 $X2=0
+ $Y2=0
cc_120 N_A_187_244#_c_105_n N_A_32_368#_c_204_n 0.00630425f $X=1.525 $Y=1.385
+ $X2=0 $Y2=0
cc_121 N_A_187_244#_c_111_n N_A_32_368#_c_204_n 0.0183437f $X=2.22 $Y=2.225
+ $X2=0 $Y2=0
cc_122 N_A_187_244#_c_111_n N_A_32_368#_c_249_n 0.0174709f $X=2.22 $Y=2.225
+ $X2=0 $Y2=0
cc_123 N_A_187_244#_c_100_n N_A_32_368#_c_205_n 0.00105802f $X=1.185 $Y=1.22
+ $X2=0 $Y2=0
cc_124 N_A_187_244#_c_103_n N_A1_M1010_g 0.00286552f $X=2.47 $Y=1.76 $X2=0 $Y2=0
cc_125 N_A_187_244#_c_104_n N_A1_M1010_g 0.0111096f $X=2.645 $Y=0.515 $X2=0
+ $Y2=0
cc_126 N_A_187_244#_c_121_p N_A1_M1010_g 0.00346711f $X=2.597 $Y=1.005 $X2=0
+ $Y2=0
cc_127 N_A_187_244#_c_103_n N_A1_c_294_n 4.44452e-19 $X=2.47 $Y=1.76 $X2=0 $Y2=0
cc_128 N_A_187_244#_c_111_n N_A1_c_294_n 0.00228162f $X=2.22 $Y=2.225 $X2=0
+ $Y2=0
cc_129 N_A_187_244#_c_111_n N_A1_c_298_n 0.00173306f $X=2.22 $Y=2.225 $X2=0
+ $Y2=0
cc_130 N_A_187_244#_c_103_n N_A1_c_295_n 0.00177514f $X=2.47 $Y=1.76 $X2=0 $Y2=0
cc_131 N_A_187_244#_c_121_p N_A1_c_295_n 7.83088e-19 $X=2.597 $Y=1.005 $X2=0
+ $Y2=0
cc_132 N_A_187_244#_c_103_n N_A1_c_296_n 0.0395719f $X=2.47 $Y=1.76 $X2=0 $Y2=0
cc_133 N_A_187_244#_c_111_n N_A1_c_296_n 0.00172161f $X=2.22 $Y=2.225 $X2=0
+ $Y2=0
cc_134 N_A_187_244#_c_121_p N_A1_c_296_n 0.00451909f $X=2.597 $Y=1.005 $X2=0
+ $Y2=0
cc_135 N_A_187_244#_c_104_n N_A2_M1006_g 0.00172432f $X=2.645 $Y=0.515 $X2=0
+ $Y2=0
cc_136 N_A_187_244#_c_121_p N_A2_M1006_g 5.12803e-19 $X=2.597 $Y=1.005 $X2=0
+ $Y2=0
cc_137 N_A_187_244#_c_107_n N_VPWR_c_364_n 0.0124521f $X=1.025 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A_187_244#_c_108_n N_VPWR_c_364_n 0.0015077f $X=1.475 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A_187_244#_c_107_n N_VPWR_c_365_n 0.0015077f $X=1.025 $Y=1.765 $X2=0
+ $Y2=0
cc_140 N_A_187_244#_c_108_n N_VPWR_c_365_n 0.0124521f $X=1.475 $Y=1.765 $X2=0
+ $Y2=0
cc_141 N_A_187_244#_c_111_n N_VPWR_c_365_n 0.031005f $X=2.22 $Y=2.225 $X2=0
+ $Y2=0
cc_142 N_A_187_244#_c_107_n N_VPWR_c_368_n 0.00413917f $X=1.025 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_A_187_244#_c_108_n N_VPWR_c_368_n 0.00413917f $X=1.475 $Y=1.765 $X2=0
+ $Y2=0
cc_144 N_A_187_244#_c_111_n N_VPWR_c_369_n 0.0158428f $X=2.22 $Y=2.225 $X2=0
+ $Y2=0
cc_145 N_A_187_244#_c_107_n N_VPWR_c_363_n 0.00817726f $X=1.025 $Y=1.765 $X2=0
+ $Y2=0
cc_146 N_A_187_244#_c_108_n N_VPWR_c_363_n 0.00817726f $X=1.475 $Y=1.765 $X2=0
+ $Y2=0
cc_147 N_A_187_244#_c_111_n N_VPWR_c_363_n 0.0130099f $X=2.22 $Y=2.225 $X2=0
+ $Y2=0
cc_148 N_A_187_244#_c_100_n N_X_c_421_n 0.0201735f $X=1.185 $Y=1.22 $X2=0 $Y2=0
cc_149 N_A_187_244#_c_101_n N_X_c_421_n 0.0101064f $X=1.615 $Y=1.22 $X2=0 $Y2=0
cc_150 N_A_187_244#_c_102_n N_X_c_421_n 0.0177631f $X=1.735 $Y=1.005 $X2=0 $Y2=0
cc_151 N_A_187_244#_c_105_n N_X_c_421_n 0.00101877f $X=1.525 $Y=1.385 $X2=0
+ $Y2=0
cc_152 N_A_187_244#_c_99_n N_X_c_422_n 0.00618282f $X=1.025 $Y=1.675 $X2=0 $Y2=0
cc_153 N_A_187_244#_c_107_n N_X_c_422_n 0.00345187f $X=1.025 $Y=1.765 $X2=0
+ $Y2=0
cc_154 N_A_187_244#_c_100_n N_X_c_422_n 0.00468919f $X=1.185 $Y=1.22 $X2=0 $Y2=0
cc_155 N_A_187_244#_c_108_n N_X_c_422_n 4.24274e-19 $X=1.475 $Y=1.765 $X2=0
+ $Y2=0
cc_156 N_A_187_244#_c_101_n N_X_c_422_n 5.48773e-19 $X=1.615 $Y=1.22 $X2=0 $Y2=0
cc_157 N_A_187_244#_c_102_n N_X_c_422_n 0.0312442f $X=1.735 $Y=1.005 $X2=0 $Y2=0
cc_158 N_A_187_244#_c_105_n N_X_c_422_n 0.0132689f $X=1.525 $Y=1.385 $X2=0 $Y2=0
cc_159 N_A_187_244#_c_107_n N_X_c_424_n 0.00515697f $X=1.025 $Y=1.765 $X2=0
+ $Y2=0
cc_160 N_A_187_244#_c_108_n N_X_c_424_n 0.00330018f $X=1.475 $Y=1.765 $X2=0
+ $Y2=0
cc_161 N_A_187_244#_c_102_n N_X_c_424_n 0.00296465f $X=1.735 $Y=1.005 $X2=0
+ $Y2=0
cc_162 N_A_187_244#_c_105_n N_X_c_424_n 0.00623749f $X=1.525 $Y=1.385 $X2=0
+ $Y2=0
cc_163 N_A_187_244#_c_111_n N_A_504_392#_c_459_n 0.0669149f $X=2.22 $Y=2.225
+ $X2=0 $Y2=0
cc_164 N_A_187_244#_c_117_p N_VGND_M1011_s 0.0154162f $X=2.385 $Y=1.005 $X2=0
+ $Y2=0
cc_165 N_A_187_244#_c_100_n N_VGND_c_482_n 0.00487752f $X=1.185 $Y=1.22 $X2=0
+ $Y2=0
cc_166 N_A_187_244#_c_105_n N_VGND_c_482_n 0.0028854f $X=1.525 $Y=1.385 $X2=0
+ $Y2=0
cc_167 N_A_187_244#_c_101_n N_VGND_c_483_n 0.00422881f $X=1.615 $Y=1.22 $X2=0
+ $Y2=0
cc_168 N_A_187_244#_c_117_p N_VGND_c_483_n 0.0448286f $X=2.385 $Y=1.005 $X2=0
+ $Y2=0
cc_169 N_A_187_244#_c_104_n N_VGND_c_483_n 0.0158686f $X=2.645 $Y=0.515 $X2=0
+ $Y2=0
cc_170 N_A_187_244#_c_104_n N_VGND_c_485_n 0.0157759f $X=2.645 $Y=0.515 $X2=0
+ $Y2=0
cc_171 N_A_187_244#_c_121_p N_VGND_c_485_n 0.00499344f $X=2.597 $Y=1.005 $X2=0
+ $Y2=0
cc_172 N_A_187_244#_c_100_n N_VGND_c_488_n 0.00421809f $X=1.185 $Y=1.22 $X2=0
+ $Y2=0
cc_173 N_A_187_244#_c_101_n N_VGND_c_488_n 0.00433139f $X=1.615 $Y=1.22 $X2=0
+ $Y2=0
cc_174 N_A_187_244#_c_104_n N_VGND_c_489_n 0.0144922f $X=2.645 $Y=0.515 $X2=0
+ $Y2=0
cc_175 N_A_187_244#_c_100_n N_VGND_c_491_n 0.00443777f $X=1.185 $Y=1.22 $X2=0
+ $Y2=0
cc_176 N_A_187_244#_c_101_n N_VGND_c_491_n 0.00819075f $X=1.615 $Y=1.22 $X2=0
+ $Y2=0
cc_177 N_A_187_244#_c_104_n N_VGND_c_491_n 0.0118826f $X=2.645 $Y=0.515 $X2=0
+ $Y2=0
cc_178 N_A_32_368#_M1002_g N_A1_M1010_g 0.0130291f $X=2.43 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A_32_368#_c_206_n N_A1_c_294_n 0.00694015f $X=2.445 $Y=1.885 $X2=0
+ $Y2=0
cc_180 N_A_32_368#_c_202_n N_A1_c_294_n 0.00571367f $X=2.445 $Y=1.73 $X2=0 $Y2=0
cc_181 N_A_32_368#_c_206_n N_A1_c_298_n 0.0179938f $X=2.445 $Y=1.885 $X2=0 $Y2=0
cc_182 N_A_32_368#_c_201_n N_A1_c_295_n 0.0206661f $X=2.43 $Y=1.425 $X2=0 $Y2=0
cc_183 N_A_32_368#_c_201_n N_A1_c_296_n 3.61775e-19 $X=2.43 $Y=1.425 $X2=0 $Y2=0
cc_184 N_A_32_368#_c_202_n N_A1_c_296_n 4.76375e-19 $X=2.445 $Y=1.73 $X2=0 $Y2=0
cc_185 N_A_32_368#_c_214_n N_VPWR_M1005_d 0.00105873f $X=0.68 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_186 N_A_32_368#_c_203_n N_VPWR_M1005_d 0.00880663f $X=0.765 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_32_368#_c_240_n N_VPWR_M1005_d 0.002049f $X=1.605 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A_32_368#_c_261_p N_VPWR_M1005_d 0.00190618f $X=0.765 $Y=2.325
+ $X2=-0.19 $Y2=-0.245
cc_189 N_A_32_368#_c_240_n N_VPWR_M1003_s 0.00498928f $X=1.605 $Y=2.325 $X2=0
+ $Y2=0
cc_190 N_A_32_368#_c_204_n N_VPWR_M1003_s 0.00117646f $X=1.707 $Y=1.89 $X2=0
+ $Y2=0
cc_191 N_A_32_368#_c_249_n N_VPWR_M1003_s 0.00717805f $X=1.707 $Y=2.24 $X2=0
+ $Y2=0
cc_192 N_A_32_368#_c_214_n N_VPWR_c_364_n 0.00305515f $X=0.68 $Y=2.325 $X2=0
+ $Y2=0
cc_193 N_A_32_368#_c_209_n N_VPWR_c_364_n 0.0049774f $X=0.45 $Y=2.325 $X2=0
+ $Y2=0
cc_194 N_A_32_368#_c_240_n N_VPWR_c_364_n 0.00448627f $X=1.605 $Y=2.325 $X2=0
+ $Y2=0
cc_195 N_A_32_368#_c_261_p N_VPWR_c_364_n 0.0152373f $X=0.765 $Y=2.325 $X2=0
+ $Y2=0
cc_196 N_A_32_368#_c_206_n N_VPWR_c_365_n 0.00356994f $X=2.445 $Y=1.885 $X2=0
+ $Y2=0
cc_197 N_A_32_368#_c_240_n N_VPWR_c_365_n 0.019347f $X=1.605 $Y=2.325 $X2=0
+ $Y2=0
cc_198 N_A_32_368#_c_206_n N_VPWR_c_366_n 7.01755e-19 $X=2.445 $Y=1.885 $X2=0
+ $Y2=0
cc_199 N_A_32_368#_c_209_n N_VPWR_c_367_n 0.00671799f $X=0.45 $Y=2.325 $X2=0
+ $Y2=0
cc_200 N_A_32_368#_c_206_n N_VPWR_c_369_n 0.00411612f $X=2.445 $Y=1.885 $X2=0
+ $Y2=0
cc_201 N_A_32_368#_c_206_n N_VPWR_c_363_n 0.00753176f $X=2.445 $Y=1.885 $X2=0
+ $Y2=0
cc_202 N_A_32_368#_c_209_n N_VPWR_c_363_n 0.0100331f $X=0.45 $Y=2.325 $X2=0
+ $Y2=0
cc_203 N_A_32_368#_c_240_n N_X_M1001_d 0.00907897f $X=1.605 $Y=2.325 $X2=0 $Y2=0
cc_204 N_A_32_368#_c_203_n N_X_c_421_n 0.00229049f $X=0.765 $Y=2.24 $X2=0 $Y2=0
cc_205 N_A_32_368#_c_205_n N_X_c_421_n 0.0187392f $X=0.435 $Y=0.775 $X2=0 $Y2=0
cc_206 N_A_32_368#_c_203_n N_X_c_422_n 0.0561377f $X=0.765 $Y=2.24 $X2=0 $Y2=0
cc_207 N_A_32_368#_c_204_n N_X_c_422_n 0.00438932f $X=1.707 $Y=1.89 $X2=0 $Y2=0
cc_208 N_A_32_368#_c_203_n N_X_c_424_n 0.0186885f $X=0.765 $Y=2.24 $X2=0 $Y2=0
cc_209 N_A_32_368#_c_240_n N_X_c_424_n 0.0204393f $X=1.605 $Y=2.325 $X2=0 $Y2=0
cc_210 N_A_32_368#_c_204_n N_X_c_424_n 0.00319333f $X=1.707 $Y=1.89 $X2=0 $Y2=0
cc_211 N_A_32_368#_c_206_n N_A_504_392#_c_459_n 0.00271725f $X=2.445 $Y=1.885
+ $X2=0 $Y2=0
cc_212 N_A_32_368#_c_203_n N_VGND_M1009_d 8.56368e-19 $X=0.765 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_213 N_A_32_368#_c_205_n N_VGND_M1009_d 0.00257106f $X=0.435 $Y=0.775
+ $X2=-0.19 $Y2=-0.245
cc_214 N_A_32_368#_c_205_n N_VGND_c_482_n 0.0124903f $X=0.435 $Y=0.775 $X2=0
+ $Y2=0
cc_215 N_A_32_368#_M1002_g N_VGND_c_483_n 0.0042292f $X=2.43 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A_32_368#_c_205_n N_VGND_c_486_n 0.00797936f $X=0.435 $Y=0.775 $X2=0
+ $Y2=0
cc_217 N_A_32_368#_M1002_g N_VGND_c_489_n 0.00434272f $X=2.43 $Y=0.74 $X2=0
+ $Y2=0
cc_218 N_A_32_368#_M1002_g N_VGND_c_491_n 0.00822841f $X=2.43 $Y=0.74 $X2=0
+ $Y2=0
cc_219 N_A_32_368#_c_205_n N_VGND_c_491_n 0.0179874f $X=0.435 $Y=0.775 $X2=0
+ $Y2=0
cc_220 N_A1_M1010_g N_A2_M1006_g 0.0375784f $X=2.86 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A1_c_295_n N_A2_M1006_g 0.019932f $X=2.88 $Y=1.425 $X2=0 $Y2=0
cc_222 N_A1_c_296_n N_A2_M1006_g 0.00865654f $X=2.88 $Y=1.425 $X2=0 $Y2=0
cc_223 N_A1_c_294_n N_A2_c_339_n 0.0139686f $X=2.895 $Y=1.795 $X2=0 $Y2=0
cc_224 N_A1_c_298_n N_A2_c_339_n 0.0324651f $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_225 N_A1_c_296_n A2 0.0270452f $X=2.88 $Y=1.425 $X2=0 $Y2=0
cc_226 N_A1_c_298_n N_VPWR_c_366_n 0.0104376f $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_227 N_A1_c_298_n N_VPWR_c_369_n 0.00413917f $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_228 N_A1_c_298_n N_VPWR_c_363_n 0.0081781f $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_229 N_A1_c_298_n N_A_504_392#_c_462_n 0.0134661f $X=2.895 $Y=1.885 $X2=0
+ $Y2=0
cc_230 N_A1_c_295_n N_A_504_392#_c_462_n 2.97896e-19 $X=2.88 $Y=1.425 $X2=0
+ $Y2=0
cc_231 N_A1_c_296_n N_A_504_392#_c_462_n 0.0204706f $X=2.88 $Y=1.425 $X2=0 $Y2=0
cc_232 N_A1_c_298_n N_A_504_392#_c_457_n 7.1333e-19 $X=2.895 $Y=1.885 $X2=0
+ $Y2=0
cc_233 N_A1_c_298_n N_A_504_392#_c_458_n 7.47301e-19 $X=2.895 $Y=1.885 $X2=0
+ $Y2=0
cc_234 N_A1_c_298_n N_A_504_392#_c_459_n 0.00392196f $X=2.895 $Y=1.885 $X2=0
+ $Y2=0
cc_235 N_A1_c_295_n N_A_504_392#_c_459_n 4.92046e-19 $X=2.88 $Y=1.425 $X2=0
+ $Y2=0
cc_236 N_A1_c_296_n N_A_504_392#_c_459_n 0.0016565f $X=2.88 $Y=1.425 $X2=0 $Y2=0
cc_237 N_A1_M1010_g N_VGND_c_485_n 0.00277908f $X=2.86 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A1_M1010_g N_VGND_c_489_n 0.00434272f $X=2.86 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A1_M1010_g N_VGND_c_491_n 0.00821825f $X=2.86 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A2_c_339_n N_VPWR_c_366_n 0.00531445f $X=3.345 $Y=1.885 $X2=0 $Y2=0
cc_241 N_A2_c_339_n N_VPWR_c_370_n 0.00445602f $X=3.345 $Y=1.885 $X2=0 $Y2=0
cc_242 N_A2_c_339_n N_VPWR_c_363_n 0.00861134f $X=3.345 $Y=1.885 $X2=0 $Y2=0
cc_243 N_A2_c_339_n N_A_504_392#_c_462_n 0.0160489f $X=3.345 $Y=1.885 $X2=0
+ $Y2=0
cc_244 N_A2_c_339_n N_A_504_392#_c_457_n 0.00608162f $X=3.345 $Y=1.885 $X2=0
+ $Y2=0
cc_245 A2 N_A_504_392#_c_457_n 0.0277331f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_246 N_A2_c_339_n N_A_504_392#_c_458_n 0.00916896f $X=3.345 $Y=1.885 $X2=0
+ $Y2=0
cc_247 N_A2_M1006_g N_VGND_c_485_n 0.0203366f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A2_c_339_n N_VGND_c_485_n 0.0019397f $X=3.345 $Y=1.885 $X2=0 $Y2=0
cc_249 A2 N_VGND_c_485_n 0.0126785f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_250 N_A2_M1006_g N_VGND_c_489_n 0.00383152f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A2_M1006_g N_VGND_c_491_n 0.00757998f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_252 N_VPWR_M1008_d N_A_504_392#_c_462_n 0.00484629f $X=2.97 $Y=1.96 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_366_n N_A_504_392#_c_462_n 0.0154669f $X=3.12 $Y=2.71 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_366_n N_A_504_392#_c_458_n 0.0362371f $X=3.12 $Y=2.71 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_370_n N_A_504_392#_c_458_n 0.0145938f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_256 N_VPWR_c_363_n N_A_504_392#_c_458_n 0.0120466f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_257 N_VPWR_c_366_n N_A_504_392#_c_459_n 0.0344602f $X=3.12 $Y=2.71 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_369_n N_A_504_392#_c_459_n 0.00749631f $X=2.955 $Y=3.33 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_363_n N_A_504_392#_c_459_n 0.0062048f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_260 N_X_c_421_n N_VGND_M1009_d 0.00215131f $X=1.105 $Y=1.04 $X2=-0.19
+ $Y2=-0.245
cc_261 N_X_c_422_n N_VGND_M1009_d 6.05713e-19 $X=1.105 $Y=1.82 $X2=-0.19
+ $Y2=-0.245
cc_262 N_X_c_421_n N_VGND_c_482_n 0.0157951f $X=1.105 $Y=1.04 $X2=0 $Y2=0
cc_263 N_X_c_421_n N_VGND_c_483_n 0.0160262f $X=1.105 $Y=1.04 $X2=0 $Y2=0
cc_264 N_X_c_421_n N_VGND_c_488_n 0.0147221f $X=1.105 $Y=1.04 $X2=0 $Y2=0
cc_265 N_X_c_421_n N_VGND_c_491_n 0.0180091f $X=1.105 $Y=1.04 $X2=0 $Y2=0
