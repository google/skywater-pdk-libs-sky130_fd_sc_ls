* File: sky130_fd_sc_ls__and2b_1.pex.spice
* Created: Wed Sep  2 10:54:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__AND2B_1%A_N 3 5 7 9 10 11 15 16
c36 16 0 4.13644e-20 $X=0.385 $Y=1.515
r37 15 18 26.3791 $w=3.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.395 $Y=1.515
+ $X2=0.395 $Y2=1.675
r38 15 17 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.395 $Y=1.515
+ $X2=0.395 $Y2=1.35
r39 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.515 $X2=0.385 $Y2=1.515
r40 10 11 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=2.035
r41 10 16 4.06745 $w=4.23e-07 $l=1.5e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.515
r42 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.225 $Y=1.765
+ $X2=1.225 $Y2=2.26
r43 6 18 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.57 $Y=1.675
+ $X2=0.395 $Y2=1.675
r44 5 7 26.9307 $w=1.5e-07 $l=1.27279e-07 $layer=POLY_cond $X=1.135 $Y=1.675
+ $X2=1.225 $Y2=1.765
r45 5 6 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.135 $Y=1.675
+ $X2=0.57 $Y2=1.675
r46 3 17 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.495 $Y=0.645
+ $X2=0.495 $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_LS__AND2B_1%A_27_74# 1 2 7 10 11 13 14 16 17 20 22 26 27
+ 29 31 32
c68 32 0 1.84498e-19 $X=0.975 $Y=1.195
c69 11 0 3.93999e-20 $X=1.675 $Y=1.765
r70 32 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.975 $Y=1.195
+ $X2=0.975 $Y2=1.285
r71 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.195 $X2=0.975 $Y2=1.195
r72 29 34 3.40825 $w=3.3e-07 $l=1.70895e-07 $layer=LI1_cond $X=0.975 $Y=2.32
+ $X2=0.987 $Y2=2.485
r73 29 31 39.2878 $w=3.28e-07 $l=1.125e-06 $layer=LI1_cond $X=0.975 $Y=2.32
+ $X2=0.975 $Y2=1.195
r74 28 31 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.975 $Y=1.18
+ $X2=0.975 $Y2=1.195
r75 26 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.81 $Y=1.095
+ $X2=0.975 $Y2=1.18
r76 26 27 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.81 $Y=1.095
+ $X2=0.445 $Y2=1.095
r77 22 34 3.40825 $w=3.3e-07 $l=1.77e-07 $layer=LI1_cond $X=0.81 $Y=2.485
+ $X2=0.987 $Y2=2.485
r78 22 24 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.81 $Y=2.485
+ $X2=0.64 $Y2=2.485
r79 18 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r80 18 20 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.645
r81 14 17 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.69 $Y=1.21
+ $X2=1.675 $Y2=1.285
r82 14 16 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.69 $Y=1.21 $X2=1.69
+ $Y2=0.81
r83 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.675 $Y=1.765
+ $X2=1.675 $Y2=2.26
r84 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.675 $Y=1.675
+ $X2=1.675 $Y2=1.765
r85 9 17 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.675 $Y=1.36
+ $X2=1.675 $Y2=1.285
r86 9 10 122.444 $w=1.8e-07 $l=3.15e-07 $layer=POLY_cond $X=1.675 $Y=1.36
+ $X2=1.675 $Y2=1.675
r87 8 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.285
+ $X2=0.975 $Y2=1.285
r88 7 17 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.585 $Y=1.285
+ $X2=1.675 $Y2=1.285
r89 7 8 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.585 $Y=1.285
+ $X2=1.14 $Y2=1.285
r90 2 34 600 $w=1.7e-07 $l=1.14287e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=1 $Y2=2.485
r91 2 24 300 $w=1.7e-07 $l=8.61249e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.64 $Y2=2.485
r92 1 20 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LS__AND2B_1%B 3 5 7 8 12
c34 12 0 3.93999e-20 $X=2.21 $Y=1.515
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.515 $X2=2.21 $Y2=1.515
r36 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.21 $Y=1.665
+ $X2=2.21 $Y2=1.515
r37 5 11 50.9845 $w=3.31e-07 $l=2.80624e-07 $layer=POLY_cond $X=2.125 $Y=1.765
+ $X2=2.19 $Y2=1.515
r38 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.125 $Y=1.765
+ $X2=2.125 $Y2=2.26
r39 1 11 38.6069 $w=3.31e-07 $l=2.13014e-07 $layer=POLY_cond $X=2.08 $Y=1.35
+ $X2=2.19 $Y2=1.515
r40 1 3 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.08 $Y=1.35 $X2=2.08
+ $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LS__AND2B_1%A_266_98# 1 2 7 9 12 16 22 23 25 30 31 35
c73 31 0 1.43133e-19 $X=1.885 $Y=1.95
r74 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.75
+ $Y=1.485 $X2=2.75 $Y2=1.485
r75 32 35 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.66 $Y=1.485 $X2=2.75
+ $Y2=1.485
r76 30 31 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=2.115
+ $X2=1.885 $Y2=1.95
r77 25 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.66 $Y=1.32
+ $X2=2.66 $Y2=1.485
r78 24 25 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.66 $Y=1.15
+ $X2=2.66 $Y2=1.32
r79 23 28 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=1.065
+ $X2=1.79 $Y2=1.065
r80 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=1.065
+ $X2=2.66 $Y2=1.15
r81 22 23 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.575 $Y=1.065
+ $X2=1.875 $Y2=1.065
r82 18 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=1.15
+ $X2=1.79 $Y2=1.065
r83 18 31 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=1.79 $Y=1.15 $X2=1.79
+ $Y2=1.95
r84 14 28 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.475 $Y=1.065
+ $X2=1.79 $Y2=1.065
r85 14 16 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.475 $Y=0.98
+ $X2=1.475 $Y2=0.635
r86 10 36 38.532 $w=3.09e-07 $l=2.10286e-07 $layer=POLY_cond $X=2.865 $Y=1.32
+ $X2=2.762 $Y2=1.485
r87 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.865 $Y=1.32
+ $X2=2.865 $Y2=0.76
r88 7 36 56.4705 $w=3.09e-07 $l=3.04893e-07 $layer=POLY_cond $X=2.71 $Y=1.765
+ $X2=2.762 $Y2=1.485
r89 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.71 $Y=1.765
+ $X2=2.71 $Y2=2.4
r90 2 30 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=1.75
+ $Y=1.84 $X2=1.9 $Y2=2.115
r91 1 16 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.33
+ $Y=0.49 $X2=1.475 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LS__AND2B_1%VPWR 1 2 9 13 18 19 21 22 23 36 37
r38 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 27 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r43 26 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 23 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 21 33 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.27 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=3.33
+ $X2=2.435 $Y2=3.33
r49 20 36 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.6 $Y=3.33 $X2=3.12
+ $Y2=3.33
r50 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=3.33
+ $X2=2.435 $Y2=3.33
r51 18 30 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 18 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=3.33
+ $X2=1.45 $Y2=3.33
r53 17 33 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.535 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 17 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=3.33
+ $X2=1.45 $Y2=3.33
r55 13 16 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=2.435 $Y=2.045
+ $X2=2.435 $Y2=2.795
r56 11 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=3.245
+ $X2=2.435 $Y2=3.33
r57 11 16 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.435 $Y=3.245
+ $X2=2.435 $Y2=2.795
r58 7 19 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.45 $Y=3.245 $X2=1.45
+ $Y2=3.33
r59 7 9 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=1.45 $Y=3.245
+ $X2=1.45 $Y2=1.985
r60 2 16 600 $w=1.7e-07 $l=1.06604e-06 $layer=licon1_PDIFF $count=1 $X=2.2
+ $Y=1.84 $X2=2.435 $Y2=2.795
r61 2 13 300 $w=1.7e-07 $l=3.21559e-07 $layer=licon1_PDIFF $count=2 $X=2.2
+ $Y=1.84 $X2=2.435 $Y2=2.045
r62 1 9 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.3
+ $Y=1.84 $X2=1.45 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LS__AND2B_1%X 1 2 9 13 14 15 16 31 32 35
r23 31 32 9.42615 $w=4.83e-07 $l=1.65e-07 $layer=LI1_cond $X=3.012 $Y=1.985
+ $X2=3.012 $Y2=1.82
r24 21 35 0.665858 $w=4.83e-07 $l=2.7e-08 $layer=LI1_cond $X=3.012 $Y=2.062
+ $X2=3.012 $Y2=2.035
r25 16 28 0.986456 $w=4.83e-07 $l=4e-08 $layer=LI1_cond $X=3.012 $Y=2.775
+ $X2=3.012 $Y2=2.815
r26 15 16 9.12472 $w=4.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.012 $Y=2.405
+ $X2=3.012 $Y2=2.775
r27 14 35 0.715181 $w=4.83e-07 $l=2.9e-08 $layer=LI1_cond $X=3.012 $Y=2.006
+ $X2=3.012 $Y2=2.035
r28 14 31 0.51789 $w=4.83e-07 $l=2.1e-08 $layer=LI1_cond $X=3.012 $Y=2.006
+ $X2=3.012 $Y2=1.985
r29 14 15 7.74368 $w=4.83e-07 $l=3.14e-07 $layer=LI1_cond $X=3.012 $Y=2.091
+ $X2=3.012 $Y2=2.405
r30 14 21 0.715181 $w=4.83e-07 $l=2.9e-08 $layer=LI1_cond $X=3.012 $Y=2.091
+ $X2=3.012 $Y2=2.062
r31 13 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.17 $Y=1.15
+ $X2=3.17 $Y2=1.82
r32 7 13 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=3.085 $Y=0.98
+ $X2=3.085 $Y2=1.15
r33 7 9 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=3.085 $Y=0.98
+ $X2=3.085 $Y2=0.535
r34 2 31 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.785
+ $Y=1.84 $X2=2.935 $Y2=1.985
r35 2 28 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.785
+ $Y=1.84 $X2=2.935 $Y2=2.815
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.39 $X2=3.08 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LS__AND2B_1%VGND 1 2 9 13 16 18 23 30 31 34 37
r36 38 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r37 37 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r39 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 31 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r41 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r42 28 37 12.7338 $w=1.7e-07 $l=3.08e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.437
+ $Y2=0
r43 28 30 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=3.12
+ $Y2=0
r44 27 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r45 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r46 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r47 24 26 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r48 23 37 12.7338 $w=1.7e-07 $l=3.07e-07 $layer=LI1_cond $X=2.13 $Y=0 $X2=2.437
+ $Y2=0
r49 23 26 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.13 $Y=0 $X2=1.2
+ $Y2=0
r50 21 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r51 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r52 18 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r53 18 20 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r54 16 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r55 16 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r56 11 37 2.57756 $w=6.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.437 $Y=0.085
+ $X2=2.437 $Y2=0
r57 11 13 10.8911 $w=6.13e-07 $l=5.6e-07 $layer=LI1_cond $X=2.437 $Y=0.085
+ $X2=2.437 $Y2=0.645
r58 7 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r59 7 9 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0.595
r60 2 13 182 $w=1.7e-07 $l=5.6723e-07 $layer=licon1_NDIFF $count=1 $X=2.155
+ $Y=0.49 $X2=2.65 $Y2=0.645
r61 2 13 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.155
+ $Y=0.49 $X2=2.295 $Y2=0.645
r62 1 9 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.595
.ends

