* File: sky130_fd_sc_ls__o41ai_2.pxi.spice
* Created: Wed Sep  2 11:23:50 2020
* 
x_PM_SKY130_FD_SC_LS__O41AI_2%B1 N_B1_c_120_n N_B1_M1015_g N_B1_c_121_n
+ N_B1_M1016_g N_B1_c_112_n N_B1_M1003_g N_B1_c_113_n N_B1_c_114_n N_B1_c_115_n
+ N_B1_M1019_g N_B1_c_116_n N_B1_c_117_n N_B1_c_118_n B1 B1 N_B1_c_119_n
+ PM_SKY130_FD_SC_LS__O41AI_2%B1
x_PM_SKY130_FD_SC_LS__O41AI_2%A4 N_A4_c_177_n N_A4_M1011_g N_A4_M1000_g
+ N_A4_c_178_n N_A4_M1017_g N_A4_M1001_g A4 N_A4_c_175_n N_A4_c_176_n
+ PM_SKY130_FD_SC_LS__O41AI_2%A4
x_PM_SKY130_FD_SC_LS__O41AI_2%A3 N_A3_M1004_g N_A3_c_234_n N_A3_M1006_g
+ N_A3_M1005_g N_A3_c_235_n N_A3_M1012_g A3 N_A3_c_232_n N_A3_c_233_n
+ PM_SKY130_FD_SC_LS__O41AI_2%A3
x_PM_SKY130_FD_SC_LS__O41AI_2%A2 N_A2_M1007_g N_A2_c_286_n N_A2_M1002_g
+ N_A2_M1018_g N_A2_c_280_n N_A2_c_288_n N_A2_M1009_g N_A2_c_281_n N_A2_c_282_n
+ N_A2_c_283_n A2 N_A2_c_285_n PM_SKY130_FD_SC_LS__O41AI_2%A2
x_PM_SKY130_FD_SC_LS__O41AI_2%A1 N_A1_c_350_n N_A1_M1008_g N_A1_c_351_n
+ N_A1_c_352_n N_A1_c_356_n N_A1_M1010_g N_A1_c_353_n N_A1_M1013_g N_A1_c_357_n
+ N_A1_M1014_g A1 A1 N_A1_c_355_n PM_SKY130_FD_SC_LS__O41AI_2%A1
x_PM_SKY130_FD_SC_LS__O41AI_2%VPWR N_VPWR_M1015_s N_VPWR_M1016_s N_VPWR_M1010_d
+ N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_406_n N_VPWR_c_407_n VPWR
+ N_VPWR_c_408_n N_VPWR_c_409_n N_VPWR_c_410_n N_VPWR_c_403_n N_VPWR_c_412_n
+ N_VPWR_c_413_n PM_SKY130_FD_SC_LS__O41AI_2%VPWR
x_PM_SKY130_FD_SC_LS__O41AI_2%Y N_Y_M1003_s N_Y_M1015_d N_Y_M1011_d N_Y_c_473_n
+ N_Y_c_474_n N_Y_c_475_n N_Y_c_470_n N_Y_c_498_n N_Y_c_471_n Y Y
+ PM_SKY130_FD_SC_LS__O41AI_2%Y
x_PM_SKY130_FD_SC_LS__O41AI_2%A_314_368# N_A_314_368#_M1011_s
+ N_A_314_368#_M1017_s N_A_314_368#_M1012_s N_A_314_368#_c_522_n
+ N_A_314_368#_c_523_n N_A_314_368#_c_524_n N_A_314_368#_c_533_n
+ N_A_314_368#_c_536_n N_A_314_368#_c_540_n N_A_314_368#_c_525_n
+ PM_SKY130_FD_SC_LS__O41AI_2%A_314_368#
x_PM_SKY130_FD_SC_LS__O41AI_2%A_607_368# N_A_607_368#_M1006_d
+ N_A_607_368#_M1002_d N_A_607_368#_c_571_n N_A_607_368#_c_569_n
+ N_A_607_368#_c_570_n N_A_607_368#_c_589_p
+ PM_SKY130_FD_SC_LS__O41AI_2%A_607_368#
x_PM_SKY130_FD_SC_LS__O41AI_2%A_807_368# N_A_807_368#_M1002_s
+ N_A_807_368#_M1009_s N_A_807_368#_M1014_s N_A_807_368#_c_599_n
+ N_A_807_368#_c_594_n N_A_807_368#_c_614_n N_A_807_368#_c_595_n
+ N_A_807_368#_c_596_n N_A_807_368#_c_597_n N_A_807_368#_c_609_n
+ PM_SKY130_FD_SC_LS__O41AI_2%A_807_368#
x_PM_SKY130_FD_SC_LS__O41AI_2%A_132_74# N_A_132_74#_M1003_d N_A_132_74#_M1019_d
+ N_A_132_74#_M1001_d N_A_132_74#_M1005_s N_A_132_74#_M1018_d
+ N_A_132_74#_M1013_d N_A_132_74#_c_641_n N_A_132_74#_c_642_n
+ N_A_132_74#_c_643_n N_A_132_74#_c_666_n N_A_132_74#_c_644_n
+ N_A_132_74#_c_645_n N_A_132_74#_c_646_n N_A_132_74#_c_647_n
+ N_A_132_74#_c_648_n N_A_132_74#_c_649_n N_A_132_74#_c_650_n
+ N_A_132_74#_c_651_n N_A_132_74#_c_652_n N_A_132_74#_c_653_n
+ N_A_132_74#_c_654_n N_A_132_74#_c_655_n PM_SKY130_FD_SC_LS__O41AI_2%A_132_74#
x_PM_SKY130_FD_SC_LS__O41AI_2%VGND N_VGND_M1000_s N_VGND_M1004_d N_VGND_M1007_s
+ N_VGND_M1008_s N_VGND_c_739_n N_VGND_c_740_n N_VGND_c_741_n N_VGND_c_742_n
+ N_VGND_c_743_n VGND N_VGND_c_744_n N_VGND_c_745_n N_VGND_c_746_n
+ N_VGND_c_747_n N_VGND_c_748_n N_VGND_c_749_n N_VGND_c_750_n N_VGND_c_751_n
+ N_VGND_c_752_n PM_SKY130_FD_SC_LS__O41AI_2%VGND
cc_1 VNB N_B1_c_112_n 0.0171093f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.22
cc_2 VNB N_B1_c_113_n 0.0249789f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.295
cc_3 VNB N_B1_c_114_n 0.0801735f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.295
cc_4 VNB N_B1_c_115_n 0.0165423f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.22
cc_5 VNB N_B1_c_116_n 0.0207396f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.18
cc_6 VNB N_B1_c_117_n 0.00249471f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.445
cc_7 VNB N_B1_c_118_n 0.126101f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.445
cc_8 VNB N_B1_c_119_n 0.00506713f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.385
cc_9 VNB N_A4_M1000_g 0.0249123f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_10 VNB N_A4_M1001_g 0.0248722f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=0.74
cc_11 VNB N_A4_c_175_n 0.0572219f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.125
cc_12 VNB N_A4_c_176_n 0.0042113f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_13 VNB N_A3_M1004_g 0.023979f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_14 VNB N_A3_M1005_g 0.023493f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.295
cc_15 VNB N_A3_c_232_n 0.00144259f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.125
cc_16 VNB N_A3_c_233_n 0.0339998f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.125
cc_17 VNB N_A2_M1007_g 0.0258128f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_18 VNB N_A2_M1018_g 0.0255771f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.295
cc_19 VNB N_A2_c_280_n 0.0150084f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.22
cc_20 VNB N_A2_c_281_n 0.00917539f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.445
cc_21 VNB N_A2_c_282_n 0.0186415f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.445
cc_22 VNB N_A2_c_283_n 0.011298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB A2 0.00394594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A2_c_285_n 0.00634113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_c_350_n 0.0153172f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_26 VNB N_A1_c_351_n 0.0150084f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.765
cc_27 VNB N_A1_c_352_n 0.00811352f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_28 VNB N_A1_c_353_n 0.0191321f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=0.74
cc_29 VNB A1 0.0162419f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.445
cc_30 VNB N_A1_c_355_n 0.0896288f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.125
cc_31 VNB N_VPWR_c_403_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_470_n 0.00339034f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.125
cc_33 VNB N_Y_c_471_n 0.00758498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB Y 0.00183105f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.22
cc_35 VNB N_A_132_74#_c_641_n 0.00407315f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.125
cc_36 VNB N_A_132_74#_c_642_n 0.0049117f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_37 VNB N_A_132_74#_c_643_n 0.0042908f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_38 VNB N_A_132_74#_c_644_n 0.00596568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_132_74#_c_645_n 0.00444342f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.125
cc_40 VNB N_A_132_74#_c_646_n 0.00252769f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.492
cc_41 VNB N_A_132_74#_c_647_n 0.00443579f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.385
cc_42 VNB N_A_132_74#_c_648_n 0.00234642f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_43 VNB N_A_132_74#_c_649_n 0.00323083f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.365
cc_44 VNB N_A_132_74#_c_650_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_132_74#_c_651_n 0.0145494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_132_74#_c_652_n 0.0281704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_132_74#_c_653_n 0.00446657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_132_74#_c_654_n 0.0103855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_132_74#_c_655_n 0.00194064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_739_n 0.0053606f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.18
cc_51 VNB N_VGND_c_740_n 0.00273364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_741_n 0.00823296f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_53 VNB N_VGND_c_742_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_743_n 0.00571618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_744_n 0.0528354f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.492
cc_56 VNB N_VGND_c_745_n 0.0167762f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.365
cc_57 VNB N_VGND_c_746_n 0.0176545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_747_n 0.0296539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_748_n 0.361198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_749_n 0.00615422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_750_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_751_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_752_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VPB N_B1_c_120_n 0.018686f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_65 VPB N_B1_c_121_n 0.0173788f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_66 VPB N_B1_c_114_n 0.0170446f $X=-0.19 $Y=1.66 $X2=1.095 $Y2=1.295
cc_67 VPB N_A4_c_177_n 0.017024f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_68 VPB N_A4_c_178_n 0.0157017f $X=-0.19 $Y=1.66 $X2=1.02 $Y2=0.74
cc_69 VPB N_A4_c_175_n 0.0199377f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.125
cc_70 VPB N_A4_c_176_n 0.00362871f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_71 VPB N_A3_c_234_n 0.0163877f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_72 VPB N_A3_c_235_n 0.0189067f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.22
cc_73 VPB N_A3_c_232_n 0.00280044f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.125
cc_74 VPB N_A3_c_233_n 0.0215083f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.125
cc_75 VPB N_A2_c_286_n 0.0189603f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_76 VPB N_A2_c_280_n 0.0128229f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.22
cc_77 VPB N_A2_c_288_n 0.0159156f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=0.74
cc_78 VPB N_A2_c_281_n 0.00944818f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.445
cc_79 VPB N_A2_c_282_n 0.0148433f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.445
cc_80 VPB N_A2_c_283_n 0.00537823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB A2 0.00315823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A1_c_356_n 0.0158584f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_83 VPB N_A1_c_357_n 0.0208611f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.22
cc_84 VPB A1 0.0103954f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.445
cc_85 VPB N_A1_c_355_n 0.0268073f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.125
cc_86 VPB N_VPWR_c_404_n 0.0116916f $X=-0.19 $Y=1.66 $X2=1.375 $Y2=1.295
cc_87 VPB N_VPWR_c_405_n 0.0558665f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.22
cc_88 VPB N_VPWR_c_406_n 0.0141083f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.445
cc_89 VPB N_VPWR_c_407_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.125
cc_90 VPB N_VPWR_c_408_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_409_n 0.0997305f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=1.492
cc_92 VPB N_VPWR_c_410_n 0.0197879f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=1.365
cc_93 VPB N_VPWR_c_403_n 0.09416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_412_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_413_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_Y_c_473_n 0.00180921f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.22
cc_97 VPB N_Y_c_474_n 8.2974e-19 $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.445
cc_98 VPB N_Y_c_475_n 0.00267017f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.445
cc_99 VPB N_Y_c_471_n 0.00875991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB Y 0.00506644f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=1.22
cc_101 VPB N_A_314_368#_c_522_n 0.00787077f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.22
cc_102 VPB N_A_314_368#_c_523_n 0.0057859f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=0.74
cc_103 VPB N_A_314_368#_c_524_n 0.00425971f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.18
cc_104 VPB N_A_314_368#_c_525_n 0.00763687f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=1.22
cc_105 VPB N_A_607_368#_c_569_n 0.0197091f $X=-0.19 $Y=1.66 $X2=1.095 $Y2=1.295
cc_106 VPB N_A_607_368#_c_570_n 0.00171072f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.22
cc_107 VPB N_A_807_368#_c_594_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.445
cc_108 VPB N_A_807_368#_c_595_n 0.00802076f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.125
cc_109 VPB N_A_807_368#_c_596_n 0.0357063f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.125
cc_110 VPB N_A_807_368#_c_597_n 0.00889141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 N_B1_c_115_n N_A4_M1000_g 0.0238637f $X=1.45 $Y=1.22 $X2=0 $Y2=0
cc_112 N_B1_c_113_n N_A4_c_175_n 0.00104192f $X=1.375 $Y=1.295 $X2=0 $Y2=0
cc_113 N_B1_c_120_n N_VPWR_c_405_n 0.0182126f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_114 N_B1_c_121_n N_VPWR_c_405_n 6.87691e-19 $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_115 N_B1_c_114_n N_VPWR_c_405_n 0.00263517f $X=1.095 $Y=1.295 $X2=0 $Y2=0
cc_116 N_B1_c_116_n N_VPWR_c_405_n 0.0252545f $X=0.29 $Y=1.18 $X2=0 $Y2=0
cc_117 N_B1_c_120_n N_VPWR_c_406_n 6.05899e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_118 N_B1_c_121_n N_VPWR_c_406_n 0.0184383f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_119 N_B1_c_114_n N_VPWR_c_406_n 7.47062e-19 $X=1.095 $Y=1.295 $X2=0 $Y2=0
cc_120 N_B1_c_120_n N_VPWR_c_408_n 0.00413917f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_121 N_B1_c_121_n N_VPWR_c_408_n 0.00413917f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_122 N_B1_c_120_n N_VPWR_c_403_n 0.00817726f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_123 N_B1_c_121_n N_VPWR_c_403_n 0.00817726f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_124 N_B1_c_120_n N_Y_c_473_n 0.00374174f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_125 N_B1_c_121_n N_Y_c_473_n 0.0064943f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_126 N_B1_c_121_n N_Y_c_474_n 0.0115681f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_127 N_B1_c_114_n N_Y_c_474_n 0.0104714f $X=1.095 $Y=1.295 $X2=0 $Y2=0
cc_128 N_B1_c_119_n N_Y_c_474_n 0.00699753f $X=0.735 $Y=1.385 $X2=0 $Y2=0
cc_129 N_B1_c_120_n N_Y_c_475_n 0.00212373f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_130 N_B1_c_114_n N_Y_c_475_n 0.00353119f $X=1.095 $Y=1.295 $X2=0 $Y2=0
cc_131 N_B1_c_119_n N_Y_c_475_n 0.0144515f $X=0.735 $Y=1.385 $X2=0 $Y2=0
cc_132 N_B1_c_112_n N_Y_c_470_n 0.0104314f $X=1.02 $Y=1.22 $X2=0 $Y2=0
cc_133 N_B1_c_113_n N_Y_c_470_n 0.0159874f $X=1.375 $Y=1.295 $X2=0 $Y2=0
cc_134 N_B1_c_114_n N_Y_c_470_n 0.00863317f $X=1.095 $Y=1.295 $X2=0 $Y2=0
cc_135 N_B1_c_115_n N_Y_c_470_n 0.00916866f $X=1.45 $Y=1.22 $X2=0 $Y2=0
cc_136 N_B1_c_117_n N_Y_c_470_n 0.00437927f $X=0.29 $Y=0.445 $X2=0 $Y2=0
cc_137 N_B1_c_118_n N_Y_c_470_n 7.61813e-19 $X=0.29 $Y=0.445 $X2=0 $Y2=0
cc_138 N_B1_c_119_n N_Y_c_470_n 0.0302432f $X=0.735 $Y=1.385 $X2=0 $Y2=0
cc_139 N_B1_c_113_n N_Y_c_471_n 0.00548316f $X=1.375 $Y=1.295 $X2=0 $Y2=0
cc_140 N_B1_c_114_n Y 0.00695651f $X=1.095 $Y=1.295 $X2=0 $Y2=0
cc_141 N_B1_c_116_n Y 0.00253276f $X=0.29 $Y=1.18 $X2=0 $Y2=0
cc_142 N_B1_c_121_n N_A_314_368#_c_522_n 0.0017837f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_B1_c_121_n N_A_314_368#_c_524_n 5.80628e-19 $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_144 N_B1_c_114_n N_A_132_74#_c_641_n 0.0012734f $X=1.095 $Y=1.295 $X2=0 $Y2=0
cc_145 N_B1_c_117_n N_A_132_74#_c_641_n 0.0424601f $X=0.29 $Y=0.445 $X2=0 $Y2=0
cc_146 N_B1_c_118_n N_A_132_74#_c_641_n 0.00586749f $X=0.29 $Y=0.445 $X2=0 $Y2=0
cc_147 N_B1_c_119_n N_A_132_74#_c_641_n 0.0216688f $X=0.735 $Y=1.385 $X2=0 $Y2=0
cc_148 N_B1_c_112_n N_A_132_74#_c_642_n 0.0125991f $X=1.02 $Y=1.22 $X2=0 $Y2=0
cc_149 N_B1_c_115_n N_A_132_74#_c_642_n 0.0134151f $X=1.45 $Y=1.22 $X2=0 $Y2=0
cc_150 N_B1_c_117_n N_A_132_74#_c_643_n 0.0114723f $X=0.29 $Y=0.445 $X2=0 $Y2=0
cc_151 N_B1_c_118_n N_A_132_74#_c_643_n 0.00158635f $X=0.29 $Y=0.445 $X2=0 $Y2=0
cc_152 N_B1_c_115_n N_A_132_74#_c_645_n 0.00116009f $X=1.45 $Y=1.22 $X2=0 $Y2=0
cc_153 N_B1_c_112_n N_VGND_c_744_n 0.00278271f $X=1.02 $Y=1.22 $X2=0 $Y2=0
cc_154 N_B1_c_115_n N_VGND_c_744_n 0.00278271f $X=1.45 $Y=1.22 $X2=0 $Y2=0
cc_155 N_B1_c_117_n N_VGND_c_744_n 0.0191905f $X=0.29 $Y=0.445 $X2=0 $Y2=0
cc_156 N_B1_c_118_n N_VGND_c_744_n 0.00683346f $X=0.29 $Y=0.445 $X2=0 $Y2=0
cc_157 N_B1_c_112_n N_VGND_c_748_n 0.00358427f $X=1.02 $Y=1.22 $X2=0 $Y2=0
cc_158 N_B1_c_115_n N_VGND_c_748_n 0.0035414f $X=1.45 $Y=1.22 $X2=0 $Y2=0
cc_159 N_B1_c_117_n N_VGND_c_748_n 0.012382f $X=0.29 $Y=0.445 $X2=0 $Y2=0
cc_160 N_B1_c_118_n N_VGND_c_748_n 0.00469111f $X=0.29 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A4_M1001_g N_A3_M1004_g 0.0242448f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A4_c_178_n N_A3_c_234_n 0.0175322f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A4_c_175_n N_A3_c_232_n 3.49546e-19 $X=2.45 $Y=1.557 $X2=0 $Y2=0
cc_164 N_A4_c_176_n N_A3_c_232_n 0.0261548f $X=2.495 $Y=1.515 $X2=0 $Y2=0
cc_165 N_A4_c_175_n N_A3_c_233_n 0.0235416f $X=2.45 $Y=1.557 $X2=0 $Y2=0
cc_166 N_A4_c_176_n N_A3_c_233_n 0.00347328f $X=2.495 $Y=1.515 $X2=0 $Y2=0
cc_167 N_A4_c_177_n N_VPWR_c_406_n 0.00264796f $X=1.925 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A4_c_177_n N_VPWR_c_409_n 0.00278257f $X=1.925 $Y=1.765 $X2=0 $Y2=0
cc_169 N_A4_c_178_n N_VPWR_c_409_n 0.00278257f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A4_c_177_n N_VPWR_c_403_n 0.00358623f $X=1.925 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A4_c_178_n N_VPWR_c_403_n 0.00354984f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A4_M1000_g N_Y_c_470_n 9.84918e-19 $X=1.95 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A4_c_175_n N_Y_c_470_n 0.00613813f $X=2.45 $Y=1.557 $X2=0 $Y2=0
cc_174 N_A4_c_178_n N_Y_c_498_n 0.00461325f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_175 N_A4_c_177_n N_Y_c_471_n 0.012072f $X=1.925 $Y=1.765 $X2=0 $Y2=0
cc_176 N_A4_c_178_n N_Y_c_471_n 0.00336536f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A4_c_175_n N_Y_c_471_n 0.0273814f $X=2.45 $Y=1.557 $X2=0 $Y2=0
cc_178 N_A4_c_176_n N_Y_c_471_n 0.019097f $X=2.495 $Y=1.515 $X2=0 $Y2=0
cc_179 N_A4_c_177_n N_A_314_368#_c_522_n 0.0136157f $X=1.925 $Y=1.765 $X2=0
+ $Y2=0
cc_180 N_A4_c_178_n N_A_314_368#_c_522_n 6.12174e-19 $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_181 N_A4_c_177_n N_A_314_368#_c_523_n 0.0108414f $X=1.925 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A4_c_178_n N_A_314_368#_c_523_n 0.0127176f $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A4_c_177_n N_A_314_368#_c_524_n 0.00262934f $X=1.925 $Y=1.765 $X2=0
+ $Y2=0
cc_184 N_A4_c_178_n N_A_314_368#_c_533_n 0.00193523f $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A4_c_175_n N_A_314_368#_c_533_n 0.00109032f $X=2.45 $Y=1.557 $X2=0
+ $Y2=0
cc_186 N_A4_c_176_n N_A_314_368#_c_533_n 0.0256132f $X=2.495 $Y=1.515 $X2=0
+ $Y2=0
cc_187 N_A4_c_177_n N_A_314_368#_c_536_n 6.22492e-19 $X=1.925 $Y=1.765 $X2=0
+ $Y2=0
cc_188 N_A4_c_178_n N_A_314_368#_c_536_n 0.00919154f $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_A4_M1000_g N_A_132_74#_c_642_n 0.00346618f $X=1.95 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A4_M1000_g N_A_132_74#_c_666_n 0.00862682f $X=1.95 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A4_M1001_g N_A_132_74#_c_666_n 0.00103499f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A4_M1000_g N_A_132_74#_c_644_n 0.0124437f $X=1.95 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A4_M1001_g N_A_132_74#_c_644_n 0.0145948f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A4_c_175_n N_A_132_74#_c_644_n 0.00507755f $X=2.45 $Y=1.557 $X2=0 $Y2=0
cc_195 N_A4_c_176_n N_A_132_74#_c_644_n 0.0129287f $X=2.495 $Y=1.515 $X2=0 $Y2=0
cc_196 N_A4_M1000_g N_A_132_74#_c_645_n 0.00177665f $X=1.95 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A4_c_175_n N_A_132_74#_c_645_n 0.00116995f $X=2.45 $Y=1.557 $X2=0 $Y2=0
cc_198 N_A4_M1001_g N_A_132_74#_c_646_n 4.64401e-19 $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A4_c_175_n N_A_132_74#_c_653_n 6.33179e-19 $X=2.45 $Y=1.557 $X2=0 $Y2=0
cc_200 N_A4_c_176_n N_A_132_74#_c_653_n 0.0154186f $X=2.495 $Y=1.515 $X2=0 $Y2=0
cc_201 N_A4_M1000_g N_VGND_c_739_n 0.00358845f $X=1.95 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A4_M1001_g N_VGND_c_739_n 0.00993236f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A4_M1001_g N_VGND_c_740_n 4.40104e-19 $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A4_M1000_g N_VGND_c_744_n 0.00430908f $X=1.95 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A4_M1001_g N_VGND_c_745_n 0.00383152f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A4_M1000_g N_VGND_c_748_n 0.00816828f $X=1.95 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A4_M1001_g N_VGND_c_748_n 0.0075821f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A3_M1005_g N_A2_M1007_g 0.0123368f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A3_c_232_n N_A2_c_281_n 7.15378e-19 $X=3.29 $Y=1.515 $X2=0 $Y2=0
cc_210 N_A3_c_233_n N_A2_c_281_n 0.0222324f $X=3.38 $Y=1.557 $X2=0 $Y2=0
cc_211 N_A3_c_232_n N_A2_c_285_n 0.0165751f $X=3.29 $Y=1.515 $X2=0 $Y2=0
cc_212 N_A3_c_233_n N_A2_c_285_n 8.82993e-19 $X=3.38 $Y=1.557 $X2=0 $Y2=0
cc_213 N_A3_c_234_n N_VPWR_c_409_n 0.0044313f $X=2.96 $Y=1.765 $X2=0 $Y2=0
cc_214 N_A3_c_235_n N_VPWR_c_409_n 0.00278271f $X=3.41 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A3_c_234_n N_VPWR_c_403_n 0.00855285f $X=2.96 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A3_c_235_n N_VPWR_c_403_n 0.00358624f $X=3.41 $Y=1.765 $X2=0 $Y2=0
cc_217 N_A3_c_234_n N_A_314_368#_c_523_n 0.0017442f $X=2.96 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A3_c_234_n N_A_314_368#_c_536_n 0.0103412f $X=2.96 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A3_c_234_n N_A_314_368#_c_540_n 0.0191394f $X=2.96 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A3_c_235_n N_A_314_368#_c_540_n 0.0123917f $X=3.41 $Y=1.765 $X2=0 $Y2=0
cc_221 N_A3_c_232_n N_A_314_368#_c_540_n 0.0306997f $X=3.29 $Y=1.515 $X2=0 $Y2=0
cc_222 N_A3_c_233_n N_A_314_368#_c_540_n 0.00130895f $X=3.38 $Y=1.557 $X2=0
+ $Y2=0
cc_223 N_A3_c_234_n N_A_314_368#_c_525_n 7.3898e-19 $X=2.96 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A3_c_235_n N_A_314_368#_c_525_n 0.00993868f $X=3.41 $Y=1.765 $X2=0
+ $Y2=0
cc_225 N_A3_c_234_n N_A_607_368#_c_571_n 0.00736507f $X=2.96 $Y=1.765 $X2=0
+ $Y2=0
cc_226 N_A3_c_235_n N_A_607_368#_c_569_n 0.0147555f $X=3.41 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A3_c_234_n N_A_607_368#_c_570_n 0.00351848f $X=2.96 $Y=1.765 $X2=0
+ $Y2=0
cc_228 N_A3_c_235_n N_A_807_368#_c_597_n 0.00335288f $X=3.41 $Y=1.765 $X2=0
+ $Y2=0
cc_229 N_A3_M1004_g N_A_132_74#_c_646_n 0.00349332f $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A3_M1004_g N_A_132_74#_c_647_n 0.0187835f $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A3_M1005_g N_A_132_74#_c_647_n 0.0132161f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A3_c_232_n N_A_132_74#_c_647_n 0.0339034f $X=3.29 $Y=1.515 $X2=0 $Y2=0
cc_233 N_A3_c_233_n N_A_132_74#_c_647_n 0.00382903f $X=3.38 $Y=1.557 $X2=0 $Y2=0
cc_234 N_A3_M1005_g N_A_132_74#_c_648_n 4.30451e-19 $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A3_M1004_g N_VGND_c_739_n 4.50471e-19 $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A3_M1004_g N_VGND_c_740_n 0.0094116f $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A3_M1005_g N_VGND_c_740_n 0.00995981f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A3_M1004_g N_VGND_c_745_n 0.00398535f $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A3_M1005_g N_VGND_c_746_n 0.00383152f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A3_M1004_g N_VGND_c_748_n 0.00788205f $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A3_M1005_g N_VGND_c_748_n 0.0075791f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A2_M1018_g N_A1_c_350_n 0.0202553f $X=4.41 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_243 A2 N_A1_c_351_n 0.00369725f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_244 N_A2_c_280_n N_A1_c_352_n 0.00933586f $X=4.755 $Y=1.65 $X2=0 $Y2=0
cc_245 N_A2_c_285_n N_A1_c_352_n 0.00369725f $X=4.925 $Y=1.565 $X2=0 $Y2=0
cc_246 N_A2_c_288_n N_A1_c_356_n 0.0123235f $X=4.845 $Y=1.765 $X2=0 $Y2=0
cc_247 A2 A1 0.0337104f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_248 N_A2_M1018_g N_A1_c_355_n 0.00248938f $X=4.41 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A2_c_280_n N_A1_c_355_n 0.00859121f $X=4.755 $Y=1.65 $X2=0 $Y2=0
cc_250 A2 N_A1_c_355_n 0.00564956f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_251 N_A2_c_286_n N_VPWR_c_409_n 0.00278271f $X=4.395 $Y=1.765 $X2=0 $Y2=0
cc_252 N_A2_c_288_n N_VPWR_c_409_n 0.00445602f $X=4.845 $Y=1.765 $X2=0 $Y2=0
cc_253 N_A2_c_286_n N_VPWR_c_403_n 0.00358624f $X=4.395 $Y=1.765 $X2=0 $Y2=0
cc_254 N_A2_c_288_n N_VPWR_c_403_n 0.00858435f $X=4.845 $Y=1.765 $X2=0 $Y2=0
cc_255 N_A2_c_286_n N_A_314_368#_c_525_n 0.00135275f $X=4.395 $Y=1.765 $X2=0
+ $Y2=0
cc_256 N_A2_c_281_n N_A_314_368#_c_525_n 9.44376e-19 $X=3.915 $Y=1.537 $X2=0
+ $Y2=0
cc_257 N_A2_c_285_n N_A_314_368#_c_525_n 0.00209089f $X=4.925 $Y=1.565 $X2=0
+ $Y2=0
cc_258 N_A2_c_286_n N_A_607_368#_c_569_n 0.0144245f $X=4.395 $Y=1.765 $X2=0
+ $Y2=0
cc_259 N_A2_c_288_n N_A_607_368#_c_569_n 0.00341066f $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_260 N_A2_c_286_n N_A_807_368#_c_599_n 0.012525f $X=4.395 $Y=1.765 $X2=0 $Y2=0
cc_261 N_A2_c_280_n N_A_807_368#_c_599_n 0.00482685f $X=4.755 $Y=1.65 $X2=0
+ $Y2=0
cc_262 N_A2_c_288_n N_A_807_368#_c_599_n 0.012432f $X=4.845 $Y=1.765 $X2=0 $Y2=0
cc_263 N_A2_c_285_n N_A_807_368#_c_599_n 0.0258073f $X=4.925 $Y=1.565 $X2=0
+ $Y2=0
cc_264 N_A2_c_286_n N_A_807_368#_c_594_n 6.54425e-19 $X=4.395 $Y=1.765 $X2=0
+ $Y2=0
cc_265 N_A2_c_288_n N_A_807_368#_c_594_n 0.0103267f $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_266 N_A2_c_286_n N_A_807_368#_c_597_n 0.013251f $X=4.395 $Y=1.765 $X2=0 $Y2=0
cc_267 N_A2_c_288_n N_A_807_368#_c_597_n 0.00104667f $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_268 N_A2_c_282_n N_A_807_368#_c_597_n 0.00761339f $X=4.305 $Y=1.537 $X2=0
+ $Y2=0
cc_269 N_A2_c_285_n N_A_807_368#_c_597_n 0.0246245f $X=4.925 $Y=1.565 $X2=0
+ $Y2=0
cc_270 N_A2_c_288_n N_A_807_368#_c_609_n 4.74495e-19 $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_271 A2 N_A_807_368#_c_609_n 0.0179976f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_272 N_A2_c_285_n N_A_807_368#_c_609_n 9.00871e-19 $X=4.925 $Y=1.565 $X2=0
+ $Y2=0
cc_273 N_A2_M1007_g N_A_132_74#_c_648_n 0.0100056f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A2_M1018_g N_A_132_74#_c_648_n 7.61734e-19 $X=4.41 $Y=0.74 $X2=0 $Y2=0
cc_275 N_A2_M1007_g N_A_132_74#_c_649_n 0.0118691f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A2_M1018_g N_A_132_74#_c_649_n 0.0118691f $X=4.41 $Y=0.74 $X2=0 $Y2=0
cc_277 N_A2_c_282_n N_A_132_74#_c_649_n 0.00552458f $X=4.305 $Y=1.537 $X2=0
+ $Y2=0
cc_278 N_A2_c_285_n N_A_132_74#_c_649_n 0.049279f $X=4.925 $Y=1.565 $X2=0 $Y2=0
cc_279 N_A2_M1007_g N_A_132_74#_c_650_n 7.60766e-19 $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A2_M1018_g N_A_132_74#_c_650_n 0.0101129f $X=4.41 $Y=0.74 $X2=0 $Y2=0
cc_281 N_A2_c_285_n N_A_132_74#_c_651_n 0.0287688f $X=4.925 $Y=1.565 $X2=0 $Y2=0
cc_282 N_A2_M1007_g N_A_132_74#_c_654_n 0.00162843f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A2_c_285_n N_A_132_74#_c_654_n 0.00199562f $X=4.925 $Y=1.565 $X2=0
+ $Y2=0
cc_284 N_A2_M1018_g N_A_132_74#_c_655_n 0.00155819f $X=4.41 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A2_c_280_n N_A_132_74#_c_655_n 0.00136108f $X=4.755 $Y=1.65 $X2=0 $Y2=0
cc_286 N_A2_c_285_n N_A_132_74#_c_655_n 0.0288617f $X=4.925 $Y=1.565 $X2=0 $Y2=0
cc_287 N_A2_M1007_g N_VGND_c_740_n 5.00531e-19 $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_288 N_A2_M1007_g N_VGND_c_741_n 0.00452037f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_289 N_A2_M1018_g N_VGND_c_741_n 0.00457079f $X=4.41 $Y=0.74 $X2=0 $Y2=0
cc_290 N_A2_M1018_g N_VGND_c_742_n 0.00434272f $X=4.41 $Y=0.74 $X2=0 $Y2=0
cc_291 N_A2_M1007_g N_VGND_c_746_n 0.00434272f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_292 N_A2_M1007_g N_VGND_c_748_n 0.00821664f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_293 N_A2_M1018_g N_VGND_c_748_n 0.00821391f $X=4.41 $Y=0.74 $X2=0 $Y2=0
cc_294 N_A1_c_356_n N_VPWR_c_407_n 0.00486623f $X=5.295 $Y=1.765 $X2=0 $Y2=0
cc_295 N_A1_c_357_n N_VPWR_c_407_n 0.00486623f $X=5.745 $Y=1.765 $X2=0 $Y2=0
cc_296 N_A1_c_356_n N_VPWR_c_409_n 0.00445602f $X=5.295 $Y=1.765 $X2=0 $Y2=0
cc_297 N_A1_c_357_n N_VPWR_c_410_n 0.00445602f $X=5.745 $Y=1.765 $X2=0 $Y2=0
cc_298 N_A1_c_356_n N_VPWR_c_403_n 0.00857673f $X=5.295 $Y=1.765 $X2=0 $Y2=0
cc_299 N_A1_c_357_n N_VPWR_c_403_n 0.0086105f $X=5.745 $Y=1.765 $X2=0 $Y2=0
cc_300 N_A1_c_356_n N_A_807_368#_c_594_n 0.0103374f $X=5.295 $Y=1.765 $X2=0
+ $Y2=0
cc_301 N_A1_c_357_n N_A_807_368#_c_594_n 6.45594e-19 $X=5.745 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_A1_c_356_n N_A_807_368#_c_614_n 0.0154891f $X=5.295 $Y=1.765 $X2=0
+ $Y2=0
cc_303 N_A1_c_357_n N_A_807_368#_c_614_n 0.0120074f $X=5.745 $Y=1.765 $X2=0
+ $Y2=0
cc_304 A1 N_A_807_368#_c_614_n 0.0310306f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_305 N_A1_c_355_n N_A_807_368#_c_614_n 0.00130963f $X=5.745 $Y=1.475 $X2=0
+ $Y2=0
cc_306 N_A1_c_357_n N_A_807_368#_c_595_n 4.27055e-19 $X=5.745 $Y=1.765 $X2=0
+ $Y2=0
cc_307 A1 N_A_807_368#_c_595_n 0.0247152f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_308 N_A1_c_355_n N_A_807_368#_c_595_n 0.0010282f $X=5.745 $Y=1.475 $X2=0
+ $Y2=0
cc_309 N_A1_c_356_n N_A_807_368#_c_596_n 6.45594e-19 $X=5.295 $Y=1.765 $X2=0
+ $Y2=0
cc_310 N_A1_c_357_n N_A_807_368#_c_596_n 0.0104891f $X=5.745 $Y=1.765 $X2=0
+ $Y2=0
cc_311 N_A1_c_351_n N_A_807_368#_c_609_n 0.0010207f $X=5.205 $Y=1.26 $X2=0 $Y2=0
cc_312 N_A1_c_356_n N_A_807_368#_c_609_n 9.50925e-19 $X=5.295 $Y=1.765 $X2=0
+ $Y2=0
cc_313 N_A1_c_350_n N_A_132_74#_c_650_n 0.00998742f $X=4.84 $Y=1.185 $X2=0 $Y2=0
cc_314 N_A1_c_353_n N_A_132_74#_c_650_n 7.48402e-19 $X=5.34 $Y=1.185 $X2=0 $Y2=0
cc_315 N_A1_c_350_n N_A_132_74#_c_651_n 0.0109137f $X=4.84 $Y=1.185 $X2=0 $Y2=0
cc_316 N_A1_c_351_n N_A_132_74#_c_651_n 0.00432085f $X=5.205 $Y=1.26 $X2=0 $Y2=0
cc_317 N_A1_c_353_n N_A_132_74#_c_651_n 0.0189246f $X=5.34 $Y=1.185 $X2=0 $Y2=0
cc_318 A1 N_A_132_74#_c_651_n 0.0364957f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_319 N_A1_c_355_n N_A_132_74#_c_651_n 0.0118315f $X=5.745 $Y=1.475 $X2=0 $Y2=0
cc_320 N_A1_c_353_n N_A_132_74#_c_652_n 0.0128452f $X=5.34 $Y=1.185 $X2=0 $Y2=0
cc_321 N_A1_c_350_n N_A_132_74#_c_655_n 0.0014099f $X=4.84 $Y=1.185 $X2=0 $Y2=0
cc_322 N_A1_c_350_n N_VGND_c_742_n 0.00434272f $X=4.84 $Y=1.185 $X2=0 $Y2=0
cc_323 N_A1_c_350_n N_VGND_c_743_n 0.00409384f $X=4.84 $Y=1.185 $X2=0 $Y2=0
cc_324 N_A1_c_353_n N_VGND_c_743_n 0.0126272f $X=5.34 $Y=1.185 $X2=0 $Y2=0
cc_325 N_A1_c_353_n N_VGND_c_747_n 0.00383152f $X=5.34 $Y=1.185 $X2=0 $Y2=0
cc_326 N_A1_c_350_n N_VGND_c_748_n 0.00820816f $X=4.84 $Y=1.185 $X2=0 $Y2=0
cc_327 N_A1_c_353_n N_VGND_c_748_n 0.00762539f $X=5.34 $Y=1.185 $X2=0 $Y2=0
cc_328 N_VPWR_c_405_n N_Y_c_473_n 0.0709943f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_329 N_VPWR_c_406_n N_Y_c_473_n 0.0599532f $X=1.17 $Y=2.225 $X2=0 $Y2=0
cc_330 N_VPWR_c_408_n N_Y_c_473_n 0.00749631f $X=1.005 $Y=3.33 $X2=0 $Y2=0
cc_331 N_VPWR_c_403_n N_Y_c_473_n 0.0062048f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_332 N_VPWR_c_406_n N_Y_c_474_n 0.00102433f $X=1.17 $Y=2.225 $X2=0 $Y2=0
cc_333 N_VPWR_c_405_n N_Y_c_475_n 0.00513432f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_334 N_VPWR_M1016_s Y 0.00270301f $X=1.02 $Y=1.84 $X2=0 $Y2=0
cc_335 N_VPWR_c_406_n Y 0.0232918f $X=1.17 $Y=2.225 $X2=0 $Y2=0
cc_336 N_VPWR_c_406_n N_A_314_368#_c_522_n 0.0627384f $X=1.17 $Y=2.225 $X2=0
+ $Y2=0
cc_337 N_VPWR_c_409_n N_A_314_368#_c_523_n 0.0594839f $X=5.435 $Y=3.33 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_403_n N_A_314_368#_c_523_n 0.0329562f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_339 N_VPWR_c_406_n N_A_314_368#_c_524_n 0.0134078f $X=1.17 $Y=2.225 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_409_n N_A_314_368#_c_524_n 0.0236039f $X=5.435 $Y=3.33 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_403_n N_A_314_368#_c_524_n 0.012761f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_342 N_VPWR_c_409_n N_A_607_368#_c_569_n 0.0927443f $X=5.435 $Y=3.33 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_403_n N_A_607_368#_c_569_n 0.0527972f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_344 N_VPWR_c_409_n N_A_607_368#_c_570_n 0.017869f $X=5.435 $Y=3.33 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_403_n N_A_607_368#_c_570_n 0.00965079f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_346 N_VPWR_c_407_n N_A_807_368#_c_594_n 0.0449718f $X=5.52 $Y=2.455 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_409_n N_A_807_368#_c_594_n 0.014552f $X=5.435 $Y=3.33 $X2=0
+ $Y2=0
cc_348 N_VPWR_c_403_n N_A_807_368#_c_594_n 0.0119791f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_349 N_VPWR_M1010_d N_A_807_368#_c_614_n 0.00408911f $X=5.37 $Y=1.84 $X2=0
+ $Y2=0
cc_350 N_VPWR_c_407_n N_A_807_368#_c_614_n 0.0136682f $X=5.52 $Y=2.455 $X2=0
+ $Y2=0
cc_351 N_VPWR_c_407_n N_A_807_368#_c_596_n 0.0449718f $X=5.52 $Y=2.455 $X2=0
+ $Y2=0
cc_352 N_VPWR_c_410_n N_A_807_368#_c_596_n 0.0145938f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_353 N_VPWR_c_403_n N_A_807_368#_c_596_n 0.0120466f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_354 N_Y_c_471_n N_A_314_368#_M1011_s 0.00265217f $X=2.035 $Y=1.72 $X2=-0.19
+ $Y2=-0.245
cc_355 N_Y_c_471_n N_A_314_368#_c_522_n 0.0231236f $X=2.035 $Y=1.72 $X2=0 $Y2=0
cc_356 N_Y_M1011_d N_A_314_368#_c_523_n 0.00218679f $X=2 $Y=1.84 $X2=0 $Y2=0
cc_357 N_Y_c_498_n N_A_314_368#_c_523_n 0.013472f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_358 N_Y_c_498_n N_A_314_368#_c_533_n 0.0119113f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_359 N_Y_c_498_n N_A_314_368#_c_536_n 0.0405146f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_360 N_Y_M1003_s N_A_132_74#_c_642_n 0.00197509f $X=1.095 $Y=0.37 $X2=0 $Y2=0
cc_361 N_Y_c_470_n N_A_132_74#_c_642_n 0.0127602f $X=1.235 $Y=0.81 $X2=0 $Y2=0
cc_362 N_Y_c_471_n N_A_132_74#_c_644_n 0.0140717f $X=2.035 $Y=1.72 $X2=0 $Y2=0
cc_363 N_Y_c_470_n N_A_132_74#_c_645_n 0.00962585f $X=1.235 $Y=0.81 $X2=0 $Y2=0
cc_364 N_Y_c_471_n N_A_132_74#_c_645_n 0.0166545f $X=2.035 $Y=1.72 $X2=0 $Y2=0
cc_365 N_A_314_368#_c_540_n N_A_607_368#_M1006_d 0.00384138f $X=3.47 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_366 N_A_314_368#_c_536_n N_A_607_368#_c_571_n 0.03423f $X=2.6 $Y=2.815 $X2=0
+ $Y2=0
cc_367 N_A_314_368#_c_540_n N_A_607_368#_c_571_n 0.0154248f $X=3.47 $Y=2.035
+ $X2=0 $Y2=0
cc_368 N_A_314_368#_c_525_n N_A_607_368#_c_571_n 0.0298377f $X=3.635 $Y=2.115
+ $X2=0 $Y2=0
cc_369 N_A_314_368#_M1012_s N_A_607_368#_c_569_n 0.00266942f $X=3.485 $Y=1.84
+ $X2=0 $Y2=0
cc_370 N_A_314_368#_c_525_n N_A_607_368#_c_569_n 0.0206198f $X=3.635 $Y=2.115
+ $X2=0 $Y2=0
cc_371 N_A_314_368#_c_523_n N_A_607_368#_c_570_n 0.0110653f $X=2.435 $Y=2.99
+ $X2=0 $Y2=0
cc_372 N_A_314_368#_c_525_n N_A_807_368#_c_597_n 0.058783f $X=3.635 $Y=2.115
+ $X2=0 $Y2=0
cc_373 N_A_607_368#_c_569_n N_A_807_368#_M1002_s 0.00273752f $X=4.535 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_374 N_A_607_368#_M1002_d N_A_807_368#_c_599_n 0.00438683f $X=4.47 $Y=1.84
+ $X2=0 $Y2=0
cc_375 N_A_607_368#_c_589_p N_A_807_368#_c_599_n 0.0136682f $X=4.62 $Y=2.455
+ $X2=0 $Y2=0
cc_376 N_A_607_368#_c_569_n N_A_807_368#_c_594_n 0.00549849f $X=4.535 $Y=2.99
+ $X2=0 $Y2=0
cc_377 N_A_607_368#_c_589_p N_A_807_368#_c_594_n 0.040027f $X=4.62 $Y=2.455
+ $X2=0 $Y2=0
cc_378 N_A_607_368#_c_569_n N_A_807_368#_c_597_n 0.0206053f $X=4.535 $Y=2.99
+ $X2=0 $Y2=0
cc_379 N_A_607_368#_c_589_p N_A_807_368#_c_597_n 0.0289859f $X=4.62 $Y=2.455
+ $X2=0 $Y2=0
cc_380 N_A_132_74#_c_644_n N_VGND_M1000_s 0.00277863f $X=2.58 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_381 N_A_132_74#_c_647_n N_VGND_M1004_d 0.00201333f $X=3.51 $Y=1.095 $X2=0
+ $Y2=0
cc_382 N_A_132_74#_c_649_n N_VGND_M1007_s 0.00393158f $X=4.46 $Y=1.095 $X2=0
+ $Y2=0
cc_383 N_A_132_74#_c_651_n N_VGND_M1008_s 0.00277863f $X=5.46 $Y=1.095 $X2=0
+ $Y2=0
cc_384 N_A_132_74#_c_642_n N_VGND_c_739_n 0.011924f $X=1.57 $Y=0.34 $X2=0 $Y2=0
cc_385 N_A_132_74#_c_644_n N_VGND_c_739_n 0.0176026f $X=2.58 $Y=1.095 $X2=0
+ $Y2=0
cc_386 N_A_132_74#_c_646_n N_VGND_c_739_n 0.0166774f $X=2.665 $Y=0.515 $X2=0
+ $Y2=0
cc_387 N_A_132_74#_c_646_n N_VGND_c_740_n 0.0174554f $X=2.665 $Y=0.515 $X2=0
+ $Y2=0
cc_388 N_A_132_74#_c_647_n N_VGND_c_740_n 0.0143251f $X=3.51 $Y=1.095 $X2=0
+ $Y2=0
cc_389 N_A_132_74#_c_648_n N_VGND_c_740_n 0.01669f $X=3.61 $Y=0.515 $X2=0 $Y2=0
cc_390 N_A_132_74#_c_648_n N_VGND_c_741_n 0.0170729f $X=3.61 $Y=0.515 $X2=0
+ $Y2=0
cc_391 N_A_132_74#_c_649_n N_VGND_c_741_n 0.0209063f $X=4.46 $Y=1.095 $X2=0
+ $Y2=0
cc_392 N_A_132_74#_c_650_n N_VGND_c_741_n 0.017488f $X=4.625 $Y=0.515 $X2=0
+ $Y2=0
cc_393 N_A_132_74#_c_650_n N_VGND_c_742_n 0.0144922f $X=4.625 $Y=0.515 $X2=0
+ $Y2=0
cc_394 N_A_132_74#_c_650_n N_VGND_c_743_n 0.017488f $X=4.625 $Y=0.515 $X2=0
+ $Y2=0
cc_395 N_A_132_74#_c_651_n N_VGND_c_743_n 0.0176026f $X=5.46 $Y=1.095 $X2=0
+ $Y2=0
cc_396 N_A_132_74#_c_652_n N_VGND_c_743_n 0.017488f $X=5.625 $Y=0.515 $X2=0
+ $Y2=0
cc_397 N_A_132_74#_c_642_n N_VGND_c_744_n 0.0664416f $X=1.57 $Y=0.34 $X2=0 $Y2=0
cc_398 N_A_132_74#_c_643_n N_VGND_c_744_n 0.0179217f $X=0.89 $Y=0.34 $X2=0 $Y2=0
cc_399 N_A_132_74#_c_646_n N_VGND_c_745_n 0.011066f $X=2.665 $Y=0.515 $X2=0
+ $Y2=0
cc_400 N_A_132_74#_c_648_n N_VGND_c_746_n 0.0123329f $X=3.61 $Y=0.515 $X2=0
+ $Y2=0
cc_401 N_A_132_74#_c_652_n N_VGND_c_747_n 0.0146357f $X=5.625 $Y=0.515 $X2=0
+ $Y2=0
cc_402 N_A_132_74#_c_642_n N_VGND_c_748_n 0.0369085f $X=1.57 $Y=0.34 $X2=0 $Y2=0
cc_403 N_A_132_74#_c_643_n N_VGND_c_748_n 0.00971942f $X=0.89 $Y=0.34 $X2=0
+ $Y2=0
cc_404 N_A_132_74#_c_646_n N_VGND_c_748_n 0.00915947f $X=2.665 $Y=0.515 $X2=0
+ $Y2=0
cc_405 N_A_132_74#_c_648_n N_VGND_c_748_n 0.0101517f $X=3.61 $Y=0.515 $X2=0
+ $Y2=0
cc_406 N_A_132_74#_c_650_n N_VGND_c_748_n 0.0118826f $X=4.625 $Y=0.515 $X2=0
+ $Y2=0
cc_407 N_A_132_74#_c_652_n N_VGND_c_748_n 0.0121141f $X=5.625 $Y=0.515 $X2=0
+ $Y2=0
