* NGSPICE file created from sky130_fd_sc_ls__decap_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__decap_4 VGND VNB VPB VPWR
M1000 VPWR VGND VPWR VPB phighvt w=1e+06u l=1e+06u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1001 VGND VPWR VGND VNB nshort w=420000u l=1e+06u
+  ad=2.352e+11p pd=2.8e+06u as=0p ps=0u
.ends

