* File: sky130_fd_sc_ls__clkbuf_4.spice
* Created: Wed Sep  2 10:57:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__clkbuf_4.pex.spice"
.subckt sky130_fd_sc_ls__clkbuf_4  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_83_270#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_83_270#_M1004_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1004_d N_A_83_270#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_83_270#_M1009_g N_X_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.0672 PD=0.8 PS=0.74 NRD=8.568 NRS=11.424 M=1 R=2.8 SA=75001.5
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1003 N_A_83_270#_M1003_d N_A_M1003_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.126 AS=0.0798 PD=1.44 PS=0.8 NRD=1.428 NRS=19.992 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_83_270#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_A_83_270#_M1005_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1005_d N_A_83_270#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1007_d N_A_83_270#_M1007_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1002 N_A_83_270#_M1002_d N_A_M1002_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ls__clkbuf_4.pxi.spice"
*
.ends
*
*
