* File: sky130_fd_sc_ls__einvp_8.spice
* Created: Wed Sep  2 11:07:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__einvp_8.pex.spice"
.subckt sky130_fd_sc_ls__einvp_8  VNB VPB A TE Z VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Z	Z
* TE	TE
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_A_27_74#_M1005_d N_A_M1005_g N_Z_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75007.2 A=0.111 P=1.78 MULT=1
MM1009 N_A_27_74#_M1009_d N_A_M1009_g N_Z_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75006.8 A=0.111 P=1.78 MULT=1
MM1014 N_A_27_74#_M1009_d N_A_M1014_g N_Z_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75006.3 A=0.111 P=1.78 MULT=1
MM1016 N_A_27_74#_M1016_d N_A_M1016_g N_Z_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75005.8 A=0.111 P=1.78 MULT=1
MM1020 N_A_27_74#_M1016_d N_A_M1020_g N_Z_M1020_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.1
+ SB=75005.3 A=0.111 P=1.78 MULT=1
MM1023 N_A_27_74#_M1023_d N_A_M1023_g N_Z_M1020_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75004.8 A=0.111 P=1.78 MULT=1
MM1026 N_A_27_74#_M1023_d N_A_M1026_g N_Z_M1026_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.1
+ SB=75004.3 A=0.111 P=1.78 MULT=1
MM1027 N_A_27_74#_M1027_d N_A_M1027_g N_Z_M1026_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75003.8 A=0.111 P=1.78 MULT=1
MM1004 N_A_27_74#_M1027_d N_TE_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.1
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1012 N_A_27_74#_M1012_d N_TE_M1012_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75004.6
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1015 N_A_27_74#_M1012_d N_TE_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1017 N_A_27_74#_M1017_d N_TE_M1017_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.4
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1024 N_A_27_74#_M1017_d N_TE_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.9
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1029 N_A_27_74#_M1029_d N_TE_M1029_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1030 N_A_27_74#_M1029_d N_TE_M1030_g N_VGND_M1030_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75006.7
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1032 N_A_27_74#_M1032_d N_TE_M1032_g N_VGND_M1030_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75007.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1033 N_VGND_M1033_d N_TE_M1033_g N_A_802_323#_M1033_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.2146 PD=2.05 PS=2.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_27_368#_M1000_d N_A_M1000_g N_Z_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3248 AS=0.168 PD=2.82 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75007 A=0.168 P=2.54 MULT=1
MM1003 N_A_27_368#_M1003_d N_A_M1003_g N_Z_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75006.5 A=0.168 P=2.54 MULT=1
MM1010 N_A_27_368#_M1003_d N_A_M1010_g N_Z_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75006.1 A=0.168 P=2.54 MULT=1
MM1018 N_A_27_368#_M1018_d N_A_M1018_g N_Z_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75005.6 A=0.168 P=2.54 MULT=1
MM1021 N_A_27_368#_M1018_d N_A_M1021_g N_Z_M1021_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75005.2 A=0.168 P=2.54 MULT=1
MM1022 N_A_27_368#_M1022_d N_A_M1022_g N_Z_M1021_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75004.7 A=0.168 P=2.54 MULT=1
MM1025 N_A_27_368#_M1022_d N_A_M1025_g N_Z_M1025_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.9 SB=75004.3 A=0.168 P=2.54 MULT=1
MM1031 N_A_27_368#_M1031_d N_A_M1031_g N_Z_M1025_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.4 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1001 N_A_27_368#_M1031_d N_A_802_323#_M1001_g N_VPWR_M1001_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75003.8 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1002 N_A_27_368#_M1002_d N_A_802_323#_M1002_g N_VPWR_M1001_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75004.3 SB=75002.9 A=0.168 P=2.54 MULT=1
MM1006 N_A_27_368#_M1002_d N_A_802_323#_M1006_g N_VPWR_M1006_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75004.7 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1007 N_A_27_368#_M1007_d N_A_802_323#_M1007_g N_VPWR_M1006_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75005.2 SB=75002 A=0.168 P=2.54 MULT=1
MM1008 N_A_27_368#_M1007_d N_A_802_323#_M1008_g N_VPWR_M1008_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75005.6 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1011 N_A_27_368#_M1011_d N_A_802_323#_M1011_g N_VPWR_M1008_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75006.1 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1019 N_A_27_368#_M1011_d N_A_802_323#_M1019_g N_VPWR_M1019_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75006.5 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1028 N_A_27_368#_M1028_d N_A_802_323#_M1028_g N_VPWR_M1019_s VPB PHIGHVT
+ L=0.15 W=1.12 AD=0.3248 AS=0.168 PD=2.82 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75007 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1013_d N_TE_M1013_g N_A_802_323#_M1013_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3192 AS=0.3192 PD=2.81 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX34_noxref VNB VPB NWDIODE A=17.67 P=22.72
*
.include "sky130_fd_sc_ls__einvp_8.pxi.spice"
*
.ends
*
*
