* File: sky130_fd_sc_ls__o21ai_2.spice
* Created: Wed Sep  2 11:18:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o21ai_2.pex.spice"
.subckt sky130_fd_sc_ls__o21ai_2  VNB VPB A1 A2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1008 N_A_27_74#_M1008_d N_A1_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1003 N_A_27_74#_M1003_d N_A2_M1003_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.74
+ AD=0.10915 AS=0.1295 PD=1.035 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1011 N_A_27_74#_M1003_d N_A2_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.10915 AS=0.12395 PD=1.035 PS=1.075 NRD=2.424 NRS=8.916 M=1 R=4.93333
+ SA=75001.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1010 N_A_27_74#_M1010_d N_A1_M1010_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.74
+ AD=0.12025 AS=0.12395 PD=1.065 PS=1.075 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_A_27_74#_M1010_d VNB NSHORT L=0.15 W=0.74
+ AD=0.11655 AS=0.12025 PD=1.055 PS=1.065 NRD=4.86 NRS=7.296 M=1 R=4.93333
+ SA=75002.1 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1002_d N_B1_M1005_g N_A_27_74#_M1005_s VNB NSHORT L=0.15 W=0.74
+ AD=0.11655 AS=0.2109 PD=1.055 PS=2.05 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_116_368#_M1000_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1007_d N_A2_M1007_g N_A_116_368#_M1000_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1009 N_Y_M1007_d N_A2_M1009_g N_A_116_368#_M1009_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_116_368#_M1009_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1001_d N_B1_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ls__o21ai_2.pxi.spice"
*
.ends
*
*
