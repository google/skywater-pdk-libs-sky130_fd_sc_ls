# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__nor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__nor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 1.795000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.180000 4.195000 1.550000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.793600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.640000 0.340000 1.690000 0.840000 ;
        RECT 0.640000 0.840000 2.690000 1.010000 ;
        RECT 2.360000 0.350000 2.690000 0.840000 ;
        RECT 2.360000 1.010000 2.690000 1.130000 ;
        RECT 2.365000 1.130000 2.690000 1.180000 ;
        RECT 2.365000 1.180000 2.755000 1.410000 ;
        RECT 2.365000 1.410000 2.695000 1.720000 ;
        RECT 2.365000 1.720000 3.695000 1.890000 ;
        RECT 2.365000 1.890000 2.695000 2.735000 ;
        RECT 3.365000 1.890000 3.695000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.085000 0.470000 1.010000 ;
      RECT 0.115000  1.720000 2.195000 1.890000 ;
      RECT 0.115000  1.890000 0.445000 2.980000 ;
      RECT 0.645000  2.060000 0.815000 3.245000 ;
      RECT 1.015000  1.890000 1.345000 2.980000 ;
      RECT 1.545000  2.060000 1.715000 3.245000 ;
      RECT 1.860000  0.085000 2.190000 0.670000 ;
      RECT 1.915000  1.890000 2.195000 2.905000 ;
      RECT 1.915000  2.905000 4.145000 3.075000 ;
      RECT 2.860000  0.085000 4.205000 1.010000 ;
      RECT 2.865000  2.060000 3.195000 2.905000 ;
      RECT 3.865000  1.820000 4.145000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_ls__nor2_4
END LIBRARY
