* File: sky130_fd_sc_ls__a221o_4.spice
* Created: Wed Sep  2 10:49:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__a221o_4.pex.spice"
.subckt sky130_fd_sc_ls__a221o_4  VNB VPB A1 A2 C1 B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* C1	C1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1004 N_A_154_135#_M1004_d N_A1_M1004_g N_A_71_135#_M1004_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1006 N_A_154_135#_M1004_d N_A1_M1006_g N_A_71_135#_M1006_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1022 N_A_71_135#_M1022_d N_A2_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75004.7 A=0.096 P=1.58 MULT=1
MM1026 N_A_71_135#_M1022_d N_A2_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.114423 PD=0.92 PS=1.01565 NRD=0 NRS=12.18 M=1 R=4.26667
+ SA=75000.6 SB=75004.3 A=0.096 P=1.58 MULT=1
MM1003 N_X_M1003_d N_A_154_135#_M1003_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.132302 PD=1.02 PS=1.17435 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1003_d N_A_154_135#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1020 N_X_M1020_d N_A_154_135#_M1020_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1023 N_X_M1020_d N_A_154_135#_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.26817 PD=1.02 PS=1.58725 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1024 N_A_154_135#_M1024_d N_C1_M1024_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.23193 PD=0.92 PS=1.37275 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.3
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1025 N_A_154_135#_M1024_d N_C1_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1648 PD=0.92 PS=1.17 NRD=0 NRS=30.468 M=1 R=4.26667 SA=75003.7
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1015 N_A_1346_123#_M1015_d N_B2_M1015_g N_VGND_M1025_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1648 PD=0.92 PS=1.17 NRD=0 NRS=13.584 M=1 R=4.26667
+ SA=75004.3 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1016 N_A_1346_123#_M1015_d N_B2_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 N_A_154_135#_M1009_d N_B1_M1009_g N_A_1346_123#_M1009_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1019 N_A_154_135#_M1009_d N_B1_M1019_g N_A_1346_123#_M1019_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.2144 PD=0.92 PS=1.95 NRD=0 NRS=4.68 M=1 R=4.26667
+ SA=75000.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1000 N_A_157_376#_M1000_d N_A1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.21 AS=0.275 PD=1.42 PS=2.55 NRD=25.5903 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75004.1 A=0.15 P=2.3 MULT=1
MM1017 N_A_157_376#_M1000_d N_A1_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.21 AS=0.3725 PD=1.42 PS=1.745 NRD=1.9503 NRS=12.7853 M=1 R=6.66667
+ SA=75000.8 SB=75003.5 A=0.15 P=2.3 MULT=1
MM1005 N_A_157_376#_M1005_d N_A2_M1005_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.3725 PD=1.3 PS=1.745 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75001.7 SB=75002.6 A=0.15 P=2.3 MULT=1
MM1010 N_A_157_376#_M1005_d N_A2_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.232547 PD=1.3 PS=1.49057 NRD=1.9503 NRS=34.4553 M=1 R=6.66667
+ SA=75002.1 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1001 N_X_M1001_d N_A_154_135#_M1001_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.260453 PD=1.42 PS=1.66943 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1007 N_X_M1001_d N_A_154_135#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.9 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1011 N_X_M1011_d N_A_154_135#_M1011_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.4 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1018 N_X_M1011_d N_A_154_135#_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.8 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1014 N_A_154_135#_M1014_d N_C1_M1014_g N_A_1102_392#_M1014_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.8 A=0.15 P=2.3 MULT=1
MM1021 N_A_154_135#_M1014_d N_C1_M1021_g N_A_1102_392#_M1021_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.6 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1002 N_A_157_376#_M1002_d N_B2_M1002_g N_A_1102_392#_M1021_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1008 N_A_157_376#_M1002_d N_B2_M1008_g N_A_1102_392#_M1008_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.15 AS=0.295 PD=1.3 PS=1.59 NRD=1.9503 NRS=32.4853 M=1
+ R=6.66667 SA=75001.5 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1012 N_A_157_376#_M1012_d N_B1_M1012_g N_A_1102_392#_M1008_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.17 AS=0.295 PD=1.34 PS=1.59 NRD=5.8903 NRS=28.565 M=1
+ R=6.66667 SA=75002.3 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1027 N_A_157_376#_M1012_d N_B1_M1027_g N_A_1102_392#_M1027_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.17 AS=0.275 PD=1.34 PS=2.55 NRD=5.8903 NRS=1.9503 M=1
+ R=6.66667 SA=75002.8 SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=18.5628 P=23.68
c_158 VPB 0 2.11319e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ls__a221o_4.pxi.spice"
*
.ends
*
*
