* File: sky130_fd_sc_ls__clkinv_2.pex.spice
* Created: Wed Sep  2 10:58:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__CLKINV_2%A 3 5 7 8 10 11 13 16 18 19 20 30
r49 30 31 1.94355 $w=3.72e-07 $l=1.5e-08 $layer=POLY_cond $X=1.41 $Y=1.557
+ $X2=1.425 $Y2=1.557
r50 29 30 58.3064 $w=3.72e-07 $l=4.5e-07 $layer=POLY_cond $X=0.96 $Y=1.557
+ $X2=1.41 $Y2=1.557
r51 27 29 4.53495 $w=3.72e-07 $l=3.5e-08 $layer=POLY_cond $X=0.925 $Y=1.557
+ $X2=0.96 $Y2=1.557
r52 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.925
+ $Y=1.515 $X2=0.925 $Y2=1.515
r53 25 27 53.7715 $w=3.72e-07 $l=4.15e-07 $layer=POLY_cond $X=0.51 $Y=1.557
+ $X2=0.925 $Y2=1.557
r54 24 25 1.94355 $w=3.72e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.51 $Y2=1.557
r55 20 28 7.37028 $w=4.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.925 $Y2=1.565
r56 19 28 5.4942 $w=4.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.925 $Y2=1.565
r57 18 19 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.72 $Y2=1.565
r58 14 31 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=1.557
r59 14 16 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=0.61
r60 11 30 24.0971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.41 $Y2=1.557
r61 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.41 $Y2=2.4
r62 8 29 24.0971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=1.557
r63 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=2.4
r64 5 25 24.0971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.557
r65 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r66 1 24 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r67 1 3 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_2%Y 1 2 3 10 12 14 18 20 22 29 31 34
r49 33 34 32.8196 $w=2.28e-07 $l=6.55e-07 $layer=LI1_cond $X=1.68 $Y=1.95
+ $X2=1.68 $Y2=1.295
r50 32 34 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.18
+ $X2=1.68 $Y2=1.295
r51 27 29 10.6117 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.14 $Y=0.845
+ $X2=1.305 $Y2=0.845
r52 23 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=2.035
+ $X2=1.185 $Y2=2.035
r53 22 33 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.565 $Y=2.035
+ $X2=1.68 $Y2=1.95
r54 22 23 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.565 $Y=2.035
+ $X2=1.35 $Y2=2.035
r55 20 32 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.565 $Y=1.095
+ $X2=1.68 $Y2=1.18
r56 20 29 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.565 $Y=1.095
+ $X2=1.305 $Y2=1.095
r57 16 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.12
+ $X2=1.185 $Y2=2.035
r58 16 18 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.185 $Y=2.12
+ $X2=1.185 $Y2=2.815
r59 15 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=2.035
+ $X2=0.285 $Y2=2.035
r60 14 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=2.035
+ $X2=1.185 $Y2=2.035
r61 14 15 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.02 $Y=2.035
+ $X2=0.45 $Y2=2.035
r62 10 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=2.12
+ $X2=0.285 $Y2=2.035
r63 10 12 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.285 $Y=2.12
+ $X2=0.285 $Y2=2.815
r64 3 31 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.115
r65 3 18 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.815
r66 2 25 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.115
r67 2 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.815
r68 1 27 91 $w=1.7e-07 $l=6.9401e-07 $layer=licon1_NDIFF $count=2 $X=0.57 $Y=0.4
+ $X2=1.14 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_2%VPWR 1 2 11 13 15 17 19 25 29
r28 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 23 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r31 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r32 20 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=0.735 $Y2=3.33
r33 20 22 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=3.33 $X2=1.2
+ $Y2=3.33
r34 19 28 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.55 $Y=3.33
+ $X2=1.735 $Y2=3.33
r35 19 22 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.55 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 17 23 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r37 17 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 13 28 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=1.675 $Y=3.245
+ $X2=1.735 $Y2=3.33
r39 13 15 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=1.675 $Y=3.245
+ $X2=1.675 $Y2=2.455
r40 9 25 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=3.33
r41 9 11 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=2.455
r42 2 15 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.84 $X2=1.635 $Y2=2.455
r43 1 11 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_2%VGND 1 2 7 9 11 13 15 17 27
r18 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r19 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r20 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r21 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r22 18 23 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r23 18 20 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=1.2
+ $Y2=0
r24 17 26 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.697
+ $Y2=0
r25 17 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.2
+ $Y2=0
r26 15 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r27 15 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.24
+ $Y2=0
r28 11 26 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=1.64 $Y=0.085
+ $X2=1.697 $Y2=0
r29 11 13 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=1.64 $Y=0.085
+ $X2=1.64 $Y2=0.61
r30 7 23 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r31 7 9 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.61
r32 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.4 $X2=1.64 $Y2=0.61
r33 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.4 $X2=0.28 $Y2=0.61
.ends

