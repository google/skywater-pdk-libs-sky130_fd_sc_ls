# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__a32o_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__a32o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 2.915000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.015000 1.350000 2.345000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 1.350000 1.775000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.155000 1.350000 3.715000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885000 1.300000 4.215000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.550600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.820000 0.935000 2.150000 ;
        RECT 0.615000 0.330000 0.935000 1.150000 ;
        RECT 0.725000 1.150000 0.935000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.320000 0.085000 ;
        RECT 0.115000  0.085000 0.445000 1.130000 ;
        RECT 1.185000  0.085000 1.515000 0.840000 ;
        RECT 3.850000  0.085000 4.180000 1.130000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 4.320000 3.415000 ;
        RECT 0.115000 2.660000 0.445000 3.245000 ;
        RECT 1.100000 2.660000 1.510000 3.245000 ;
        RECT 2.265000 2.630000 2.645000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.225000 1.320000 0.555000 1.650000 ;
      RECT 0.225000 1.650000 0.395000 2.320000 ;
      RECT 0.225000 2.320000 1.275000 2.490000 ;
      RECT 1.105000 1.010000 3.105000 1.180000 ;
      RECT 1.105000 1.180000 1.275000 1.950000 ;
      RECT 1.105000 1.950000 3.705000 2.120000 ;
      RECT 1.105000 2.120000 1.275000 2.320000 ;
      RECT 1.715000 2.290000 3.205000 2.460000 ;
      RECT 1.715000 2.460000 2.045000 2.860000 ;
      RECT 2.775000 0.350000 3.105000 1.010000 ;
      RECT 2.875000 2.460000 3.205000 2.905000 ;
      RECT 2.875000 2.905000 4.205000 3.075000 ;
      RECT 3.375000 2.120000 3.705000 2.735000 ;
      RECT 3.875000 1.950000 4.205000 2.905000 ;
  END
END sky130_fd_sc_ls__a32o_2
