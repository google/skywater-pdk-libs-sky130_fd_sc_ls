# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__a41oi_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__a41oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.285000 1.350000 3.295000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.320000 5.620000 1.650000 ;
        RECT 3.965000 1.650000 4.675000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.350000 8.035000 1.780000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285000 1.350000 9.955000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.430000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.447600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.350000 0.875000 1.010000 ;
        RECT 0.545000 1.010000 2.435000 1.180000 ;
        RECT 0.615000 1.950000 3.715000 2.120000 ;
        RECT 0.615000 2.120000 0.945000 2.735000 ;
        RECT 1.645000 1.820000 2.105000 1.950000 ;
        RECT 1.645000 2.120000 1.815000 2.735000 ;
        RECT 1.815000 1.180000 2.105000 1.820000 ;
        RECT 2.105000 0.595000 2.435000 1.010000 ;
        RECT 3.305000 0.595000 3.635000 1.000000 ;
        RECT 3.465000 1.000000 3.635000 1.550000 ;
        RECT 3.465000 1.550000 3.715000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.080000 0.085000 ;
        RECT 0.115000  0.085000  0.365000 1.130000 ;
        RECT 1.045000  0.085000  1.375000 0.840000 ;
        RECT 8.305000  0.085000  8.635000 0.840000 ;
        RECT 9.165000  0.085000  9.495000 0.840000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
        RECT 9.755000 -0.085000 9.925000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 10.080000 3.415000 ;
        RECT 2.515000 2.630000  2.845000 3.245000 ;
        RECT 3.545000 2.630000  3.795000 3.245000 ;
        RECT 4.500000 2.290000  4.750000 3.245000 ;
        RECT 5.460000 2.290000  5.710000 3.245000 ;
        RECT 6.410000 2.290000  6.660000 3.245000 ;
        RECT 7.360000 2.290000  7.610000 3.245000 ;
        RECT 8.280000 2.290000  8.530000 3.245000 ;
        RECT 9.260000 2.290000  9.430000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
        RECT 9.755000 3.245000 9.925000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 1.950000 0.445000 2.905000 ;
      RECT 0.115000 2.905000 2.345000 3.075000 ;
      RECT 1.115000 2.290000 1.445000 2.905000 ;
      RECT 1.605000 0.255000 5.925000 0.425000 ;
      RECT 1.605000 0.425000 1.935000 0.840000 ;
      RECT 2.015000 2.290000 4.300000 2.460000 ;
      RECT 2.015000 2.460000 2.345000 2.905000 ;
      RECT 2.605000 0.425000 3.135000 1.130000 ;
      RECT 3.015000 2.460000 3.345000 2.980000 ;
      RECT 3.805000 0.425000 5.925000 0.620000 ;
      RECT 3.805000 0.620000 4.135000 1.130000 ;
      RECT 3.970000 1.950000 9.960000 2.120000 ;
      RECT 3.970000 2.120000 4.300000 2.290000 ;
      RECT 3.970000 2.460000 4.300000 2.980000 ;
      RECT 4.305000 0.790000 7.775000 1.130000 ;
      RECT 4.930000 1.820000 5.260000 1.950000 ;
      RECT 4.930000 2.120000 5.260000 2.980000 ;
      RECT 5.880000 2.120000 6.210000 2.980000 ;
      RECT 6.155000 0.350000 8.125000 0.600000 ;
      RECT 6.155000 0.600000 6.485000 0.620000 ;
      RECT 6.830000 2.120000 7.160000 2.980000 ;
      RECT 7.445000 0.770000 7.775000 0.790000 ;
      RECT 7.780000 2.120000 8.110000 2.980000 ;
      RECT 7.955000 0.600000 8.125000 1.010000 ;
      RECT 7.955000 1.010000 9.965000 1.180000 ;
      RECT 8.730000 2.120000 9.060000 2.980000 ;
      RECT 8.815000 0.350000 8.985000 1.010000 ;
      RECT 9.630000 2.120000 9.960000 2.980000 ;
      RECT 9.715000 0.350000 9.965000 1.010000 ;
  END
END sky130_fd_sc_ls__a41oi_4
