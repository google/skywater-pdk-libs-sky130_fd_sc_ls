* File: sky130_fd_sc_ls__o21ba_1.spice
* Created: Wed Sep  2 11:18:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__o21ba_1.pex.spice"
.subckt sky130_fd_sc_ls__o21ba_1  VNB VPB A1 A2 B1_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1_N	B1_N
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A1_M1007_g N_A_27_74#_M1007_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1344 AS=0.1824 PD=1.06 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1008 N_A_27_74#_M1008_d N_A2_M1008_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0944 AS=0.1344 PD=0.935 PS=1.06 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75000.8
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1003 N_A_200_392#_M1003_d N_A_281_244#_M1003_g N_A_27_74#_M1008_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.2176 AS=0.0944 PD=1.96 PS=0.935 NRD=10.308 NRS=2.808 M=1
+ R=4.26667 SA=75001.2 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1004_d N_B1_N_M1004_g N_A_281_244#_M1004_s VNB NSHORT L=0.15
+ W=0.55 AD=0.123601 AS=0.275 PD=0.989147 PS=2.1 NRD=23.448 NRS=0 M=1 R=3.66667
+ SA=75000.4 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1009 N_X_M1009_d N_A_200_392#_M1009_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.166299 PD=2.05 PS=1.33085 NRD=0 NRS=5.664 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 A_116_392# N_A1_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1002 N_A_200_392#_M1002_d N_A2_M1002_g A_116_392# VPB PHIGHVT L=0.15 W=1
+ AD=0.21 AS=0.135 PD=1.42 PS=1.27 NRD=15.7403 NRS=15.7403 M=1 R=6.66667
+ SA=75000.6 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A_281_244#_M1001_g N_A_200_392#_M1002_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.295 AS=0.21 PD=2.59 PS=1.42 NRD=1.9503 NRS=11.8003 M=1
+ R=6.66667 SA=75001.2 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_B1_N_M1005_g N_A_281_244#_M1005_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.198 AS=0.3108 PD=1.33286 PS=2.42 NRD=42.3747 NRS=3.5066 M=1 R=5.6
+ SA=75000.3 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1000 N_X_M1000_d N_A_200_392#_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.3304 AS=0.264 PD=2.83 PS=1.77714 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ls__o21ba_1.pxi.spice"
*
.ends
*
*
