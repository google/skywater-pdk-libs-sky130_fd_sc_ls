* NGSPICE file created from sky130_fd_sc_ls__nand3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_ls__nand3b_4 A_N B C VGND VNB VPB VPWR Y
M1000 VPWR A_N a_89_172# VPB phighvt w=840000u l=150000u
+  ad=4.9686e+12p pd=1.99e+07u as=2.52e+11p ps=2.28e+06u
M1001 a_744_74# B a_297_82# VNB nshort w=740000u l=150000u
+  ad=1.0672e+12p pd=1.036e+07u as=8.806e+11p ps=8.3e+06u
M1002 Y C VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=1.4336e+12p pd=9.28e+06u as=0p ps=0u
M1003 a_297_82# C VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=1.1492e+12p ps=8.02e+06u
M1004 a_744_74# a_89_172# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=4.329e+11p ps=4.13e+06u
M1005 a_744_74# B a_297_82# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y a_89_172# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR C Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND C a_297_82# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND C a_297_82# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_297_82# C VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y a_89_172# a_744_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_89_172# a_744_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_297_82# B a_744_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_89_172# Y VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_297_82# B a_744_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_89_172# A_N VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_744_74# a_89_172# Y VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A_N a_89_172# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=1.9515e+11p ps=2.05e+06u
.ends

