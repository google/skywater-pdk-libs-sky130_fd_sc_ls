* File: sky130_fd_sc_ls__fa_2.spice
* Created: Fri Aug 28 13:25:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__fa_2.pex.spice"
.subckt sky130_fd_sc_ls__fa_2  VNB VPB A CIN B VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* B	B
* CIN	CIN
* A	A
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_A_M1015_g N_A_27_79#_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.18315 AS=0.2109 PD=1.235 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75008.3 A=0.111 P=1.78 MULT=1
MM1003 N_A_27_79#_M1003_d N_B_M1003_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.74
+ AD=0.2109 AS=0.18315 PD=1.31 PS=1.235 NRD=23.508 NRS=23.508 M=1 R=4.93333
+ SA=75000.9 SB=75007.7 A=0.111 P=1.78 MULT=1
MM1028 N_A_336_347#_M1028_d N_CIN_M1028_g N_A_27_79#_M1003_d VNB NSHORT L=0.15
+ W=0.74 AD=0.1295 AS=0.2109 PD=1.09 PS=1.31 NRD=11.34 NRS=23.508 M=1 R=4.93333
+ SA=75001.6 SB=75007 A=0.111 P=1.78 MULT=1
MM1021 A_487_79# N_B_M1021_g N_A_336_347#_M1028_d VNB NSHORT L=0.15 W=0.74
+ AD=0.0888 AS=0.1295 PD=0.98 PS=1.09 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75006.5 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1019_d N_A_M1019_g A_487_79# VNB NSHORT L=0.15 W=0.74 AD=0.1961
+ AS=0.0888 PD=1.27 PS=0.98 NRD=14.592 NRS=10.536 M=1 R=4.93333 SA=75002.5
+ SB=75006.1 A=0.111 P=1.78 MULT=1
MM1029 N_A_701_79#_M1029_d N_CIN_M1029_g N_VGND_M1019_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=1.27 NRD=0 NRS=25.944 M=1 R=4.93333 SA=75003.1
+ SB=75005.4 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_B_M1011_g N_A_701_79#_M1029_d VNB NSHORT L=0.15 W=0.74
+ AD=0.193975 AS=0.1036 PD=1.395 PS=1.02 NRD=33.588 NRS=0 M=1 R=4.93333
+ SA=75003.6 SB=75005 A=0.111 P=1.78 MULT=1
MM1013 N_A_701_79#_M1013_d N_A_M1013_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1554 AS=0.193975 PD=1.16 PS=1.395 NRD=1.212 NRS=33.588 M=1 R=4.93333
+ SA=75004.2 SB=75004.4 A=0.111 P=1.78 MULT=1
MM1031 N_A_992_347#_M1031_d N_A_336_347#_M1031_g N_A_701_79#_M1013_d VNB NSHORT
+ L=0.15 W=0.74 AD=0.1295 AS=0.1554 PD=1.09 PS=1.16 NRD=11.34 NRS=11.34 M=1
+ R=4.93333 SA=75004.7 SB=75003.8 A=0.111 P=1.78 MULT=1
MM1017 A_1119_79# N_CIN_M1017_g N_A_992_347#_M1031_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=13.776 NRS=0 M=1 R=4.93333 SA=75005.2
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1000 A_1205_79# N_B_M1000_g A_1119_79# VNB NSHORT L=0.15 W=0.74 AD=0.0888
+ AS=0.1036 PD=0.98 PS=1.02 NRD=10.536 NRS=13.776 M=1 R=4.93333 SA=75005.7
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g A_1205_79# VNB NSHORT L=0.15 W=0.74
+ AD=0.253662 AS=0.0888 PD=1.52 PS=0.98 NRD=23.508 NRS=10.536 M=1 R=4.93333
+ SA=75006.1 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1002 N_COUT_M1002_d N_A_336_347#_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.253662 PD=1.02 PS=1.52 NRD=0 NRS=46.668 M=1 R=4.93333
+ SA=75006.8 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1008 N_COUT_M1002_d N_A_336_347#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.251275 PD=1.02 PS=1.515 NRD=0 NRS=46.14 M=1 R=4.93333
+ SA=75007.2 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1004 N_SUM_M1004_d N_A_992_347#_M1004_g N_VGND_M1008_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.251275 PD=1.02 PS=1.515 NRD=0 NRS=46.14 M=1 R=4.93333
+ SA=75007.9 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1010 N_SUM_M1004_d N_A_992_347#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75008.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_27_378#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.263562 AS=0.295 PD=1.655 PS=2.59 NRD=17.73 NRS=3.2702 M=1 R=6.66667
+ SA=75000.2 SB=75007.1 A=0.15 P=2.3 MULT=1
MM1005 N_A_27_378#_M1005_d N_B_M1005_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.263562 PD=1.3 PS=1.655 NRD=1.9503 NRS=26.5753 M=1 R=6.66667
+ SA=75000.8 SB=75006.9 A=0.15 P=2.3 MULT=1
MM1012 N_A_336_347#_M1012_d N_CIN_M1012_g N_A_27_378#_M1005_d VPB PHIGHVT L=0.15
+ W=1 AD=0.295 AS=0.15 PD=1.59 PS=1.3 NRD=35.4403 NRS=1.9503 M=1 R=6.66667
+ SA=75001.2 SB=75006.4 A=0.15 P=2.3 MULT=1
MM1022 A_484_347# N_B_M1022_g N_A_336_347#_M1012_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.295 PD=1.27 PS=1.59 NRD=15.7403 NRS=25.5903 M=1 R=6.66667
+ SA=75002 SB=75005.7 A=0.15 P=2.3 MULT=1
MM1016 N_VPWR_M1016_d N_A_M1016_g A_484_347# VPB PHIGHVT L=0.15 W=1 AD=0.2125
+ AS=0.135 PD=1.425 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667 SA=75002.4
+ SB=75005.2 A=0.15 P=2.3 MULT=1
MM1006 N_A_683_347#_M1006_d N_CIN_M1006_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=1
+ AD=0.191062 AS=0.2125 PD=1.51 PS=1.425 NRD=2.9353 NRS=26.5753 M=1 R=6.66667
+ SA=75002.9 SB=75004.7 A=0.15 P=2.3 MULT=1
MM1023 N_VPWR_M1023_d N_B_M1023_g N_A_683_347#_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.233562 AS=0.191062 PD=1.595 PS=1.51 NRD=6.8753 NRS=11.8003 M=1 R=6.66667
+ SA=75003 SB=75004.3 A=0.15 P=2.3 MULT=1
MM1018 N_A_683_347#_M1018_d N_A_M1018_g N_VPWR_M1023_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.233562 PD=1.3 PS=1.595 NRD=1.9503 NRS=25.5903 M=1 R=6.66667
+ SA=75003.5 SB=75004.1 A=0.15 P=2.3 MULT=1
MM1030 N_A_992_347#_M1030_d N_A_336_347#_M1030_g N_A_683_347#_M1018_d VPB
+ PHIGHVT L=0.15 W=1 AD=0.18 AS=0.15 PD=1.36 PS=1.3 NRD=13.7703 NRS=1.9503 M=1
+ R=6.66667 SA=75004 SB=75003.6 A=0.15 P=2.3 MULT=1
MM1025 A_1094_347# N_CIN_M1025_g N_A_992_347#_M1030_d VPB PHIGHVT L=0.15 W=1
+ AD=0.20235 AS=0.18 PD=1.495 PS=1.36 NRD=29.0181 NRS=1.9503 M=1 R=6.66667
+ SA=75004.5 SB=75003.1 A=0.15 P=2.3 MULT=1
MM1026 A_1202_368# N_B_M1026_g A_1094_347# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.20235 PD=1.27 PS=1.495 NRD=15.7403 NRS=29.0181 M=1 R=6.66667 SA=75004.9
+ SB=75002.9 A=0.15 P=2.3 MULT=1
MM1020 N_VPWR_M1020_d N_A_M1020_g A_1202_368# VPB PHIGHVT L=0.15 W=1 AD=0.214811
+ AS=0.135 PD=1.45283 PS=1.27 NRD=26.5753 NRS=15.7403 M=1 R=6.66667 SA=75005.3
+ SB=75002.5 A=0.15 P=2.3 MULT=1
MM1009 N_COUT_M1009_d N_A_336_347#_M1009_g N_VPWR_M1020_d VPB PHIGHVT L=0.15
+ W=1.12 AD=0.2212 AS=0.240589 PD=1.515 PS=1.62717 NRD=9.6727 NRS=1.7533 M=1
+ R=7.46667 SA=75005.3 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1027 N_COUT_M1009_d N_A_336_347#_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.2212 AS=0.3024 PD=1.515 PS=1.66 NRD=10.5395 NRS=18.4589 M=1
+ R=7.46667 SA=75005.8 SB=75001.4 A=0.168 P=2.54 MULT=1
MM1014 N_SUM_M1014_d N_A_992_347#_M1014_g N_VPWR_M1027_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3024 PD=1.42 PS=1.66 NRD=1.7533 NRS=27.2451 M=1 R=7.46667
+ SA=75006.5 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1024 N_SUM_M1014_d N_A_992_347#_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.9 SB=75000.2 A=0.168 P=2.54 MULT=1
DX32_noxref VNB VPB NWDIODE A=18.2244 P=22.93
c_83 VNB 0 1.3983e-19 $X=0 $Y=0
c_1274 A_1094_347# 0 1.35287e-19 $X=5.47 $Y=1.735
*
.include "sky130_fd_sc_ls__fa_2.pxi.spice"
*
.ends
*
*
