* File: sky130_fd_sc_ls__sdfxtp_4.pxi.spice
* Created: Fri Aug 28 14:06:02 2020
* 
x_PM_SKY130_FD_SC_LS__SDFXTP_4%A_36_74# N_A_36_74#_M1036_s N_A_36_74#_M1024_s
+ N_A_36_74#_M1020_g N_A_36_74#_c_255_n N_A_36_74#_M1016_g N_A_36_74#_c_249_n
+ N_A_36_74#_c_257_n N_A_36_74#_c_250_n N_A_36_74#_c_258_n N_A_36_74#_c_259_n
+ N_A_36_74#_c_251_n N_A_36_74#_c_252_n N_A_36_74#_c_253_n N_A_36_74#_c_254_n
+ PM_SKY130_FD_SC_LS__SDFXTP_4%A_36_74#
x_PM_SKY130_FD_SC_LS__SDFXTP_4%SCE N_SCE_c_343_n N_SCE_c_351_n N_SCE_c_352_n
+ N_SCE_M1036_g N_SCE_c_353_n N_SCE_M1024_g N_SCE_c_354_n N_SCE_c_355_n
+ N_SCE_M1031_g N_SCE_c_345_n N_SCE_M1009_g N_SCE_c_356_n SCE N_SCE_c_346_n
+ N_SCE_c_347_n N_SCE_c_348_n N_SCE_c_349_n PM_SKY130_FD_SC_LS__SDFXTP_4%SCE
x_PM_SKY130_FD_SC_LS__SDFXTP_4%D N_D_M1021_g N_D_c_427_n N_D_c_428_n N_D_M1007_g
+ D N_D_c_425_n N_D_c_426_n PM_SKY130_FD_SC_LS__SDFXTP_4%D
x_PM_SKY130_FD_SC_LS__SDFXTP_4%SCD N_SCD_c_469_n N_SCD_c_470_n N_SCD_M1029_g
+ N_SCD_M1008_g SCD SCD N_SCD_c_468_n PM_SKY130_FD_SC_LS__SDFXTP_4%SCD
x_PM_SKY130_FD_SC_LS__SDFXTP_4%CLK N_CLK_c_514_n N_CLK_M1001_g N_CLK_c_515_n
+ N_CLK_M1023_g CLK PM_SKY130_FD_SC_LS__SDFXTP_4%CLK
x_PM_SKY130_FD_SC_LS__SDFXTP_4%A_828_74# N_A_828_74#_M1019_d N_A_828_74#_M1017_d
+ N_A_828_74#_c_575_n N_A_828_74#_M1000_g N_A_828_74#_c_555_n
+ N_A_828_74#_M1012_g N_A_828_74#_M1030_g N_A_828_74#_c_576_n
+ N_A_828_74#_c_577_n N_A_828_74#_M1005_g N_A_828_74#_c_557_n
+ N_A_828_74#_c_558_n N_A_828_74#_c_559_n N_A_828_74#_c_560_n
+ N_A_828_74#_c_561_n N_A_828_74#_c_562_n N_A_828_74#_c_563_n
+ N_A_828_74#_c_564_n N_A_828_74#_c_565_n N_A_828_74#_c_633_p
+ N_A_828_74#_c_566_n N_A_828_74#_c_567_n N_A_828_74#_c_568_n
+ N_A_828_74#_c_569_n N_A_828_74#_c_579_n N_A_828_74#_c_570_n
+ N_A_828_74#_c_660_p N_A_828_74#_c_571_n N_A_828_74#_c_572_n
+ N_A_828_74#_c_573_n N_A_828_74#_c_574_n PM_SKY130_FD_SC_LS__SDFXTP_4%A_828_74#
x_PM_SKY130_FD_SC_LS__SDFXTP_4%A_630_74# N_A_630_74#_M1001_d N_A_630_74#_M1023_d
+ N_A_630_74#_M1019_g N_A_630_74#_c_754_n N_A_630_74#_c_773_n
+ N_A_630_74#_M1017_g N_A_630_74#_c_755_n N_A_630_74#_M1025_g
+ N_A_630_74#_c_774_n N_A_630_74#_c_775_n N_A_630_74#_c_776_n
+ N_A_630_74#_M1011_g N_A_630_74#_c_757_n N_A_630_74#_M1022_g
+ N_A_630_74#_c_758_n N_A_630_74#_c_759_n N_A_630_74#_c_760_n
+ N_A_630_74#_M1018_g N_A_630_74#_c_762_n N_A_630_74#_c_763_n
+ N_A_630_74#_c_764_n N_A_630_74#_c_765_n N_A_630_74#_c_766_n
+ N_A_630_74#_c_767_n N_A_630_74#_c_781_n N_A_630_74#_c_768_n
+ N_A_630_74#_c_769_n N_A_630_74#_c_770_n N_A_630_74#_c_783_n
+ N_A_630_74#_c_784_n N_A_630_74#_c_878_p N_A_630_74#_c_785_n
+ N_A_630_74#_c_786_n N_A_630_74#_c_771_n N_A_630_74#_c_787_n
+ N_A_630_74#_c_772_n PM_SKY130_FD_SC_LS__SDFXTP_4%A_630_74#
x_PM_SKY130_FD_SC_LS__SDFXTP_4%A_1257_74# N_A_1257_74#_M1035_d
+ N_A_1257_74#_M1004_d N_A_1257_74#_M1034_g N_A_1257_74#_c_958_n
+ N_A_1257_74#_c_965_n N_A_1257_74#_M1026_g N_A_1257_74#_c_959_n
+ N_A_1257_74#_c_960_n N_A_1257_74#_c_961_n N_A_1257_74#_c_1004_n
+ N_A_1257_74#_c_984_n N_A_1257_74#_c_962_n N_A_1257_74#_c_963_n
+ PM_SKY130_FD_SC_LS__SDFXTP_4%A_1257_74#
x_PM_SKY130_FD_SC_LS__SDFXTP_4%A_1026_100# N_A_1026_100#_M1025_d
+ N_A_1026_100#_M1000_d N_A_1026_100#_c_1038_n N_A_1026_100#_M1004_g
+ N_A_1026_100#_M1035_g N_A_1026_100#_c_1034_n N_A_1026_100#_c_1035_n
+ N_A_1026_100#_c_1036_n N_A_1026_100#_c_1040_n N_A_1026_100#_c_1041_n
+ N_A_1026_100#_c_1037_n PM_SKY130_FD_SC_LS__SDFXTP_4%A_1026_100#
x_PM_SKY130_FD_SC_LS__SDFXTP_4%A_1814_48# N_A_1814_48#_M1027_s
+ N_A_1814_48#_M1010_d N_A_1814_48#_c_1114_n N_A_1814_48#_M1014_g
+ N_A_1814_48#_c_1115_n N_A_1814_48#_c_1116_n N_A_1814_48#_c_1129_n
+ N_A_1814_48#_M1037_g N_A_1814_48#_M1003_g N_A_1814_48#_c_1130_n
+ N_A_1814_48#_M1002_g N_A_1814_48#_c_1131_n N_A_1814_48#_M1006_g
+ N_A_1814_48#_M1013_g N_A_1814_48#_c_1132_n N_A_1814_48#_M1032_g
+ N_A_1814_48#_M1015_g N_A_1814_48#_c_1133_n N_A_1814_48#_M1033_g
+ N_A_1814_48#_M1028_g N_A_1814_48#_c_1121_n N_A_1814_48#_c_1122_n
+ N_A_1814_48#_c_1123_n N_A_1814_48#_c_1124_n N_A_1814_48#_c_1125_n
+ N_A_1814_48#_c_1126_n N_A_1814_48#_c_1134_n N_A_1814_48#_c_1135_n
+ N_A_1814_48#_c_1127_n PM_SKY130_FD_SC_LS__SDFXTP_4%A_1814_48#
x_PM_SKY130_FD_SC_LS__SDFXTP_4%A_1587_74# N_A_1587_74#_M1030_d
+ N_A_1587_74#_M1022_d N_A_1587_74#_c_1267_n N_A_1587_74#_M1010_g
+ N_A_1587_74#_c_1268_n N_A_1587_74#_c_1269_n N_A_1587_74#_c_1280_n
+ N_A_1587_74#_M1038_g N_A_1587_74#_M1027_g N_A_1587_74#_c_1271_n
+ N_A_1587_74#_c_1281_n N_A_1587_74#_c_1272_n N_A_1587_74#_c_1282_n
+ N_A_1587_74#_c_1283_n N_A_1587_74#_c_1273_n N_A_1587_74#_c_1274_n
+ N_A_1587_74#_c_1275_n N_A_1587_74#_c_1284_n N_A_1587_74#_c_1276_n
+ N_A_1587_74#_c_1277_n PM_SKY130_FD_SC_LS__SDFXTP_4%A_1587_74#
x_PM_SKY130_FD_SC_LS__SDFXTP_4%VPWR N_VPWR_M1024_d N_VPWR_M1029_d N_VPWR_M1017_s
+ N_VPWR_M1026_d N_VPWR_M1037_d N_VPWR_M1038_s N_VPWR_M1006_d N_VPWR_M1033_d
+ N_VPWR_c_1381_n N_VPWR_c_1382_n N_VPWR_c_1383_n N_VPWR_c_1384_n
+ N_VPWR_c_1385_n N_VPWR_c_1386_n N_VPWR_c_1387_n N_VPWR_c_1388_n
+ N_VPWR_c_1389_n N_VPWR_c_1390_n N_VPWR_c_1391_n VPWR N_VPWR_c_1392_n
+ N_VPWR_c_1393_n N_VPWR_c_1394_n N_VPWR_c_1395_n N_VPWR_c_1396_n
+ N_VPWR_c_1397_n N_VPWR_c_1398_n N_VPWR_c_1399_n N_VPWR_c_1400_n
+ N_VPWR_c_1401_n N_VPWR_c_1402_n N_VPWR_c_1380_n
+ PM_SKY130_FD_SC_LS__SDFXTP_4%VPWR
x_PM_SKY130_FD_SC_LS__SDFXTP_4%A_301_74# N_A_301_74#_M1021_d N_A_301_74#_M1025_s
+ N_A_301_74#_M1007_d N_A_301_74#_M1000_s N_A_301_74#_c_1540_n
+ N_A_301_74#_c_1541_n N_A_301_74#_c_1527_n N_A_301_74#_c_1528_n
+ N_A_301_74#_c_1529_n N_A_301_74#_c_1530_n N_A_301_74#_c_1535_n
+ N_A_301_74#_c_1531_n N_A_301_74#_c_1532_n N_A_301_74#_c_1533_n
+ N_A_301_74#_c_1537_n N_A_301_74#_c_1592_n N_A_301_74#_c_1538_n
+ N_A_301_74#_c_1644_n N_A_301_74#_c_1539_n
+ PM_SKY130_FD_SC_LS__SDFXTP_4%A_301_74#
x_PM_SKY130_FD_SC_LS__SDFXTP_4%Q N_Q_M1003_s N_Q_M1015_s N_Q_M1002_s N_Q_M1032_s
+ N_Q_c_1666_n N_Q_c_1660_n N_Q_c_1661_n N_Q_c_1662_n N_Q_c_1667_n N_Q_c_1668_n
+ N_Q_c_1669_n N_Q_c_1663_n N_Q_c_1670_n N_Q_c_1664_n Q
+ PM_SKY130_FD_SC_LS__SDFXTP_4%Q
x_PM_SKY130_FD_SC_LS__SDFXTP_4%VGND N_VGND_M1036_d N_VGND_M1008_d N_VGND_M1019_s
+ N_VGND_M1034_d N_VGND_M1014_d N_VGND_M1027_d N_VGND_M1013_d N_VGND_M1028_d
+ N_VGND_c_1733_n N_VGND_c_1734_n N_VGND_c_1735_n N_VGND_c_1736_n
+ N_VGND_c_1737_n N_VGND_c_1738_n N_VGND_c_1739_n N_VGND_c_1740_n
+ N_VGND_c_1741_n N_VGND_c_1742_n N_VGND_c_1743_n N_VGND_c_1744_n
+ N_VGND_c_1745_n N_VGND_c_1746_n N_VGND_c_1747_n VGND N_VGND_c_1748_n
+ N_VGND_c_1749_n N_VGND_c_1750_n N_VGND_c_1751_n N_VGND_c_1752_n
+ N_VGND_c_1753_n N_VGND_c_1754_n N_VGND_c_1755_n N_VGND_c_1756_n
+ PM_SKY130_FD_SC_LS__SDFXTP_4%VGND
cc_1 VNB N_A_36_74#_M1020_g 0.0490151f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_2 VNB N_A_36_74#_c_249_n 0.0188181f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.69
cc_3 VNB N_A_36_74#_c_250_n 0.0296807f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.525
cc_4 VNB N_A_36_74#_c_251_n 0.00213926f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_5 VNB N_A_36_74#_c_252_n 0.0173623f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_6 VNB N_A_36_74#_c_253_n 0.0216588f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=0.565
cc_7 VNB N_A_36_74#_c_254_n 0.00785153f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.825
cc_8 VNB N_SCE_c_343_n 0.0226362f $X=-0.19 $Y=-0.245 $X2=0.245 $Y2=2.32
cc_9 VNB N_SCE_M1036_g 0.0254968f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.525
cc_10 VNB N_SCE_c_345_n 0.0194158f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.525
cc_11 VNB N_SCE_c_346_n 0.0491505f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.567
cc_12 VNB N_SCE_c_347_n 0.0129414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_SCE_c_348_n 0.0394959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_SCE_c_349_n 0.0174105f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.69
cc_15 VNB N_D_M1021_g 0.0517509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_D_c_425_n 0.0161794f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=2.64
cc_17 VNB N_D_c_426_n 0.00377665f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.69
cc_18 VNB N_SCD_M1008_g 0.0593729f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_19 VNB SCD 0.00260181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_SCD_c_468_n 0.00891463f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.975
cc_21 VNB N_CLK_c_514_n 0.021694f $X=-0.19 $Y=-0.245 $X2=0.18 $Y2=0.37
cc_22 VNB N_CLK_c_515_n 0.0628877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB CLK 0.00720769f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.525
cc_24 VNB N_A_828_74#_c_555_n 0.0186508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_828_74#_M1030_g 0.0224561f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.975
cc_26 VNB N_A_828_74#_c_557_n 0.00968753f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.955
cc_27 VNB N_A_828_74#_c_558_n 0.0189124f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_28 VNB N_A_828_74#_c_559_n 0.00361019f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_29 VNB N_A_828_74#_c_560_n 0.0063862f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.567
cc_30 VNB N_A_828_74#_c_561_n 0.0175796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_828_74#_c_562_n 7.46964e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_828_74#_c_563_n 0.0031908f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.825
cc_33 VNB N_A_828_74#_c_564_n 0.0434008f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.825
cc_34 VNB N_A_828_74#_c_565_n 0.00948655f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.69
cc_35 VNB N_A_828_74#_c_566_n 0.00633546f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_36 VNB N_A_828_74#_c_567_n 0.00212722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_828_74#_c_568_n 0.00236499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_828_74#_c_569_n 0.00709406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_828_74#_c_570_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_828_74#_c_571_n 0.0326894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_828_74#_c_572_n 0.00870836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_828_74#_c_573_n 0.00308014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_828_74#_c_574_n 0.0229954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_630_74#_M1019_g 0.0265784f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_45 VNB N_A_630_74#_c_754_n 0.0220514f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=2.245
cc_46 VNB N_A_630_74#_c_755_n 0.0285836f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.785
cc_47 VNB N_A_630_74#_M1025_g 0.0460728f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=2.465
cc_48 VNB N_A_630_74#_c_757_n 0.00296197f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.567
cc_49 VNB N_A_630_74#_c_758_n 0.0289595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_630_74#_c_759_n 0.0301128f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.825
cc_51 VNB N_A_630_74#_c_760_n 0.0124319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_630_74#_M1018_g 0.0252697f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.69
cc_53 VNB N_A_630_74#_c_762_n 0.014598f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.825
cc_54 VNB N_A_630_74#_c_763_n 0.00855852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_630_74#_c_764_n 0.00858623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_630_74#_c_765_n 0.00806055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_630_74#_c_766_n 0.00801141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_630_74#_c_767_n 2.44598e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_630_74#_c_768_n 9.79198e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_630_74#_c_769_n 6.00443e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_630_74#_c_770_n 0.0386652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_630_74#_c_771_n 0.00328989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_630_74#_c_772_n 0.00268376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1257_74#_M1034_g 0.0277707f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_65 VNB N_A_1257_74#_c_958_n 0.0191132f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=2.64
cc_66 VNB N_A_1257_74#_c_959_n 0.0127069f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.785
cc_67 VNB N_A_1257_74#_c_960_n 0.00153902f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=2.04
cc_68 VNB N_A_1257_74#_c_961_n 0.00299466f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.955
cc_69 VNB N_A_1257_74#_c_962_n 0.00239652f $X=-0.19 $Y=-0.245 $X2=0.325
+ $Y2=0.565
cc_70 VNB N_A_1257_74#_c_963_n 0.0351021f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.825
cc_71 VNB N_A_1026_100#_M1035_g 0.0581128f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=2.64
cc_72 VNB N_A_1026_100#_c_1034_n 0.0177526f $X=-0.19 $Y=-0.245 $X2=0.17
+ $Y2=0.785
cc_73 VNB N_A_1026_100#_c_1035_n 0.011868f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=2.465
cc_74 VNB N_A_1026_100#_c_1036_n 0.00359387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1026_100#_c_1037_n 0.0147487f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.825
cc_76 VNB N_A_1814_48#_c_1114_n 0.0199283f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.525
cc_77 VNB N_A_1814_48#_c_1115_n 0.00716699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1814_48#_c_1116_n 0.0072661f $X=-0.19 $Y=-0.245 $X2=1.985
+ $Y2=2.245
cc_79 VNB N_A_1814_48#_M1003_g 0.0233037f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.465
cc_80 VNB N_A_1814_48#_M1013_g 0.0213942f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.567
cc_81 VNB N_A_1814_48#_M1015_g 0.0203016f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.825
cc_82 VNB N_A_1814_48#_M1028_g 0.0237682f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_83 VNB N_A_1814_48#_c_1121_n 0.0127275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1814_48#_c_1122_n 0.0122313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1814_48#_c_1123_n 0.00213324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1814_48#_c_1124_n 0.024907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1814_48#_c_1125_n 0.0123136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1814_48#_c_1126_n 0.0392798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1814_48#_c_1127_n 0.105142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1587_74#_c_1267_n 0.0159226f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.525
cc_91 VNB N_A_1587_74#_c_1268_n 0.0154092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1587_74#_c_1269_n 0.00194393f $X=-0.19 $Y=-0.245 $X2=1.985
+ $Y2=2.64
cc_93 VNB N_A_1587_74#_M1027_g 0.0338567f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.465
cc_94 VNB N_A_1587_74#_c_1271_n 0.00597846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1587_74#_c_1272_n 0.00443001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1587_74#_c_1273_n 0.0158525f $X=-0.19 $Y=-0.245 $X2=0.325
+ $Y2=0.565
cc_97 VNB N_A_1587_74#_c_1274_n 5.09778e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1587_74#_c_1275_n 0.00376591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1587_74#_c_1276_n 0.0020424f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=1.825
cc_100 VNB N_A_1587_74#_c_1277_n 0.0011566f $X=-0.19 $Y=-0.245 $X2=2.03
+ $Y2=1.635
cc_101 VNB N_VPWR_c_1380_n 0.521925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_301_74#_c_1527_n 0.00234674f $X=-0.19 $Y=-0.245 $X2=1.865
+ $Y2=2.04
cc_103 VNB N_A_301_74#_c_1528_n 0.0134907f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.04
cc_104 VNB N_A_301_74#_c_1529_n 0.00681672f $X=-0.19 $Y=-0.245 $X2=2.03
+ $Y2=1.955
cc_105 VNB N_A_301_74#_c_1530_n 0.0054408f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_106 VNB N_A_301_74#_c_1531_n 2.93026e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_301_74#_c_1532_n 0.00461118f $X=-0.19 $Y=-0.245 $X2=0.325
+ $Y2=0.567
cc_108 VNB N_A_301_74#_c_1533_n 0.0154088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_Q_c_1660_n 0.00201266f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.465
cc_110 VNB N_Q_c_1661_n 0.0025518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_Q_c_1662_n 0.00343767f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.04
cc_112 VNB N_Q_c_1663_n 0.00195975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_Q_c_1664_n 0.0114845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB Q 0.0254971f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_115 VNB N_VGND_c_1733_n 0.00641221f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.567
cc_116 VNB N_VGND_c_1734_n 0.00956899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1735_n 0.0098347f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.825
cc_118 VNB N_VGND_c_1736_n 0.0120465f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.69
cc_119 VNB N_VGND_c_1737_n 0.00973411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1738_n 0.00520205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1739_n 0.00267297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1740_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1741_n 0.022631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1742_n 0.046746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1743_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1744_n 0.0206041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1745_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1746_n 0.0620957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1747_n 0.00632182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1748_n 0.0629321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1749_n 0.0194685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1750_n 0.0188435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1751_n 0.0150174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1752_n 0.0261461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1753_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1754_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1755_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1756_n 0.681112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VPB N_A_36_74#_c_255_n 0.0168561f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.245
cc_140 VPB N_A_36_74#_c_249_n 0.0234124f $X=-0.19 $Y=1.66 $X2=0.965 $Y2=1.69
cc_141 VPB N_A_36_74#_c_257_n 0.0209674f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.975
cc_142 VPB N_A_36_74#_c_258_n 0.0408284f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=2.465
cc_143 VPB N_A_36_74#_c_259_n 0.0216748f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=2.04
cc_144 VPB N_A_36_74#_c_252_n 0.0218206f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_145 VPB N_A_36_74#_c_254_n 0.0207696f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=1.825
cc_146 VPB N_SCE_c_343_n 0.0258923f $X=-0.19 $Y=1.66 $X2=0.245 $Y2=2.32
cc_147 VPB N_SCE_c_351_n 0.0141272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_SCE_c_352_n 0.010921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_SCE_c_353_n 0.0201282f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.58
cc_150 VPB N_SCE_c_354_n 0.0224948f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.64
cc_151 VPB N_SCE_c_355_n 0.0154896f $X=-0.19 $Y=1.66 $X2=0.965 $Y2=1.69
cc_152 VPB N_SCE_c_356_n 0.00488727f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=2.465
cc_153 VPB N_D_c_427_n 0.0217105f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_D_c_428_n 0.0221933f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.525
cc_155 VPB N_D_c_425_n 0.0107067f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.64
cc_156 VPB N_D_c_426_n 0.00253078f $X=-0.19 $Y=1.66 $X2=0.965 $Y2=1.69
cc_157 VPB N_SCD_c_469_n 0.0124229f $X=-0.19 $Y=1.66 $X2=0.245 $Y2=2.32
cc_158 VPB N_SCD_c_470_n 0.0248549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB SCD 0.00304953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_SCD_c_468_n 0.0257778f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.975
cc_161 VPB N_CLK_c_515_n 0.0270292f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_828_74#_c_575_n 0.0185475f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.525
cc_163 VPB N_A_828_74#_c_576_n 0.0272614f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=2.125
cc_164 VPB N_A_828_74#_c_577_n 0.0230089f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=2.465
cc_165 VPB N_A_828_74#_c_560_n 0.0167142f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=0.567
cc_166 VPB N_A_828_74#_c_579_n 0.0540169f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_828_74#_c_573_n 0.00149822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_828_74#_c_574_n 0.00797126f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_630_74#_c_773_n 0.0214384f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.64
cc_170 VPB N_A_630_74#_c_774_n 0.0651691f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=2.04
cc_171 VPB N_A_630_74#_c_775_n 0.0205374f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_172 VPB N_A_630_74#_c_776_n 0.0431587f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_173 VPB N_A_630_74#_c_757_n 0.043006f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=0.567
cc_174 VPB N_A_630_74#_c_762_n 0.00806617f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=1.825
cc_175 VPB N_A_630_74#_c_763_n 0.0108427f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_630_74#_c_764_n 0.0281562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_630_74#_c_781_n 0.0113727f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_630_74#_c_769_n 0.0033331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_630_74#_c_783_n 0.00440291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_630_74#_c_784_n 0.0126187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_630_74#_c_785_n 0.00304474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_630_74#_c_786_n 0.012145f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_630_74#_c_787_n 0.00393484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_630_74#_c_772_n 0.00215264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_1257_74#_c_958_n 0.0395338f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.64
cc_186 VPB N_A_1257_74#_c_965_n 0.0234006f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.64
cc_187 VPB N_A_1257_74#_c_961_n 0.00549227f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.955
cc_188 VPB N_A_1026_100#_c_1038_n 0.0211162f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.525
cc_189 VPB N_A_1026_100#_c_1035_n 0.017023f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=2.465
cc_190 VPB N_A_1026_100#_c_1040_n 0.00544024f $X=-0.19 $Y=1.66 $X2=2.03
+ $Y2=1.635
cc_191 VPB N_A_1026_100#_c_1041_n 0.00856705f $X=-0.19 $Y=1.66 $X2=2.03
+ $Y2=1.635
cc_192 VPB N_A_1026_100#_c_1037_n 0.0414634f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.825
cc_193 VPB N_A_1814_48#_c_1116_n 0.0273109f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.245
cc_194 VPB N_A_1814_48#_c_1129_n 0.0213806f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.64
cc_195 VPB N_A_1814_48#_c_1130_n 0.0161879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_1814_48#_c_1131_n 0.0152283f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.955
cc_197 VPB N_A_1814_48#_c_1132_n 0.0147072f $X=-0.19 $Y=1.66 $X2=0.325 $Y2=0.567
cc_198 VPB N_A_1814_48#_c_1133_n 0.0173358f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.69
cc_199 VPB N_A_1814_48#_c_1134_n 0.00333712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_1814_48#_c_1135_n 0.00241715f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_1814_48#_c_1127_n 0.0270437f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_1587_74#_c_1267_n 0.0344f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.525
cc_203 VPB N_A_1587_74#_c_1269_n 0.00689445f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.64
cc_204 VPB N_A_1587_74#_c_1280_n 0.0212508f $X=-0.19 $Y=1.66 $X2=0.965 $Y2=1.69
cc_205 VPB N_A_1587_74#_c_1281_n 0.00227012f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.955
cc_206 VPB N_A_1587_74#_c_1282_n 0.0162864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_1587_74#_c_1283_n 0.00429246f $X=-0.19 $Y=1.66 $X2=0.325
+ $Y2=0.567
cc_208 VPB N_A_1587_74#_c_1284_n 0.00210678f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.825
cc_209 VPB N_A_1587_74#_c_1276_n 0.00414731f $X=-0.19 $Y=1.66 $X2=0.915
+ $Y2=1.825
cc_210 VPB N_A_1587_74#_c_1277_n 0.00130798f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_211 VPB N_VPWR_c_1381_n 0.00875225f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_212 VPB N_VPWR_c_1382_n 0.00810949f $X=-0.19 $Y=1.66 $X2=0.325 $Y2=0.567
cc_213 VPB N_VPWR_c_1383_n 0.021301f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1384_n 0.0215047f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.825
cc_215 VPB N_VPWR_c_1385_n 0.0112021f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.69
cc_216 VPB N_VPWR_c_1386_n 0.0209223f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_217 VPB N_VPWR_c_1387_n 0.00504372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1388_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1389_n 0.0393005f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1390_n 0.0215455f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1391_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1392_n 0.0457766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1393_n 0.0214801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1394_n 0.0604843f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1395_n 0.063807f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1396_n 0.0162902f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1397_n 0.0179897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1398_n 0.0252449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1399_n 0.00631504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1400_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1401_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1402_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1380_n 0.163242f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_301_74#_c_1530_n 0.00370565f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_235 VPB N_A_301_74#_c_1535_n 0.00931039f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_236 VPB N_A_301_74#_c_1531_n 0.00165322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_301_74#_c_1537_n 0.00744679f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_301_74#_c_1538_n 0.00519454f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.69
cc_239 VPB N_A_301_74#_c_1539_n 0.00688331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_Q_c_1666_n 0.00257348f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.975
cc_241 VPB N_Q_c_1667_n 0.00236302f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_242 VPB N_Q_c_1668_n 0.00183475f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_243 VPB N_Q_c_1669_n 0.00198541f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=0.567
cc_244 VPB N_Q_c_1670_n 0.00992123f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.69
cc_245 VPB Q 0.0076623f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_246 N_A_36_74#_M1020_g N_SCE_c_343_n 0.00365204f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_247 N_A_36_74#_c_249_n N_SCE_c_343_n 0.0181319f $X=0.965 $Y=1.69 $X2=0 $Y2=0
cc_248 N_A_36_74#_c_250_n N_SCE_c_343_n 0.0150312f $X=0.17 $Y=1.525 $X2=0 $Y2=0
cc_249 N_A_36_74#_c_254_n N_SCE_c_343_n 0.02872f $X=0.915 $Y=1.825 $X2=0 $Y2=0
cc_250 N_A_36_74#_c_258_n N_SCE_c_351_n 0.00743868f $X=0.39 $Y=2.465 $X2=0 $Y2=0
cc_251 N_A_36_74#_c_254_n N_SCE_c_351_n 0.00558688f $X=0.915 $Y=1.825 $X2=0
+ $Y2=0
cc_252 N_A_36_74#_c_258_n N_SCE_c_352_n 0.00791271f $X=0.39 $Y=2.465 $X2=0 $Y2=0
cc_253 N_A_36_74#_c_254_n N_SCE_c_352_n 0.00136027f $X=0.915 $Y=1.825 $X2=0
+ $Y2=0
cc_254 N_A_36_74#_M1020_g N_SCE_M1036_g 0.0165198f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_255 N_A_36_74#_c_250_n N_SCE_M1036_g 0.00555867f $X=0.17 $Y=1.525 $X2=0 $Y2=0
cc_256 N_A_36_74#_c_253_n N_SCE_M1036_g 0.00594445f $X=0.325 $Y=0.565 $X2=0
+ $Y2=0
cc_257 N_A_36_74#_c_258_n N_SCE_c_353_n 0.00970192f $X=0.39 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A_36_74#_c_259_n N_SCE_c_354_n 0.0121527f $X=1.865 $Y=2.04 $X2=0 $Y2=0
cc_259 N_A_36_74#_c_254_n N_SCE_c_354_n 0.00663735f $X=0.915 $Y=1.825 $X2=0
+ $Y2=0
cc_260 N_A_36_74#_c_258_n N_SCE_c_355_n 4.2278e-19 $X=0.39 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A_36_74#_c_249_n N_SCE_c_356_n 0.0290107f $X=0.965 $Y=1.69 $X2=0 $Y2=0
cc_262 N_A_36_74#_c_258_n N_SCE_c_356_n 0.0059435f $X=0.39 $Y=2.465 $X2=0 $Y2=0
cc_263 N_A_36_74#_c_254_n N_SCE_c_356_n 0.00954427f $X=0.915 $Y=1.825 $X2=0
+ $Y2=0
cc_264 N_A_36_74#_M1020_g N_SCE_c_346_n 0.0213665f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_265 N_A_36_74#_c_249_n N_SCE_c_346_n 0.00889754f $X=0.965 $Y=1.69 $X2=0 $Y2=0
cc_266 N_A_36_74#_c_250_n N_SCE_c_346_n 0.00782677f $X=0.17 $Y=1.525 $X2=0 $Y2=0
cc_267 N_A_36_74#_c_253_n N_SCE_c_346_n 0.00584522f $X=0.325 $Y=0.565 $X2=0
+ $Y2=0
cc_268 N_A_36_74#_c_254_n N_SCE_c_346_n 0.00761616f $X=0.915 $Y=1.825 $X2=0
+ $Y2=0
cc_269 N_A_36_74#_c_251_n N_SCE_c_347_n 0.0265176f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_270 N_A_36_74#_c_252_n N_SCE_c_347_n 0.00120449f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_271 N_A_36_74#_c_251_n N_SCE_c_348_n 3.72097e-19 $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_272 N_A_36_74#_c_252_n N_SCE_c_348_n 0.018258f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_273 N_A_36_74#_M1020_g N_SCE_c_349_n 0.020864f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_274 N_A_36_74#_c_249_n N_SCE_c_349_n 0.00540176f $X=0.965 $Y=1.69 $X2=0 $Y2=0
cc_275 N_A_36_74#_c_250_n N_SCE_c_349_n 0.0256551f $X=0.17 $Y=1.525 $X2=0 $Y2=0
cc_276 N_A_36_74#_c_259_n N_SCE_c_349_n 0.0111746f $X=1.865 $Y=2.04 $X2=0 $Y2=0
cc_277 N_A_36_74#_c_253_n N_SCE_c_349_n 0.00341751f $X=0.325 $Y=0.565 $X2=0
+ $Y2=0
cc_278 N_A_36_74#_c_254_n N_SCE_c_349_n 0.0306627f $X=0.915 $Y=1.825 $X2=0 $Y2=0
cc_279 N_A_36_74#_M1020_g N_D_M1021_g 0.065161f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_280 N_A_36_74#_c_249_n N_D_c_427_n 0.00308042f $X=0.965 $Y=1.69 $X2=0 $Y2=0
cc_281 N_A_36_74#_c_257_n N_D_c_427_n 0.00563966f $X=2.03 $Y=1.975 $X2=0 $Y2=0
cc_282 N_A_36_74#_c_259_n N_D_c_427_n 0.0176729f $X=1.865 $Y=2.04 $X2=0 $Y2=0
cc_283 N_A_36_74#_c_251_n N_D_c_427_n 0.00111327f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_284 N_A_36_74#_c_252_n N_D_c_427_n 0.0196508f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_285 N_A_36_74#_c_254_n N_D_c_427_n 0.00316536f $X=0.915 $Y=1.825 $X2=0 $Y2=0
cc_286 N_A_36_74#_c_255_n N_D_c_428_n 0.00953633f $X=1.985 $Y=2.245 $X2=0 $Y2=0
cc_287 N_A_36_74#_M1020_g N_D_c_425_n 0.0214207f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_288 N_A_36_74#_c_259_n N_D_c_425_n 0.00371768f $X=1.865 $Y=2.04 $X2=0 $Y2=0
cc_289 N_A_36_74#_c_251_n N_D_c_425_n 3.9661e-19 $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_290 N_A_36_74#_c_252_n N_D_c_425_n 0.0198258f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_291 N_A_36_74#_M1020_g N_D_c_426_n 0.00420444f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_292 N_A_36_74#_c_249_n N_D_c_426_n 0.00698958f $X=0.965 $Y=1.69 $X2=0 $Y2=0
cc_293 N_A_36_74#_c_259_n N_D_c_426_n 0.0430317f $X=1.865 $Y=2.04 $X2=0 $Y2=0
cc_294 N_A_36_74#_c_251_n N_D_c_426_n 0.0208514f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_295 N_A_36_74#_c_252_n N_D_c_426_n 0.00109252f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_296 N_A_36_74#_c_254_n N_D_c_426_n 0.0215506f $X=0.915 $Y=1.825 $X2=0 $Y2=0
cc_297 N_A_36_74#_c_257_n N_SCD_c_469_n 0.0178983f $X=2.03 $Y=1.975 $X2=0 $Y2=0
cc_298 N_A_36_74#_c_259_n N_SCD_c_469_n 6.06626e-19 $X=1.865 $Y=2.04 $X2=0 $Y2=0
cc_299 N_A_36_74#_c_255_n N_SCD_c_470_n 0.0259129f $X=1.985 $Y=2.245 $X2=0 $Y2=0
cc_300 N_A_36_74#_c_251_n N_SCD_M1008_g 5.61529e-19 $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_301 N_A_36_74#_c_252_n N_SCD_M1008_g 0.00579641f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_302 N_A_36_74#_c_259_n SCD 0.0111133f $X=1.865 $Y=2.04 $X2=0 $Y2=0
cc_303 N_A_36_74#_c_251_n SCD 0.0232698f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_304 N_A_36_74#_c_252_n SCD 0.00191524f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_305 N_A_36_74#_c_251_n N_SCD_c_468_n 0.00126093f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_306 N_A_36_74#_c_252_n N_SCD_c_468_n 0.0136147f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_307 N_A_36_74#_c_258_n N_VPWR_c_1381_n 0.0285143f $X=0.39 $Y=2.465 $X2=0
+ $Y2=0
cc_308 N_A_36_74#_c_254_n N_VPWR_c_1381_n 0.0271045f $X=0.915 $Y=1.825 $X2=0
+ $Y2=0
cc_309 N_A_36_74#_c_258_n N_VPWR_c_1390_n 0.0208407f $X=0.39 $Y=2.465 $X2=0
+ $Y2=0
cc_310 N_A_36_74#_c_255_n N_VPWR_c_1392_n 0.00445602f $X=1.985 $Y=2.245 $X2=0
+ $Y2=0
cc_311 N_A_36_74#_c_255_n N_VPWR_c_1397_n 0.00127463f $X=1.985 $Y=2.245 $X2=0
+ $Y2=0
cc_312 N_A_36_74#_c_255_n N_VPWR_c_1380_n 0.00438648f $X=1.985 $Y=2.245 $X2=0
+ $Y2=0
cc_313 N_A_36_74#_c_258_n N_VPWR_c_1380_n 0.0172173f $X=0.39 $Y=2.465 $X2=0
+ $Y2=0
cc_314 N_A_36_74#_M1020_g N_A_301_74#_c_1540_n 6.99132e-19 $X=1.04 $Y=0.58 $X2=0
+ $Y2=0
cc_315 N_A_36_74#_c_255_n N_A_301_74#_c_1541_n 0.009774f $X=1.985 $Y=2.245 $X2=0
+ $Y2=0
cc_316 N_A_36_74#_c_257_n N_A_301_74#_c_1541_n 6.60098e-19 $X=2.03 $Y=1.975
+ $X2=0 $Y2=0
cc_317 N_A_36_74#_c_259_n N_A_301_74#_c_1541_n 0.0138117f $X=1.865 $Y=2.04 $X2=0
+ $Y2=0
cc_318 N_A_36_74#_c_255_n N_A_301_74#_c_1538_n 0.0105369f $X=1.985 $Y=2.245
+ $X2=0 $Y2=0
cc_319 N_A_36_74#_c_257_n N_A_301_74#_c_1538_n 6.9574e-19 $X=2.03 $Y=1.975 $X2=0
+ $Y2=0
cc_320 N_A_36_74#_c_259_n N_A_301_74#_c_1538_n 0.0265031f $X=1.865 $Y=2.04 $X2=0
+ $Y2=0
cc_321 N_A_36_74#_M1020_g N_VGND_c_1733_n 0.0120744f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_322 N_A_36_74#_c_253_n N_VGND_c_1733_n 0.0176087f $X=0.325 $Y=0.565 $X2=0
+ $Y2=0
cc_323 N_A_36_74#_M1020_g N_VGND_c_1742_n 0.00383152f $X=1.04 $Y=0.58 $X2=0
+ $Y2=0
cc_324 N_A_36_74#_c_253_n N_VGND_c_1752_n 0.017355f $X=0.325 $Y=0.565 $X2=0
+ $Y2=0
cc_325 N_A_36_74#_M1020_g N_VGND_c_1756_n 0.0075725f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_326 N_A_36_74#_c_253_n N_VGND_c_1756_n 0.0146072f $X=0.325 $Y=0.565 $X2=0
+ $Y2=0
cc_327 N_SCE_c_345_n N_D_M1021_g 0.0124029f $X=2.185 $Y=0.9 $X2=0 $Y2=0
cc_328 N_SCE_c_347_n N_D_M1021_g 0.00479723f $X=2.03 $Y=1.065 $X2=0 $Y2=0
cc_329 N_SCE_c_348_n N_D_M1021_g 0.0104743f $X=2.185 $Y=1.065 $X2=0 $Y2=0
cc_330 N_SCE_c_349_n N_D_M1021_g 0.0217242f $X=1.565 $Y=1.047 $X2=0 $Y2=0
cc_331 N_SCE_c_354_n N_D_c_427_n 0.00963193f $X=1.04 $Y=2.17 $X2=0 $Y2=0
cc_332 N_SCE_c_355_n N_D_c_428_n 0.036954f $X=1.115 $Y=2.245 $X2=0 $Y2=0
cc_333 N_SCE_c_349_n N_D_c_425_n 0.00459108f $X=1.565 $Y=1.047 $X2=0 $Y2=0
cc_334 N_SCE_c_354_n N_D_c_426_n 4.96306e-19 $X=1.04 $Y=2.17 $X2=0 $Y2=0
cc_335 N_SCE_c_349_n N_D_c_426_n 0.0454102f $X=1.565 $Y=1.047 $X2=0 $Y2=0
cc_336 N_SCE_c_345_n N_SCD_M1008_g 0.051937f $X=2.185 $Y=0.9 $X2=0 $Y2=0
cc_337 N_SCE_c_347_n N_SCD_M1008_g 6.88372e-19 $X=2.03 $Y=1.065 $X2=0 $Y2=0
cc_338 N_SCE_c_353_n N_VPWR_c_1381_n 0.00688056f $X=0.615 $Y=2.245 $X2=0 $Y2=0
cc_339 N_SCE_c_354_n N_VPWR_c_1381_n 0.00393386f $X=1.04 $Y=2.17 $X2=0 $Y2=0
cc_340 N_SCE_c_355_n N_VPWR_c_1381_n 0.0157029f $X=1.115 $Y=2.245 $X2=0 $Y2=0
cc_341 N_SCE_c_353_n N_VPWR_c_1390_n 0.00445602f $X=0.615 $Y=2.245 $X2=0 $Y2=0
cc_342 N_SCE_c_355_n N_VPWR_c_1392_n 0.00413917f $X=1.115 $Y=2.245 $X2=0 $Y2=0
cc_343 N_SCE_c_353_n N_VPWR_c_1380_n 0.00861184f $X=0.615 $Y=2.245 $X2=0 $Y2=0
cc_344 N_SCE_c_355_n N_VPWR_c_1380_n 0.00817532f $X=1.115 $Y=2.245 $X2=0 $Y2=0
cc_345 N_SCE_c_345_n N_A_301_74#_c_1540_n 0.0166661f $X=2.185 $Y=0.9 $X2=0 $Y2=0
cc_346 N_SCE_c_347_n N_A_301_74#_c_1540_n 0.0476568f $X=2.03 $Y=1.065 $X2=0
+ $Y2=0
cc_347 N_SCE_c_348_n N_A_301_74#_c_1540_n 0.0012945f $X=2.185 $Y=1.065 $X2=0
+ $Y2=0
cc_348 N_SCE_c_349_n N_A_301_74#_c_1540_n 0.0027972f $X=1.565 $Y=1.047 $X2=0
+ $Y2=0
cc_349 N_SCE_c_345_n N_A_301_74#_c_1527_n 0.0060927f $X=2.185 $Y=0.9 $X2=0 $Y2=0
cc_350 N_SCE_c_347_n N_A_301_74#_c_1527_n 0.0293371f $X=2.03 $Y=1.065 $X2=0
+ $Y2=0
cc_351 N_SCE_c_347_n N_A_301_74#_c_1529_n 0.00951665f $X=2.03 $Y=1.065 $X2=0
+ $Y2=0
cc_352 N_SCE_c_348_n N_A_301_74#_c_1529_n 3.79717e-19 $X=2.185 $Y=1.065 $X2=0
+ $Y2=0
cc_353 N_SCE_c_355_n N_A_301_74#_c_1538_n 0.00193095f $X=1.115 $Y=2.245 $X2=0
+ $Y2=0
cc_354 N_SCE_M1036_g N_VGND_c_1733_n 0.00544316f $X=0.54 $Y=0.58 $X2=0 $Y2=0
cc_355 N_SCE_c_346_n N_VGND_c_1733_n 0.00215627f $X=0.54 $Y=1.12 $X2=0 $Y2=0
cc_356 N_SCE_c_349_n N_VGND_c_1733_n 0.0248315f $X=1.565 $Y=1.047 $X2=0 $Y2=0
cc_357 N_SCE_c_345_n N_VGND_c_1742_n 0.00296985f $X=2.185 $Y=0.9 $X2=0 $Y2=0
cc_358 N_SCE_M1036_g N_VGND_c_1752_n 0.00433162f $X=0.54 $Y=0.58 $X2=0 $Y2=0
cc_359 N_SCE_M1036_g N_VGND_c_1756_n 0.00820923f $X=0.54 $Y=0.58 $X2=0 $Y2=0
cc_360 N_SCE_c_345_n N_VGND_c_1756_n 0.00366123f $X=2.185 $Y=0.9 $X2=0 $Y2=0
cc_361 N_D_c_428_n N_VPWR_c_1381_n 0.00252392f $X=1.535 $Y=2.245 $X2=0 $Y2=0
cc_362 N_D_c_428_n N_VPWR_c_1392_n 0.00445602f $X=1.535 $Y=2.245 $X2=0 $Y2=0
cc_363 N_D_c_428_n N_VPWR_c_1380_n 0.00858241f $X=1.535 $Y=2.245 $X2=0 $Y2=0
cc_364 N_D_M1021_g N_A_301_74#_c_1540_n 0.00973833f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_365 N_D_c_428_n N_A_301_74#_c_1538_n 0.012472f $X=1.535 $Y=2.245 $X2=0 $Y2=0
cc_366 N_D_M1021_g N_VGND_c_1733_n 0.00218966f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_367 N_D_M1021_g N_VGND_c_1742_n 0.00434051f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_368 N_D_M1021_g N_VGND_c_1756_n 0.00820535f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_369 N_SCD_M1008_g N_CLK_c_514_n 0.0281939f $X=2.575 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_370 N_SCD_c_469_n N_CLK_c_515_n 0.00393479f $X=2.525 $Y=2.155 $X2=0 $Y2=0
cc_371 N_SCD_c_470_n N_CLK_c_515_n 0.0135342f $X=2.525 $Y=2.245 $X2=0 $Y2=0
cc_372 N_SCD_M1008_g N_CLK_c_515_n 0.00367775f $X=2.575 $Y=0.58 $X2=0 $Y2=0
cc_373 N_SCD_c_468_n N_CLK_c_515_n 0.00692543f $X=2.6 $Y=1.775 $X2=0 $Y2=0
cc_374 N_SCD_M1008_g N_A_630_74#_c_767_n 5.18837e-19 $X=2.575 $Y=0.58 $X2=0
+ $Y2=0
cc_375 N_SCD_c_470_n N_VPWR_c_1392_n 0.00415318f $X=2.525 $Y=2.245 $X2=0 $Y2=0
cc_376 N_SCD_c_470_n N_VPWR_c_1397_n 0.0145263f $X=2.525 $Y=2.245 $X2=0 $Y2=0
cc_377 N_SCD_c_470_n N_VPWR_c_1380_n 0.00399473f $X=2.525 $Y=2.245 $X2=0 $Y2=0
cc_378 N_SCD_M1008_g N_A_301_74#_c_1540_n 0.00571599f $X=2.575 $Y=0.58 $X2=0
+ $Y2=0
cc_379 N_SCD_c_470_n N_A_301_74#_c_1541_n 0.0136916f $X=2.525 $Y=2.245 $X2=0
+ $Y2=0
cc_380 SCD N_A_301_74#_c_1541_n 0.0178592f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_381 N_SCD_c_468_n N_A_301_74#_c_1541_n 5.60776e-19 $X=2.6 $Y=1.775 $X2=0
+ $Y2=0
cc_382 N_SCD_M1008_g N_A_301_74#_c_1527_n 0.0122054f $X=2.575 $Y=0.58 $X2=0
+ $Y2=0
cc_383 N_SCD_M1008_g N_A_301_74#_c_1528_n 0.0108788f $X=2.575 $Y=0.58 $X2=0
+ $Y2=0
cc_384 SCD N_A_301_74#_c_1528_n 0.0160708f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_385 N_SCD_c_468_n N_A_301_74#_c_1528_n 6.69081e-19 $X=2.6 $Y=1.775 $X2=0
+ $Y2=0
cc_386 N_SCD_M1008_g N_A_301_74#_c_1529_n 0.00345941f $X=2.575 $Y=0.58 $X2=0
+ $Y2=0
cc_387 SCD N_A_301_74#_c_1529_n 0.00786526f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_388 N_SCD_c_468_n N_A_301_74#_c_1529_n 4.24893e-19 $X=2.6 $Y=1.775 $X2=0
+ $Y2=0
cc_389 N_SCD_c_469_n N_A_301_74#_c_1530_n 0.00243312f $X=2.525 $Y=2.155 $X2=0
+ $Y2=0
cc_390 N_SCD_c_470_n N_A_301_74#_c_1530_n 0.00276684f $X=2.525 $Y=2.245 $X2=0
+ $Y2=0
cc_391 N_SCD_M1008_g N_A_301_74#_c_1530_n 0.0041215f $X=2.575 $Y=0.58 $X2=0
+ $Y2=0
cc_392 SCD N_A_301_74#_c_1530_n 0.0457958f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_393 N_SCD_c_468_n N_A_301_74#_c_1530_n 0.00259384f $X=2.6 $Y=1.775 $X2=0
+ $Y2=0
cc_394 N_SCD_c_470_n N_A_301_74#_c_1538_n 0.00190599f $X=2.525 $Y=2.245 $X2=0
+ $Y2=0
cc_395 N_SCD_M1008_g N_VGND_c_1734_n 0.00372502f $X=2.575 $Y=0.58 $X2=0 $Y2=0
cc_396 N_SCD_M1008_g N_VGND_c_1742_n 0.00423055f $X=2.575 $Y=0.58 $X2=0 $Y2=0
cc_397 N_SCD_M1008_g N_VGND_c_1756_n 0.00781486f $X=2.575 $Y=0.58 $X2=0 $Y2=0
cc_398 N_CLK_c_515_n N_A_630_74#_M1019_g 0.00234424f $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_399 CLK N_A_630_74#_M1019_g 4.4309e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_400 N_CLK_c_514_n N_A_630_74#_c_765_n 0.0062725f $X=3.075 $Y=1.22 $X2=0 $Y2=0
cc_401 N_CLK_c_515_n N_A_630_74#_c_766_n 9.4523e-19 $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_402 CLK N_A_630_74#_c_766_n 0.0183633f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_403 N_CLK_c_514_n N_A_630_74#_c_767_n 0.0042911f $X=3.075 $Y=1.22 $X2=0 $Y2=0
cc_404 N_CLK_c_515_n N_A_630_74#_c_767_n 0.00551046f $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_405 CLK N_A_630_74#_c_767_n 0.0157349f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_406 CLK N_A_630_74#_c_781_n 0.00174029f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_407 N_CLK_c_515_n N_A_630_74#_c_768_n 2.63894e-19 $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_408 N_CLK_c_515_n N_A_630_74#_c_769_n 0.00540383f $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_409 N_CLK_c_515_n N_A_630_74#_c_770_n 0.015756f $X=3.265 $Y=1.765 $X2=0 $Y2=0
cc_410 CLK N_A_630_74#_c_770_n 0.00161387f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_411 N_CLK_c_515_n N_A_630_74#_c_786_n 0.0112279f $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_412 CLK N_A_630_74#_c_786_n 0.0190511f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_413 N_CLK_c_515_n N_A_630_74#_c_771_n 2.21465e-19 $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_414 CLK N_A_630_74#_c_771_n 0.0296263f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_415 N_CLK_c_515_n N_VPWR_c_1393_n 0.00415318f $X=3.265 $Y=1.765 $X2=0 $Y2=0
cc_416 N_CLK_c_515_n N_VPWR_c_1397_n 0.0237454f $X=3.265 $Y=1.765 $X2=0 $Y2=0
cc_417 N_CLK_c_515_n N_VPWR_c_1398_n 0.00966956f $X=3.265 $Y=1.765 $X2=0 $Y2=0
cc_418 N_CLK_c_515_n N_VPWR_c_1380_n 0.00403443f $X=3.265 $Y=1.765 $X2=0 $Y2=0
cc_419 N_CLK_c_514_n N_A_301_74#_c_1527_n 0.00148975f $X=3.075 $Y=1.22 $X2=0
+ $Y2=0
cc_420 N_CLK_c_514_n N_A_301_74#_c_1528_n 0.00661351f $X=3.075 $Y=1.22 $X2=0
+ $Y2=0
cc_421 N_CLK_c_515_n N_A_301_74#_c_1528_n 0.00501474f $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_422 CLK N_A_301_74#_c_1528_n 0.0138976f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_423 N_CLK_c_515_n N_A_301_74#_c_1530_n 0.0206038f $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_424 CLK N_A_301_74#_c_1530_n 0.0151716f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_425 N_CLK_c_515_n N_A_301_74#_c_1535_n 0.0189575f $X=3.265 $Y=1.765 $X2=0
+ $Y2=0
cc_426 N_CLK_c_514_n N_VGND_c_1734_n 0.00539676f $X=3.075 $Y=1.22 $X2=0 $Y2=0
cc_427 N_CLK_c_514_n N_VGND_c_1735_n 0.0033335f $X=3.075 $Y=1.22 $X2=0 $Y2=0
cc_428 N_CLK_c_514_n N_VGND_c_1744_n 0.00434272f $X=3.075 $Y=1.22 $X2=0 $Y2=0
cc_429 N_CLK_c_514_n N_VGND_c_1756_n 0.00825771f $X=3.075 $Y=1.22 $X2=0 $Y2=0
cc_430 N_A_828_74#_c_557_n N_A_630_74#_M1019_g 0.0015901f $X=4.28 $Y=0.515 $X2=0
+ $Y2=0
cc_431 N_A_828_74#_c_559_n N_A_630_74#_M1019_g 0.00266901f $X=4.445 $Y=0.34
+ $X2=0 $Y2=0
cc_432 N_A_828_74#_c_557_n N_A_630_74#_c_754_n 0.00669668f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_433 N_A_828_74#_c_560_n N_A_630_74#_c_773_n 0.00217477f $X=5.18 $Y=2.04 $X2=0
+ $Y2=0
cc_434 N_A_828_74#_c_579_n N_A_630_74#_c_773_n 0.00521252f $X=5.24 $Y=2.205
+ $X2=0 $Y2=0
cc_435 N_A_828_74#_c_560_n N_A_630_74#_c_755_n 0.00192692f $X=5.18 $Y=2.04 $X2=0
+ $Y2=0
cc_436 N_A_828_74#_c_555_n N_A_630_74#_M1025_g 0.0134166f $X=5.735 $Y=1.03 $X2=0
+ $Y2=0
cc_437 N_A_828_74#_c_557_n N_A_630_74#_M1025_g 0.00323285f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_438 N_A_828_74#_c_558_n N_A_630_74#_M1025_g 0.00881128f $X=5.095 $Y=0.34
+ $X2=0 $Y2=0
cc_439 N_A_828_74#_c_560_n N_A_630_74#_M1025_g 0.0268052f $X=5.18 $Y=2.04 $X2=0
+ $Y2=0
cc_440 N_A_828_74#_c_570_n N_A_630_74#_M1025_g 0.00175971f $X=5.18 $Y=0.34 $X2=0
+ $Y2=0
cc_441 N_A_828_74#_c_560_n N_A_630_74#_c_774_n 0.00950878f $X=5.18 $Y=2.04 $X2=0
+ $Y2=0
cc_442 N_A_828_74#_c_563_n N_A_630_74#_c_774_n 3.40454e-19 $X=5.91 $Y=1.195
+ $X2=0 $Y2=0
cc_443 N_A_828_74#_c_564_n N_A_630_74#_c_774_n 0.0158989f $X=5.91 $Y=1.195 $X2=0
+ $Y2=0
cc_444 N_A_828_74#_c_579_n N_A_630_74#_c_774_n 0.00771818f $X=5.24 $Y=2.205
+ $X2=0 $Y2=0
cc_445 N_A_828_74#_c_579_n N_A_630_74#_c_775_n 0.00324993f $X=5.24 $Y=2.205
+ $X2=0 $Y2=0
cc_446 N_A_828_74#_c_575_n N_A_630_74#_c_776_n 0.0101337f $X=5.545 $Y=2.455
+ $X2=0 $Y2=0
cc_447 N_A_828_74#_c_579_n N_A_630_74#_c_776_n 0.0102782f $X=5.24 $Y=2.205 $X2=0
+ $Y2=0
cc_448 N_A_828_74#_c_576_n N_A_630_74#_c_757_n 0.0174736f $X=8.745 $Y=2.215
+ $X2=0 $Y2=0
cc_449 N_A_828_74#_c_577_n N_A_630_74#_c_757_n 0.00914653f $X=8.745 $Y=2.305
+ $X2=0 $Y2=0
cc_450 N_A_828_74#_c_569_n N_A_630_74#_c_757_n 0.00147398f $X=8.535 $Y=1.325
+ $X2=0 $Y2=0
cc_451 N_A_828_74#_c_569_n N_A_630_74#_c_758_n 0.0178299f $X=8.535 $Y=1.325
+ $X2=0 $Y2=0
cc_452 N_A_828_74#_c_573_n N_A_630_74#_c_758_n 0.00248381f $X=8.69 $Y=1.325
+ $X2=0 $Y2=0
cc_453 N_A_828_74#_c_574_n N_A_630_74#_c_758_n 0.0213283f $X=8.7 $Y=1.55 $X2=0
+ $Y2=0
cc_454 N_A_828_74#_c_569_n N_A_630_74#_c_759_n 0.00436518f $X=8.535 $Y=1.325
+ $X2=0 $Y2=0
cc_455 N_A_828_74#_c_573_n N_A_630_74#_c_759_n 0.00215779f $X=8.69 $Y=1.325
+ $X2=0 $Y2=0
cc_456 N_A_828_74#_c_574_n N_A_630_74#_c_759_n 0.0154685f $X=8.7 $Y=1.55 $X2=0
+ $Y2=0
cc_457 N_A_828_74#_M1030_g N_A_630_74#_c_760_n 0.00290209f $X=7.86 $Y=0.645
+ $X2=0 $Y2=0
cc_458 N_A_828_74#_c_568_n N_A_630_74#_c_760_n 4.78988e-19 $X=8.04 $Y=1.055
+ $X2=0 $Y2=0
cc_459 N_A_828_74#_c_571_n N_A_630_74#_c_760_n 0.0207468f $X=7.8 $Y=1.22 $X2=0
+ $Y2=0
cc_460 N_A_828_74#_c_572_n N_A_630_74#_c_760_n 0.00499098f $X=8.125 $Y=1.232
+ $X2=0 $Y2=0
cc_461 N_A_828_74#_c_566_n N_A_630_74#_M1018_g 0.00168666f $X=7.955 $Y=0.38
+ $X2=0 $Y2=0
cc_462 N_A_828_74#_c_568_n N_A_630_74#_M1018_g 7.82313e-19 $X=8.04 $Y=1.055
+ $X2=0 $Y2=0
cc_463 N_A_828_74#_c_560_n N_A_630_74#_c_762_n 3.90464e-19 $X=5.18 $Y=2.04 $X2=0
+ $Y2=0
cc_464 N_A_828_74#_c_560_n N_A_630_74#_c_763_n 0.0126158f $X=5.18 $Y=2.04 $X2=0
+ $Y2=0
cc_465 N_A_828_74#_c_579_n N_A_630_74#_c_763_n 0.0207943f $X=5.24 $Y=2.205 $X2=0
+ $Y2=0
cc_466 N_A_828_74#_c_571_n N_A_630_74#_c_764_n 0.0107644f $X=7.8 $Y=1.22 $X2=0
+ $Y2=0
cc_467 N_A_828_74#_c_572_n N_A_630_74#_c_764_n 0.00313968f $X=8.125 $Y=1.232
+ $X2=0 $Y2=0
cc_468 N_A_828_74#_c_557_n N_A_630_74#_c_771_n 0.0047909f $X=4.28 $Y=0.515 $X2=0
+ $Y2=0
cc_469 N_A_828_74#_c_576_n N_A_630_74#_c_772_n 0.00101223f $X=8.745 $Y=2.215
+ $X2=0 $Y2=0
cc_470 N_A_828_74#_c_571_n N_A_630_74#_c_772_n 2.34783e-19 $X=7.8 $Y=1.22 $X2=0
+ $Y2=0
cc_471 N_A_828_74#_c_572_n N_A_630_74#_c_772_n 0.0226074f $X=8.125 $Y=1.232
+ $X2=0 $Y2=0
cc_472 N_A_828_74#_c_573_n N_A_630_74#_c_772_n 0.00314277f $X=8.69 $Y=1.325
+ $X2=0 $Y2=0
cc_473 N_A_828_74#_c_574_n N_A_630_74#_c_772_n 2.24348e-19 $X=8.7 $Y=1.55 $X2=0
+ $Y2=0
cc_474 N_A_828_74#_c_566_n N_A_1257_74#_M1035_d 0.00364436f $X=7.955 $Y=0.38
+ $X2=-0.19 $Y2=-0.245
cc_475 N_A_828_74#_c_555_n N_A_1257_74#_M1034_g 0.0131205f $X=5.735 $Y=1.03
+ $X2=0 $Y2=0
cc_476 N_A_828_74#_c_561_n N_A_1257_74#_M1034_g 5.55205e-19 $X=5.775 $Y=0.34
+ $X2=0 $Y2=0
cc_477 N_A_828_74#_c_562_n N_A_1257_74#_M1034_g 0.0045554f $X=5.86 $Y=0.77 $X2=0
+ $Y2=0
cc_478 N_A_828_74#_c_563_n N_A_1257_74#_M1034_g 0.00354212f $X=5.91 $Y=1.195
+ $X2=0 $Y2=0
cc_479 N_A_828_74#_c_564_n N_A_1257_74#_M1034_g 0.0207835f $X=5.91 $Y=1.195
+ $X2=0 $Y2=0
cc_480 N_A_828_74#_c_565_n N_A_1257_74#_M1034_g 0.0146054f $X=6.99 $Y=0.855
+ $X2=0 $Y2=0
cc_481 N_A_828_74#_c_633_p N_A_1257_74#_M1034_g 0.00402963f $X=7.075 $Y=0.77
+ $X2=0 $Y2=0
cc_482 N_A_828_74#_c_563_n N_A_1257_74#_c_959_n 0.0160452f $X=5.91 $Y=1.195
+ $X2=0 $Y2=0
cc_483 N_A_828_74#_c_564_n N_A_1257_74#_c_959_n 8.89984e-19 $X=5.91 $Y=1.195
+ $X2=0 $Y2=0
cc_484 N_A_828_74#_c_565_n N_A_1257_74#_c_959_n 0.0681547f $X=6.99 $Y=0.855
+ $X2=0 $Y2=0
cc_485 N_A_828_74#_c_566_n N_A_1257_74#_c_959_n 0.00366775f $X=7.955 $Y=0.38
+ $X2=0 $Y2=0
cc_486 N_A_828_74#_M1030_g N_A_1257_74#_c_960_n 0.00138161f $X=7.86 $Y=0.645
+ $X2=0 $Y2=0
cc_487 N_A_828_74#_c_565_n N_A_1257_74#_c_960_n 0.00275859f $X=6.99 $Y=0.855
+ $X2=0 $Y2=0
cc_488 N_A_828_74#_c_568_n N_A_1257_74#_c_960_n 0.0057135f $X=8.04 $Y=1.055
+ $X2=0 $Y2=0
cc_489 N_A_828_74#_c_571_n N_A_1257_74#_c_960_n 3.77672e-19 $X=7.8 $Y=1.22 $X2=0
+ $Y2=0
cc_490 N_A_828_74#_c_572_n N_A_1257_74#_c_960_n 0.00414256f $X=8.125 $Y=1.232
+ $X2=0 $Y2=0
cc_491 N_A_828_74#_M1030_g N_A_1257_74#_c_984_n 0.00265713f $X=7.86 $Y=0.645
+ $X2=0 $Y2=0
cc_492 N_A_828_74#_c_566_n N_A_1257_74#_c_984_n 0.0240267f $X=7.955 $Y=0.38
+ $X2=0 $Y2=0
cc_493 N_A_828_74#_c_571_n N_A_1257_74#_c_984_n 0.00383634f $X=7.8 $Y=1.22 $X2=0
+ $Y2=0
cc_494 N_A_828_74#_c_572_n N_A_1257_74#_c_984_n 0.0065951f $X=8.125 $Y=1.232
+ $X2=0 $Y2=0
cc_495 N_A_828_74#_c_571_n N_A_1257_74#_c_962_n 0.00207447f $X=7.8 $Y=1.22 $X2=0
+ $Y2=0
cc_496 N_A_828_74#_c_572_n N_A_1257_74#_c_962_n 0.0264386f $X=8.125 $Y=1.232
+ $X2=0 $Y2=0
cc_497 N_A_828_74#_c_565_n N_A_1257_74#_c_963_n 0.00496909f $X=6.99 $Y=0.855
+ $X2=0 $Y2=0
cc_498 N_A_828_74#_c_560_n N_A_1026_100#_M1025_d 0.0042575f $X=5.18 $Y=2.04
+ $X2=-0.19 $Y2=-0.245
cc_499 N_A_828_74#_M1030_g N_A_1026_100#_M1035_g 0.0203971f $X=7.86 $Y=0.645
+ $X2=0 $Y2=0
cc_500 N_A_828_74#_c_565_n N_A_1026_100#_M1035_g 0.00337097f $X=6.99 $Y=0.855
+ $X2=0 $Y2=0
cc_501 N_A_828_74#_c_566_n N_A_1026_100#_M1035_g 0.0131439f $X=7.955 $Y=0.38
+ $X2=0 $Y2=0
cc_502 N_A_828_74#_c_571_n N_A_1026_100#_M1035_g 0.0140546f $X=7.8 $Y=1.22 $X2=0
+ $Y2=0
cc_503 N_A_828_74#_c_572_n N_A_1026_100#_M1035_g 4.49059e-19 $X=8.125 $Y=1.232
+ $X2=0 $Y2=0
cc_504 N_A_828_74#_c_555_n N_A_1026_100#_c_1034_n 0.00498983f $X=5.735 $Y=1.03
+ $X2=0 $Y2=0
cc_505 N_A_828_74#_c_560_n N_A_1026_100#_c_1034_n 0.0755586f $X=5.18 $Y=2.04
+ $X2=0 $Y2=0
cc_506 N_A_828_74#_c_561_n N_A_1026_100#_c_1034_n 0.012971f $X=5.775 $Y=0.34
+ $X2=0 $Y2=0
cc_507 N_A_828_74#_c_563_n N_A_1026_100#_c_1034_n 0.0312592f $X=5.91 $Y=1.195
+ $X2=0 $Y2=0
cc_508 N_A_828_74#_c_660_p N_A_1026_100#_c_1034_n 0.00787896f $X=5.925 $Y=0.855
+ $X2=0 $Y2=0
cc_509 N_A_828_74#_c_563_n N_A_1026_100#_c_1035_n 0.0177193f $X=5.91 $Y=1.195
+ $X2=0 $Y2=0
cc_510 N_A_828_74#_c_564_n N_A_1026_100#_c_1035_n 0.00103095f $X=5.91 $Y=1.195
+ $X2=0 $Y2=0
cc_511 N_A_828_74#_c_565_n N_A_1026_100#_c_1035_n 0.00630202f $X=6.99 $Y=0.855
+ $X2=0 $Y2=0
cc_512 N_A_828_74#_c_560_n N_A_1026_100#_c_1036_n 0.0133687f $X=5.18 $Y=2.04
+ $X2=0 $Y2=0
cc_513 N_A_828_74#_c_564_n N_A_1026_100#_c_1036_n 0.00236559f $X=5.91 $Y=1.195
+ $X2=0 $Y2=0
cc_514 N_A_828_74#_c_579_n N_A_1026_100#_c_1036_n 9.11699e-19 $X=5.24 $Y=2.205
+ $X2=0 $Y2=0
cc_515 N_A_828_74#_c_575_n N_A_1026_100#_c_1040_n 0.00783432f $X=5.545 $Y=2.455
+ $X2=0 $Y2=0
cc_516 N_A_828_74#_c_575_n N_A_1026_100#_c_1041_n 0.00260822f $X=5.545 $Y=2.455
+ $X2=0 $Y2=0
cc_517 N_A_828_74#_c_560_n N_A_1026_100#_c_1041_n 0.0376527f $X=5.18 $Y=2.04
+ $X2=0 $Y2=0
cc_518 N_A_828_74#_c_579_n N_A_1026_100#_c_1041_n 0.00994071f $X=5.24 $Y=2.205
+ $X2=0 $Y2=0
cc_519 N_A_828_74#_c_573_n N_A_1814_48#_c_1115_n 3.57139e-19 $X=8.69 $Y=1.325
+ $X2=0 $Y2=0
cc_520 N_A_828_74#_c_574_n N_A_1814_48#_c_1115_n 0.0204649f $X=8.7 $Y=1.55 $X2=0
+ $Y2=0
cc_521 N_A_828_74#_c_576_n N_A_1814_48#_c_1116_n 0.0155183f $X=8.745 $Y=2.215
+ $X2=0 $Y2=0
cc_522 N_A_828_74#_c_577_n N_A_1814_48#_c_1129_n 0.043208f $X=8.745 $Y=2.305
+ $X2=0 $Y2=0
cc_523 N_A_828_74#_c_573_n N_A_1814_48#_c_1122_n 8.55777e-19 $X=8.69 $Y=1.325
+ $X2=0 $Y2=0
cc_524 N_A_828_74#_c_566_n N_A_1587_74#_M1030_d 0.00100458f $X=7.955 $Y=0.38
+ $X2=-0.19 $Y2=-0.245
cc_525 N_A_828_74#_c_568_n N_A_1587_74#_M1030_d 0.00611407f $X=8.04 $Y=1.055
+ $X2=-0.19 $Y2=-0.245
cc_526 N_A_828_74#_c_576_n N_A_1587_74#_c_1281_n 0.00325391f $X=8.745 $Y=2.215
+ $X2=0 $Y2=0
cc_527 N_A_828_74#_c_577_n N_A_1587_74#_c_1281_n 0.00839216f $X=8.745 $Y=2.305
+ $X2=0 $Y2=0
cc_528 N_A_828_74#_M1030_g N_A_1587_74#_c_1272_n 0.00133546f $X=7.86 $Y=0.645
+ $X2=0 $Y2=0
cc_529 N_A_828_74#_c_566_n N_A_1587_74#_c_1272_n 0.0098597f $X=7.955 $Y=0.38
+ $X2=0 $Y2=0
cc_530 N_A_828_74#_c_568_n N_A_1587_74#_c_1272_n 0.033167f $X=8.04 $Y=1.055
+ $X2=0 $Y2=0
cc_531 N_A_828_74#_c_576_n N_A_1587_74#_c_1282_n 0.0181702f $X=8.745 $Y=2.215
+ $X2=0 $Y2=0
cc_532 N_A_828_74#_c_573_n N_A_1587_74#_c_1282_n 0.0115014f $X=8.69 $Y=1.325
+ $X2=0 $Y2=0
cc_533 N_A_828_74#_c_574_n N_A_1587_74#_c_1282_n 0.00107876f $X=8.7 $Y=1.55
+ $X2=0 $Y2=0
cc_534 N_A_828_74#_c_569_n N_A_1587_74#_c_1283_n 0.00885113f $X=8.535 $Y=1.325
+ $X2=0 $Y2=0
cc_535 N_A_828_74#_c_573_n N_A_1587_74#_c_1283_n 0.0035906f $X=8.69 $Y=1.325
+ $X2=0 $Y2=0
cc_536 N_A_828_74#_c_574_n N_A_1587_74#_c_1283_n 4.71321e-19 $X=8.7 $Y=1.55
+ $X2=0 $Y2=0
cc_537 N_A_828_74#_c_573_n N_A_1587_74#_c_1273_n 0.0171164f $X=8.69 $Y=1.325
+ $X2=0 $Y2=0
cc_538 N_A_828_74#_c_574_n N_A_1587_74#_c_1273_n 9.20427e-19 $X=8.7 $Y=1.55
+ $X2=0 $Y2=0
cc_539 N_A_828_74#_c_568_n N_A_1587_74#_c_1274_n 0.0127557f $X=8.04 $Y=1.055
+ $X2=0 $Y2=0
cc_540 N_A_828_74#_c_569_n N_A_1587_74#_c_1274_n 0.0191115f $X=8.535 $Y=1.325
+ $X2=0 $Y2=0
cc_541 N_A_828_74#_c_572_n N_A_1587_74#_c_1274_n 0.00120956f $X=8.125 $Y=1.232
+ $X2=0 $Y2=0
cc_542 N_A_828_74#_c_573_n N_A_1587_74#_c_1274_n 0.00774767f $X=8.69 $Y=1.325
+ $X2=0 $Y2=0
cc_543 N_A_828_74#_c_573_n N_A_1587_74#_c_1275_n 0.0177584f $X=8.69 $Y=1.325
+ $X2=0 $Y2=0
cc_544 N_A_828_74#_c_574_n N_A_1587_74#_c_1275_n 4.64187e-19 $X=8.7 $Y=1.55
+ $X2=0 $Y2=0
cc_545 N_A_828_74#_c_576_n N_A_1587_74#_c_1284_n 0.00439306f $X=8.745 $Y=2.215
+ $X2=0 $Y2=0
cc_546 N_A_828_74#_c_576_n N_A_1587_74#_c_1277_n 0.00228435f $X=8.745 $Y=2.215
+ $X2=0 $Y2=0
cc_547 N_A_828_74#_c_573_n N_A_1587_74#_c_1277_n 0.020573f $X=8.69 $Y=1.325
+ $X2=0 $Y2=0
cc_548 N_A_828_74#_c_574_n N_A_1587_74#_c_1277_n 0.00156371f $X=8.7 $Y=1.55
+ $X2=0 $Y2=0
cc_549 N_A_828_74#_c_577_n N_VPWR_c_1383_n 0.00190266f $X=8.745 $Y=2.305 $X2=0
+ $Y2=0
cc_550 N_A_828_74#_c_575_n N_VPWR_c_1394_n 0.00522247f $X=5.545 $Y=2.455 $X2=0
+ $Y2=0
cc_551 N_A_828_74#_c_577_n N_VPWR_c_1395_n 0.00469064f $X=8.745 $Y=2.305 $X2=0
+ $Y2=0
cc_552 N_A_828_74#_c_575_n N_VPWR_c_1380_n 0.00542671f $X=5.545 $Y=2.455 $X2=0
+ $Y2=0
cc_553 N_A_828_74#_c_577_n N_VPWR_c_1380_n 0.0049649f $X=8.745 $Y=2.305 $X2=0
+ $Y2=0
cc_554 N_A_828_74#_c_579_n N_VPWR_c_1380_n 3.17865e-19 $X=5.24 $Y=2.205 $X2=0
+ $Y2=0
cc_555 N_A_828_74#_c_560_n N_A_301_74#_c_1531_n 0.0383113f $X=5.18 $Y=2.04 $X2=0
+ $Y2=0
cc_556 N_A_828_74#_c_579_n N_A_301_74#_c_1531_n 2.7287e-19 $X=5.24 $Y=2.205
+ $X2=0 $Y2=0
cc_557 N_A_828_74#_c_557_n N_A_301_74#_c_1532_n 0.00515156f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_558 N_A_828_74#_c_560_n N_A_301_74#_c_1532_n 0.0329467f $X=5.18 $Y=2.04 $X2=0
+ $Y2=0
cc_559 N_A_828_74#_c_557_n N_A_301_74#_c_1533_n 0.0345841f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_560 N_A_828_74#_c_558_n N_A_301_74#_c_1533_n 0.0191962f $X=5.095 $Y=0.34
+ $X2=0 $Y2=0
cc_561 N_A_828_74#_c_560_n N_A_301_74#_c_1533_n 0.0522592f $X=5.18 $Y=2.04 $X2=0
+ $Y2=0
cc_562 N_A_828_74#_M1017_d N_A_301_74#_c_1537_n 0.00361533f $X=4.61 $Y=1.84
+ $X2=0 $Y2=0
cc_563 N_A_828_74#_c_560_n N_A_301_74#_c_1537_n 0.0195838f $X=5.18 $Y=2.04 $X2=0
+ $Y2=0
cc_564 N_A_828_74#_c_579_n N_A_301_74#_c_1537_n 5.63958e-19 $X=5.24 $Y=2.205
+ $X2=0 $Y2=0
cc_565 N_A_828_74#_M1017_d N_A_301_74#_c_1592_n 0.00795981f $X=4.61 $Y=1.84
+ $X2=0 $Y2=0
cc_566 N_A_828_74#_c_575_n N_A_301_74#_c_1592_n 0.00210767f $X=5.545 $Y=2.455
+ $X2=0 $Y2=0
cc_567 N_A_828_74#_c_560_n N_A_301_74#_c_1592_n 0.0114774f $X=5.18 $Y=2.04 $X2=0
+ $Y2=0
cc_568 N_A_828_74#_c_579_n N_A_301_74#_c_1592_n 0.00167232f $X=5.24 $Y=2.205
+ $X2=0 $Y2=0
cc_569 N_A_828_74#_c_575_n N_A_301_74#_c_1539_n 0.00203632f $X=5.545 $Y=2.455
+ $X2=0 $Y2=0
cc_570 N_A_828_74#_c_560_n N_A_301_74#_c_1539_n 0.020359f $X=5.18 $Y=2.04 $X2=0
+ $Y2=0
cc_571 N_A_828_74#_c_579_n N_A_301_74#_c_1539_n 0.00187948f $X=5.24 $Y=2.205
+ $X2=0 $Y2=0
cc_572 N_A_828_74#_c_565_n N_VGND_M1034_d 0.0110146f $X=6.99 $Y=0.855 $X2=0
+ $Y2=0
cc_573 N_A_828_74#_c_633_p N_VGND_M1034_d 0.00544097f $X=7.075 $Y=0.77 $X2=0
+ $Y2=0
cc_574 N_A_828_74#_c_567_n N_VGND_M1034_d 0.00113603f $X=7.16 $Y=0.38 $X2=0
+ $Y2=0
cc_575 N_A_828_74#_c_559_n N_VGND_c_1735_n 0.0112234f $X=4.445 $Y=0.34 $X2=0
+ $Y2=0
cc_576 N_A_828_74#_c_561_n N_VGND_c_1736_n 0.0066699f $X=5.775 $Y=0.34 $X2=0
+ $Y2=0
cc_577 N_A_828_74#_c_562_n N_VGND_c_1736_n 0.00411865f $X=5.86 $Y=0.77 $X2=0
+ $Y2=0
cc_578 N_A_828_74#_c_565_n N_VGND_c_1736_n 0.0258618f $X=6.99 $Y=0.855 $X2=0
+ $Y2=0
cc_579 N_A_828_74#_c_633_p N_VGND_c_1736_n 0.0102806f $X=7.075 $Y=0.77 $X2=0
+ $Y2=0
cc_580 N_A_828_74#_c_567_n N_VGND_c_1736_n 0.014725f $X=7.16 $Y=0.38 $X2=0 $Y2=0
cc_581 N_A_828_74#_c_555_n N_VGND_c_1746_n 7.26171e-19 $X=5.735 $Y=1.03 $X2=0
+ $Y2=0
cc_582 N_A_828_74#_c_558_n N_VGND_c_1746_n 0.0418136f $X=5.095 $Y=0.34 $X2=0
+ $Y2=0
cc_583 N_A_828_74#_c_559_n N_VGND_c_1746_n 0.0179217f $X=4.445 $Y=0.34 $X2=0
+ $Y2=0
cc_584 N_A_828_74#_c_561_n N_VGND_c_1746_n 0.0449818f $X=5.775 $Y=0.34 $X2=0
+ $Y2=0
cc_585 N_A_828_74#_c_570_n N_VGND_c_1746_n 0.0121867f $X=5.18 $Y=0.34 $X2=0
+ $Y2=0
cc_586 N_A_828_74#_M1030_g N_VGND_c_1748_n 0.00284028f $X=7.86 $Y=0.645 $X2=0
+ $Y2=0
cc_587 N_A_828_74#_c_566_n N_VGND_c_1748_n 0.0498254f $X=7.955 $Y=0.38 $X2=0
+ $Y2=0
cc_588 N_A_828_74#_c_567_n N_VGND_c_1748_n 0.00968103f $X=7.16 $Y=0.38 $X2=0
+ $Y2=0
cc_589 N_A_828_74#_M1030_g N_VGND_c_1756_n 0.00361049f $X=7.86 $Y=0.645 $X2=0
+ $Y2=0
cc_590 N_A_828_74#_c_558_n N_VGND_c_1756_n 0.0244305f $X=5.095 $Y=0.34 $X2=0
+ $Y2=0
cc_591 N_A_828_74#_c_559_n N_VGND_c_1756_n 0.00971942f $X=4.445 $Y=0.34 $X2=0
+ $Y2=0
cc_592 N_A_828_74#_c_561_n N_VGND_c_1756_n 0.025776f $X=5.775 $Y=0.34 $X2=0
+ $Y2=0
cc_593 N_A_828_74#_c_565_n N_VGND_c_1756_n 0.0222018f $X=6.99 $Y=0.855 $X2=0
+ $Y2=0
cc_594 N_A_828_74#_c_566_n N_VGND_c_1756_n 0.0342339f $X=7.955 $Y=0.38 $X2=0
+ $Y2=0
cc_595 N_A_828_74#_c_567_n N_VGND_c_1756_n 0.00646784f $X=7.16 $Y=0.38 $X2=0
+ $Y2=0
cc_596 N_A_828_74#_c_570_n N_VGND_c_1756_n 0.00660921f $X=5.18 $Y=0.34 $X2=0
+ $Y2=0
cc_597 N_A_828_74#_c_660_p N_VGND_c_1756_n 0.0053779f $X=5.925 $Y=0.855 $X2=0
+ $Y2=0
cc_598 N_A_828_74#_c_562_n A_1162_100# 0.00372609f $X=5.86 $Y=0.77 $X2=-0.19
+ $Y2=-0.245
cc_599 N_A_828_74#_c_565_n A_1162_100# 0.00299768f $X=6.99 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_600 N_A_828_74#_c_660_p A_1162_100# 0.00320575f $X=5.925 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_601 N_A_630_74#_c_784_n N_A_1257_74#_M1004_d 0.0279005f $X=7.93 $Y=2.6 $X2=0
+ $Y2=0
cc_602 N_A_630_74#_c_785_n N_A_1257_74#_M1004_d 0.0122344f $X=8.015 $Y=2.515
+ $X2=0 $Y2=0
cc_603 N_A_630_74#_c_774_n N_A_1257_74#_c_958_n 0.0380891f $X=5.905 $Y=1.755
+ $X2=0 $Y2=0
cc_604 N_A_630_74#_c_776_n N_A_1257_74#_c_958_n 0.00440286f $X=5.995 $Y=2.455
+ $X2=0 $Y2=0
cc_605 N_A_630_74#_c_783_n N_A_1257_74#_c_958_n 0.00379018f $X=6.19 $Y=2.515
+ $X2=0 $Y2=0
cc_606 N_A_630_74#_c_787_n N_A_1257_74#_c_958_n 0.00765601f $X=6.19 $Y=2.115
+ $X2=0 $Y2=0
cc_607 N_A_630_74#_c_776_n N_A_1257_74#_c_965_n 0.0179533f $X=5.995 $Y=2.455
+ $X2=0 $Y2=0
cc_608 N_A_630_74#_c_783_n N_A_1257_74#_c_965_n 0.00126251f $X=6.19 $Y=2.515
+ $X2=0 $Y2=0
cc_609 N_A_630_74#_c_784_n N_A_1257_74#_c_965_n 0.0187936f $X=7.93 $Y=2.6 $X2=0
+ $Y2=0
cc_610 N_A_630_74#_c_758_n N_A_1257_74#_c_961_n 0.00374483f $X=8.25 $Y=1.625
+ $X2=0 $Y2=0
cc_611 N_A_630_74#_c_764_n N_A_1257_74#_c_961_n 0.00265195f $X=8.115 $Y=1.79
+ $X2=0 $Y2=0
cc_612 N_A_630_74#_c_785_n N_A_1257_74#_c_961_n 0.00850637f $X=8.015 $Y=2.515
+ $X2=0 $Y2=0
cc_613 N_A_630_74#_c_772_n N_A_1257_74#_c_961_n 0.0175575f $X=7.935 $Y=1.79
+ $X2=0 $Y2=0
cc_614 N_A_630_74#_c_784_n N_A_1257_74#_c_1004_n 0.0369777f $X=7.93 $Y=2.6 $X2=0
+ $Y2=0
cc_615 N_A_630_74#_c_785_n N_A_1257_74#_c_1004_n 0.0135845f $X=8.015 $Y=2.515
+ $X2=0 $Y2=0
cc_616 N_A_630_74#_c_758_n N_A_1257_74#_c_962_n 8.555e-19 $X=8.25 $Y=1.625 $X2=0
+ $Y2=0
cc_617 N_A_630_74#_c_784_n N_A_1026_100#_c_1038_n 0.0173259f $X=7.93 $Y=2.6
+ $X2=0 $Y2=0
cc_618 N_A_630_74#_M1025_g N_A_1026_100#_c_1034_n 0.00335709f $X=5.055 $Y=0.71
+ $X2=0 $Y2=0
cc_619 N_A_630_74#_c_774_n N_A_1026_100#_c_1034_n 0.00134961f $X=5.905 $Y=1.755
+ $X2=0 $Y2=0
cc_620 N_A_630_74#_c_774_n N_A_1026_100#_c_1035_n 0.0206006f $X=5.905 $Y=1.755
+ $X2=0 $Y2=0
cc_621 N_A_630_74#_c_784_n N_A_1026_100#_c_1035_n 0.0081744f $X=7.93 $Y=2.6
+ $X2=0 $Y2=0
cc_622 N_A_630_74#_c_787_n N_A_1026_100#_c_1035_n 0.0260234f $X=6.19 $Y=2.115
+ $X2=0 $Y2=0
cc_623 N_A_630_74#_c_774_n N_A_1026_100#_c_1036_n 0.0109488f $X=5.905 $Y=1.755
+ $X2=0 $Y2=0
cc_624 N_A_630_74#_c_763_n N_A_1026_100#_c_1036_n 3.96092e-19 $X=5.055 $Y=1.555
+ $X2=0 $Y2=0
cc_625 N_A_630_74#_c_774_n N_A_1026_100#_c_1040_n 0.00365808f $X=5.905 $Y=1.755
+ $X2=0 $Y2=0
cc_626 N_A_630_74#_c_776_n N_A_1026_100#_c_1040_n 0.00910157f $X=5.995 $Y=2.455
+ $X2=0 $Y2=0
cc_627 N_A_630_74#_c_783_n N_A_1026_100#_c_1040_n 3.4062e-19 $X=6.19 $Y=2.515
+ $X2=0 $Y2=0
cc_628 N_A_630_74#_c_878_p N_A_1026_100#_c_1040_n 0.00714769f $X=6.275 $Y=2.6
+ $X2=0 $Y2=0
cc_629 N_A_630_74#_c_787_n N_A_1026_100#_c_1040_n 0.00117537f $X=6.19 $Y=2.115
+ $X2=0 $Y2=0
cc_630 N_A_630_74#_c_774_n N_A_1026_100#_c_1041_n 0.0078561f $X=5.905 $Y=1.755
+ $X2=0 $Y2=0
cc_631 N_A_630_74#_c_775_n N_A_1026_100#_c_1041_n 0.00994612f $X=6.07 $Y=2.115
+ $X2=0 $Y2=0
cc_632 N_A_630_74#_c_776_n N_A_1026_100#_c_1041_n 4.19687e-19 $X=5.995 $Y=2.455
+ $X2=0 $Y2=0
cc_633 N_A_630_74#_c_783_n N_A_1026_100#_c_1041_n 0.0102483f $X=6.19 $Y=2.515
+ $X2=0 $Y2=0
cc_634 N_A_630_74#_c_787_n N_A_1026_100#_c_1041_n 0.0248993f $X=6.19 $Y=2.115
+ $X2=0 $Y2=0
cc_635 N_A_630_74#_c_764_n N_A_1026_100#_c_1037_n 0.00850011f $X=8.115 $Y=1.79
+ $X2=0 $Y2=0
cc_636 N_A_630_74#_c_784_n N_A_1026_100#_c_1037_n 0.00118349f $X=7.93 $Y=2.6
+ $X2=0 $Y2=0
cc_637 N_A_630_74#_c_772_n N_A_1026_100#_c_1037_n 3.2502e-19 $X=7.935 $Y=1.79
+ $X2=0 $Y2=0
cc_638 N_A_630_74#_M1018_g N_A_1814_48#_c_1114_n 0.0210271f $X=8.755 $Y=0.58
+ $X2=0 $Y2=0
cc_639 N_A_630_74#_c_759_n N_A_1814_48#_c_1121_n 0.025472f $X=8.68 $Y=1.07 $X2=0
+ $Y2=0
cc_640 N_A_630_74#_c_757_n N_A_1587_74#_c_1281_n 0.0106328f $X=8.205 $Y=2.04
+ $X2=0 $Y2=0
cc_641 N_A_630_74#_M1018_g N_A_1587_74#_c_1272_n 0.0131812f $X=8.755 $Y=0.58
+ $X2=0 $Y2=0
cc_642 N_A_630_74#_c_757_n N_A_1587_74#_c_1283_n 0.00505228f $X=8.205 $Y=2.04
+ $X2=0 $Y2=0
cc_643 N_A_630_74#_c_785_n N_A_1587_74#_c_1283_n 0.0106703f $X=8.015 $Y=2.515
+ $X2=0 $Y2=0
cc_644 N_A_630_74#_c_759_n N_A_1587_74#_c_1273_n 0.00438494f $X=8.68 $Y=1.07
+ $X2=0 $Y2=0
cc_645 N_A_630_74#_M1018_g N_A_1587_74#_c_1273_n 0.0106668f $X=8.755 $Y=0.58
+ $X2=0 $Y2=0
cc_646 N_A_630_74#_c_759_n N_A_1587_74#_c_1274_n 0.0111704f $X=8.68 $Y=1.07
+ $X2=0 $Y2=0
cc_647 N_A_630_74#_c_760_n N_A_1587_74#_c_1274_n 0.00188364f $X=8.325 $Y=1.07
+ $X2=0 $Y2=0
cc_648 N_A_630_74#_c_758_n N_A_1587_74#_c_1275_n 0.00190634f $X=8.25 $Y=1.625
+ $X2=0 $Y2=0
cc_649 N_A_630_74#_c_759_n N_A_1587_74#_c_1275_n 0.00159758f $X=8.68 $Y=1.07
+ $X2=0 $Y2=0
cc_650 N_A_630_74#_c_781_n N_VPWR_M1017_s 0.00785452f $X=3.855 $Y=1.905 $X2=0
+ $Y2=0
cc_651 N_A_630_74#_c_784_n N_VPWR_M1026_d 0.0087397f $X=7.93 $Y=2.6 $X2=0 $Y2=0
cc_652 N_A_630_74#_c_784_n N_VPWR_c_1382_n 0.0250835f $X=7.93 $Y=2.6 $X2=0 $Y2=0
cc_653 N_A_630_74#_c_773_n N_VPWR_c_1394_n 0.00415318f $X=4.535 $Y=1.765 $X2=0
+ $Y2=0
cc_654 N_A_630_74#_c_776_n N_VPWR_c_1394_n 0.0055545f $X=5.995 $Y=2.455 $X2=0
+ $Y2=0
cc_655 N_A_630_74#_c_784_n N_VPWR_c_1394_n 0.00587216f $X=7.93 $Y=2.6 $X2=0
+ $Y2=0
cc_656 N_A_630_74#_c_878_p N_VPWR_c_1394_n 0.00290121f $X=6.275 $Y=2.6 $X2=0
+ $Y2=0
cc_657 N_A_630_74#_c_757_n N_VPWR_c_1395_n 0.00448506f $X=8.205 $Y=2.04 $X2=0
+ $Y2=0
cc_658 N_A_630_74#_c_784_n N_VPWR_c_1395_n 0.0176177f $X=7.93 $Y=2.6 $X2=0 $Y2=0
cc_659 N_A_630_74#_c_773_n N_VPWR_c_1398_n 0.025071f $X=4.535 $Y=1.765 $X2=0
+ $Y2=0
cc_660 N_A_630_74#_c_773_n N_VPWR_c_1380_n 0.00403216f $X=4.535 $Y=1.765 $X2=0
+ $Y2=0
cc_661 N_A_630_74#_c_776_n N_VPWR_c_1380_n 0.00580281f $X=5.995 $Y=2.455 $X2=0
+ $Y2=0
cc_662 N_A_630_74#_c_757_n N_VPWR_c_1380_n 0.00544287f $X=8.205 $Y=2.04 $X2=0
+ $Y2=0
cc_663 N_A_630_74#_c_784_n N_VPWR_c_1380_n 0.0432739f $X=7.93 $Y=2.6 $X2=0 $Y2=0
cc_664 N_A_630_74#_c_878_p N_VPWR_c_1380_n 0.00500266f $X=6.275 $Y=2.6 $X2=0
+ $Y2=0
cc_665 N_A_630_74#_c_765_n N_A_301_74#_c_1527_n 7.52944e-19 $X=3.29 $Y=0.515
+ $X2=0 $Y2=0
cc_666 N_A_630_74#_c_767_n N_A_301_74#_c_1527_n 0.00461766f $X=3.455 $Y=0.925
+ $X2=0 $Y2=0
cc_667 N_A_630_74#_c_786_n N_A_301_74#_c_1530_n 0.0242448f $X=3.49 $Y=1.905
+ $X2=0 $Y2=0
cc_668 N_A_630_74#_M1023_d N_A_301_74#_c_1535_n 0.00809453f $X=3.34 $Y=1.84
+ $X2=0 $Y2=0
cc_669 N_A_630_74#_c_781_n N_A_301_74#_c_1535_n 0.0218726f $X=3.855 $Y=1.905
+ $X2=0 $Y2=0
cc_670 N_A_630_74#_c_786_n N_A_301_74#_c_1535_n 0.0211124f $X=3.49 $Y=1.905
+ $X2=0 $Y2=0
cc_671 N_A_630_74#_c_754_n N_A_301_74#_c_1531_n 0.00156402f $X=4.445 $Y=1.555
+ $X2=0 $Y2=0
cc_672 N_A_630_74#_c_773_n N_A_301_74#_c_1531_n 0.0201921f $X=4.535 $Y=1.765
+ $X2=0 $Y2=0
cc_673 N_A_630_74#_c_762_n N_A_301_74#_c_1531_n 0.00516076f $X=4.535 $Y=1.555
+ $X2=0 $Y2=0
cc_674 N_A_630_74#_c_763_n N_A_301_74#_c_1531_n 6.79214e-19 $X=5.055 $Y=1.555
+ $X2=0 $Y2=0
cc_675 N_A_630_74#_c_781_n N_A_301_74#_c_1531_n 0.0135759f $X=3.855 $Y=1.905
+ $X2=0 $Y2=0
cc_676 N_A_630_74#_c_769_n N_A_301_74#_c_1531_n 0.0133694f $X=4.01 $Y=1.465
+ $X2=0 $Y2=0
cc_677 N_A_630_74#_c_754_n N_A_301_74#_c_1532_n 0.00624221f $X=4.445 $Y=1.555
+ $X2=0 $Y2=0
cc_678 N_A_630_74#_c_755_n N_A_301_74#_c_1532_n 0.0138473f $X=4.98 $Y=1.555
+ $X2=0 $Y2=0
cc_679 N_A_630_74#_c_762_n N_A_301_74#_c_1532_n 0.0153911f $X=4.535 $Y=1.555
+ $X2=0 $Y2=0
cc_680 N_A_630_74#_c_769_n N_A_301_74#_c_1532_n 0.0133606f $X=4.01 $Y=1.465
+ $X2=0 $Y2=0
cc_681 N_A_630_74#_M1019_g N_A_301_74#_c_1533_n 0.00351387f $X=4.065 $Y=0.74
+ $X2=0 $Y2=0
cc_682 N_A_630_74#_c_755_n N_A_301_74#_c_1533_n 0.00506057f $X=4.98 $Y=1.555
+ $X2=0 $Y2=0
cc_683 N_A_630_74#_M1025_g N_A_301_74#_c_1533_n 0.0124052f $X=5.055 $Y=0.71
+ $X2=0 $Y2=0
cc_684 N_A_630_74#_c_768_n N_A_301_74#_c_1533_n 0.00606886f $X=4.01 $Y=1.455
+ $X2=0 $Y2=0
cc_685 N_A_630_74#_c_770_n N_A_301_74#_c_1533_n 0.00320936f $X=4.01 $Y=1.465
+ $X2=0 $Y2=0
cc_686 N_A_630_74#_c_771_n N_A_301_74#_c_1533_n 0.00453071f $X=4.01 $Y=1.3 $X2=0
+ $Y2=0
cc_687 N_A_630_74#_c_773_n N_A_301_74#_c_1592_n 0.0175636f $X=4.535 $Y=1.765
+ $X2=0 $Y2=0
cc_688 N_A_630_74#_c_773_n N_A_301_74#_c_1539_n 0.00637121f $X=4.535 $Y=1.765
+ $X2=0 $Y2=0
cc_689 N_A_630_74#_c_784_n A_1214_506# 0.00227104f $X=7.93 $Y=2.6 $X2=-0.19
+ $Y2=-0.245
cc_690 N_A_630_74#_c_878_p A_1214_506# 0.00393591f $X=6.275 $Y=2.6 $X2=-0.19
+ $Y2=-0.245
cc_691 N_A_630_74#_c_766_n N_VGND_M1019_s 0.00884676f $X=3.855 $Y=0.925 $X2=0
+ $Y2=0
cc_692 N_A_630_74#_c_771_n N_VGND_M1019_s 0.0037774f $X=4.01 $Y=1.3 $X2=0 $Y2=0
cc_693 N_A_630_74#_c_765_n N_VGND_c_1734_n 0.0180182f $X=3.29 $Y=0.515 $X2=0
+ $Y2=0
cc_694 N_A_630_74#_M1019_g N_VGND_c_1735_n 0.00850533f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_695 N_A_630_74#_c_765_n N_VGND_c_1735_n 0.0215739f $X=3.29 $Y=0.515 $X2=0
+ $Y2=0
cc_696 N_A_630_74#_c_766_n N_VGND_c_1735_n 0.0222748f $X=3.855 $Y=0.925 $X2=0
+ $Y2=0
cc_697 N_A_630_74#_c_770_n N_VGND_c_1735_n 3.75969e-19 $X=4.01 $Y=1.465 $X2=0
+ $Y2=0
cc_698 N_A_630_74#_M1018_g N_VGND_c_1737_n 0.00167829f $X=8.755 $Y=0.58 $X2=0
+ $Y2=0
cc_699 N_A_630_74#_c_765_n N_VGND_c_1744_n 0.0145323f $X=3.29 $Y=0.515 $X2=0
+ $Y2=0
cc_700 N_A_630_74#_M1019_g N_VGND_c_1746_n 0.00383152f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_701 N_A_630_74#_M1025_g N_VGND_c_1746_n 7.26171e-19 $X=5.055 $Y=0.71 $X2=0
+ $Y2=0
cc_702 N_A_630_74#_M1018_g N_VGND_c_1748_n 0.00461464f $X=8.755 $Y=0.58 $X2=0
+ $Y2=0
cc_703 N_A_630_74#_M1019_g N_VGND_c_1756_n 0.00729907f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_704 N_A_630_74#_M1018_g N_VGND_c_1756_n 0.00914027f $X=8.755 $Y=0.58 $X2=0
+ $Y2=0
cc_705 N_A_630_74#_c_765_n N_VGND_c_1756_n 0.0119861f $X=3.29 $Y=0.515 $X2=0
+ $Y2=0
cc_706 N_A_630_74#_c_766_n N_VGND_c_1756_n 0.00942661f $X=3.855 $Y=0.925 $X2=0
+ $Y2=0
cc_707 N_A_1257_74#_c_958_n N_A_1026_100#_c_1038_n 0.0128668f $X=6.535 $Y=2.365
+ $X2=0 $Y2=0
cc_708 N_A_1257_74#_c_965_n N_A_1026_100#_c_1038_n 0.0145211f $X=6.535 $Y=2.455
+ $X2=0 $Y2=0
cc_709 N_A_1257_74#_c_961_n N_A_1026_100#_c_1038_n 0.00495033f $X=7.415 $Y=2.175
+ $X2=0 $Y2=0
cc_710 N_A_1257_74#_c_1004_n N_A_1026_100#_c_1038_n 0.00839121f $X=7.485 $Y=2.26
+ $X2=0 $Y2=0
cc_711 N_A_1257_74#_c_959_n N_A_1026_100#_M1035_g 0.0193438f $X=7.33 $Y=1.275
+ $X2=0 $Y2=0
cc_712 N_A_1257_74#_c_960_n N_A_1026_100#_M1035_g 0.00969358f $X=7.415 $Y=1.11
+ $X2=0 $Y2=0
cc_713 N_A_1257_74#_c_961_n N_A_1026_100#_M1035_g 0.00967622f $X=7.415 $Y=2.175
+ $X2=0 $Y2=0
cc_714 N_A_1257_74#_c_984_n N_A_1026_100#_M1035_g 0.00707154f $X=7.555 $Y=0.72
+ $X2=0 $Y2=0
cc_715 N_A_1257_74#_c_962_n N_A_1026_100#_M1035_g 0.00373289f $X=7.415 $Y=1.275
+ $X2=0 $Y2=0
cc_716 N_A_1257_74#_c_963_n N_A_1026_100#_M1035_g 0.00930171f $X=6.535 $Y=1.275
+ $X2=0 $Y2=0
cc_717 N_A_1257_74#_M1034_g N_A_1026_100#_c_1034_n 0.0017866f $X=6.36 $Y=0.71
+ $X2=0 $Y2=0
cc_718 N_A_1257_74#_c_958_n N_A_1026_100#_c_1035_n 0.0185001f $X=6.535 $Y=2.365
+ $X2=0 $Y2=0
cc_719 N_A_1257_74#_c_959_n N_A_1026_100#_c_1035_n 0.0664648f $X=7.33 $Y=1.275
+ $X2=0 $Y2=0
cc_720 N_A_1257_74#_c_961_n N_A_1026_100#_c_1035_n 0.0235372f $X=7.415 $Y=2.175
+ $X2=0 $Y2=0
cc_721 N_A_1257_74#_c_963_n N_A_1026_100#_c_1035_n 0.00422752f $X=6.535 $Y=1.275
+ $X2=0 $Y2=0
cc_722 N_A_1257_74#_c_965_n N_A_1026_100#_c_1040_n 0.00141443f $X=6.535 $Y=2.455
+ $X2=0 $Y2=0
cc_723 N_A_1257_74#_c_958_n N_A_1026_100#_c_1037_n 0.0253149f $X=6.535 $Y=2.365
+ $X2=0 $Y2=0
cc_724 N_A_1257_74#_c_959_n N_A_1026_100#_c_1037_n 0.00442607f $X=7.33 $Y=1.275
+ $X2=0 $Y2=0
cc_725 N_A_1257_74#_c_961_n N_A_1026_100#_c_1037_n 0.0128324f $X=7.415 $Y=2.175
+ $X2=0 $Y2=0
cc_726 N_A_1257_74#_c_1004_n N_A_1026_100#_c_1037_n 0.00261556f $X=7.485 $Y=2.26
+ $X2=0 $Y2=0
cc_727 N_A_1257_74#_c_965_n N_VPWR_c_1382_n 0.00649277f $X=6.535 $Y=2.455 $X2=0
+ $Y2=0
cc_728 N_A_1257_74#_c_965_n N_VPWR_c_1394_n 0.00438517f $X=6.535 $Y=2.455 $X2=0
+ $Y2=0
cc_729 N_A_1257_74#_c_965_n N_VPWR_c_1380_n 0.00542671f $X=6.535 $Y=2.455 $X2=0
+ $Y2=0
cc_730 N_A_1257_74#_M1034_g N_VGND_c_1736_n 0.00553953f $X=6.36 $Y=0.71 $X2=0
+ $Y2=0
cc_731 N_A_1257_74#_M1034_g N_VGND_c_1746_n 0.00487664f $X=6.36 $Y=0.71 $X2=0
+ $Y2=0
cc_732 N_A_1257_74#_M1034_g N_VGND_c_1756_n 0.00505379f $X=6.36 $Y=0.71 $X2=0
+ $Y2=0
cc_733 N_A_1026_100#_c_1038_n N_VPWR_c_1382_n 0.0066996f $X=7.155 $Y=2.04 $X2=0
+ $Y2=0
cc_734 N_A_1026_100#_c_1040_n N_VPWR_c_1394_n 0.0149647f $X=5.77 $Y=2.74 $X2=0
+ $Y2=0
cc_735 N_A_1026_100#_c_1038_n N_VPWR_c_1395_n 0.0032411f $X=7.155 $Y=2.04 $X2=0
+ $Y2=0
cc_736 N_A_1026_100#_c_1038_n N_VPWR_c_1380_n 0.00544287f $X=7.155 $Y=2.04 $X2=0
+ $Y2=0
cc_737 N_A_1026_100#_c_1040_n N_VPWR_c_1380_n 0.013003f $X=5.77 $Y=2.74 $X2=0
+ $Y2=0
cc_738 N_A_1026_100#_c_1040_n N_A_301_74#_c_1539_n 0.0329228f $X=5.77 $Y=2.74
+ $X2=0 $Y2=0
cc_739 N_A_1026_100#_M1035_g N_VGND_c_1736_n 0.00260166f $X=7.28 $Y=0.645 $X2=0
+ $Y2=0
cc_740 N_A_1026_100#_M1035_g N_VGND_c_1748_n 0.00284028f $X=7.28 $Y=0.645 $X2=0
+ $Y2=0
cc_741 N_A_1026_100#_M1035_g N_VGND_c_1756_n 0.00361049f $X=7.28 $Y=0.645 $X2=0
+ $Y2=0
cc_742 N_A_1814_48#_c_1115_n N_A_1587_74#_c_1267_n 0.0213701f $X=9.165 $Y=1.475
+ $X2=0 $Y2=0
cc_743 N_A_1814_48#_c_1116_n N_A_1587_74#_c_1267_n 0.0179787f $X=9.165 $Y=2.215
+ $X2=0 $Y2=0
cc_744 N_A_1814_48#_c_1129_n N_A_1587_74#_c_1267_n 0.0119201f $X=9.165 $Y=2.305
+ $X2=0 $Y2=0
cc_745 N_A_1814_48#_c_1124_n N_A_1587_74#_c_1267_n 0.00916312f $X=10.135
+ $Y=1.465 $X2=0 $Y2=0
cc_746 N_A_1814_48#_c_1126_n N_A_1587_74#_c_1267_n 0.0107699f $X=9.5 $Y=1.065
+ $X2=0 $Y2=0
cc_747 N_A_1814_48#_c_1134_n N_A_1587_74#_c_1267_n 0.0137249f $X=9.895 $Y=2.135
+ $X2=0 $Y2=0
cc_748 N_A_1814_48#_c_1135_n N_A_1587_74#_c_1267_n 0.00381127f $X=9.932 $Y=1.97
+ $X2=0 $Y2=0
cc_749 N_A_1814_48#_c_1124_n N_A_1587_74#_c_1268_n 0.00605989f $X=10.135
+ $Y=1.465 $X2=0 $Y2=0
cc_750 N_A_1814_48#_c_1134_n N_A_1587_74#_c_1268_n 0.00353734f $X=9.895 $Y=2.135
+ $X2=0 $Y2=0
cc_751 N_A_1814_48#_c_1130_n N_A_1587_74#_c_1269_n 0.0040171f $X=10.625 $Y=1.765
+ $X2=0 $Y2=0
cc_752 N_A_1814_48#_c_1125_n N_A_1587_74#_c_1269_n 0.00361976f $X=11.38 $Y=1.465
+ $X2=0 $Y2=0
cc_753 N_A_1814_48#_c_1135_n N_A_1587_74#_c_1269_n 0.00461962f $X=9.932 $Y=1.97
+ $X2=0 $Y2=0
cc_754 N_A_1814_48#_c_1130_n N_A_1587_74#_c_1280_n 0.00803968f $X=10.625
+ $Y=1.765 $X2=0 $Y2=0
cc_755 N_A_1814_48#_c_1134_n N_A_1587_74#_c_1280_n 0.0154789f $X=9.895 $Y=2.135
+ $X2=0 $Y2=0
cc_756 N_A_1814_48#_c_1135_n N_A_1587_74#_c_1280_n 0.00504194f $X=9.932 $Y=1.97
+ $X2=0 $Y2=0
cc_757 N_A_1814_48#_M1003_g N_A_1587_74#_M1027_g 0.0153489f $X=10.61 $Y=0.74
+ $X2=0 $Y2=0
cc_758 N_A_1814_48#_c_1123_n N_A_1587_74#_M1027_g 0.00205498f $X=9.92 $Y=0.515
+ $X2=0 $Y2=0
cc_759 N_A_1814_48#_c_1124_n N_A_1587_74#_M1027_g 0.0151138f $X=10.135 $Y=1.465
+ $X2=0 $Y2=0
cc_760 N_A_1814_48#_c_1125_n N_A_1587_74#_M1027_g 0.00626302f $X=11.38 $Y=1.465
+ $X2=0 $Y2=0
cc_761 N_A_1814_48#_c_1126_n N_A_1587_74#_M1027_g 0.00633351f $X=9.5 $Y=1.065
+ $X2=0 $Y2=0
cc_762 N_A_1814_48#_c_1124_n N_A_1587_74#_c_1271_n 0.00210457f $X=10.135
+ $Y=1.465 $X2=0 $Y2=0
cc_763 N_A_1814_48#_c_1125_n N_A_1587_74#_c_1271_n 0.00306956f $X=11.38 $Y=1.465
+ $X2=0 $Y2=0
cc_764 N_A_1814_48#_c_1127_n N_A_1587_74#_c_1271_n 0.0153489f $X=11.975 $Y=1.532
+ $X2=0 $Y2=0
cc_765 N_A_1814_48#_c_1116_n N_A_1587_74#_c_1282_n 0.0114703f $X=9.165 $Y=2.215
+ $X2=0 $Y2=0
cc_766 N_A_1814_48#_c_1134_n N_A_1587_74#_c_1282_n 0.0052631f $X=9.895 $Y=2.135
+ $X2=0 $Y2=0
cc_767 N_A_1814_48#_c_1121_n N_A_1587_74#_c_1273_n 0.012308f $X=9.07 $Y=0.9
+ $X2=0 $Y2=0
cc_768 N_A_1814_48#_c_1124_n N_A_1587_74#_c_1273_n 0.01358f $X=10.135 $Y=1.465
+ $X2=0 $Y2=0
cc_769 N_A_1814_48#_c_1115_n N_A_1587_74#_c_1275_n 0.00467978f $X=9.165 $Y=1.475
+ $X2=0 $Y2=0
cc_770 N_A_1814_48#_c_1121_n N_A_1587_74#_c_1275_n 0.00513059f $X=9.07 $Y=0.9
+ $X2=0 $Y2=0
cc_771 N_A_1814_48#_c_1122_n N_A_1587_74#_c_1275_n 0.00718932f $X=9.165 $Y=1.385
+ $X2=0 $Y2=0
cc_772 N_A_1814_48#_c_1124_n N_A_1587_74#_c_1275_n 0.0174825f $X=10.135 $Y=1.465
+ $X2=0 $Y2=0
cc_773 N_A_1814_48#_c_1116_n N_A_1587_74#_c_1284_n 0.00625387f $X=9.165 $Y=2.215
+ $X2=0 $Y2=0
cc_774 N_A_1814_48#_c_1134_n N_A_1587_74#_c_1284_n 0.00138238f $X=9.895 $Y=2.135
+ $X2=0 $Y2=0
cc_775 N_A_1814_48#_c_1115_n N_A_1587_74#_c_1276_n 0.00324185f $X=9.165 $Y=1.475
+ $X2=0 $Y2=0
cc_776 N_A_1814_48#_c_1116_n N_A_1587_74#_c_1276_n 0.00764798f $X=9.165 $Y=2.215
+ $X2=0 $Y2=0
cc_777 N_A_1814_48#_c_1124_n N_A_1587_74#_c_1276_n 0.0493324f $X=10.135 $Y=1.465
+ $X2=0 $Y2=0
cc_778 N_A_1814_48#_c_1126_n N_A_1587_74#_c_1276_n 0.0046291f $X=9.5 $Y=1.065
+ $X2=0 $Y2=0
cc_779 N_A_1814_48#_c_1134_n N_A_1587_74#_c_1276_n 0.00296045f $X=9.895 $Y=2.135
+ $X2=0 $Y2=0
cc_780 N_A_1814_48#_c_1135_n N_A_1587_74#_c_1276_n 0.013468f $X=9.932 $Y=1.97
+ $X2=0 $Y2=0
cc_781 N_A_1814_48#_c_1116_n N_A_1587_74#_c_1277_n 0.00444158f $X=9.165 $Y=2.215
+ $X2=0 $Y2=0
cc_782 N_A_1814_48#_c_1129_n N_VPWR_c_1383_n 0.0137754f $X=9.165 $Y=2.305 $X2=0
+ $Y2=0
cc_783 N_A_1814_48#_c_1134_n N_VPWR_c_1383_n 0.0181747f $X=9.895 $Y=2.135 $X2=0
+ $Y2=0
cc_784 N_A_1814_48#_c_1134_n N_VPWR_c_1384_n 0.0106053f $X=9.895 $Y=2.135 $X2=0
+ $Y2=0
cc_785 N_A_1814_48#_c_1130_n N_VPWR_c_1385_n 0.00963242f $X=10.625 $Y=1.765
+ $X2=0 $Y2=0
cc_786 N_A_1814_48#_c_1125_n N_VPWR_c_1385_n 0.00946188f $X=11.38 $Y=1.465 $X2=0
+ $Y2=0
cc_787 N_A_1814_48#_c_1135_n N_VPWR_c_1385_n 0.06581f $X=9.932 $Y=1.97 $X2=0
+ $Y2=0
cc_788 N_A_1814_48#_c_1130_n N_VPWR_c_1386_n 0.00445602f $X=10.625 $Y=1.765
+ $X2=0 $Y2=0
cc_789 N_A_1814_48#_c_1131_n N_VPWR_c_1386_n 0.00445602f $X=11.075 $Y=1.765
+ $X2=0 $Y2=0
cc_790 N_A_1814_48#_c_1131_n N_VPWR_c_1387_n 0.00630489f $X=11.075 $Y=1.765
+ $X2=0 $Y2=0
cc_791 N_A_1814_48#_c_1132_n N_VPWR_c_1387_n 0.0133451f $X=11.525 $Y=1.765 $X2=0
+ $Y2=0
cc_792 N_A_1814_48#_c_1133_n N_VPWR_c_1387_n 5.83721e-19 $X=11.975 $Y=1.765
+ $X2=0 $Y2=0
cc_793 N_A_1814_48#_c_1132_n N_VPWR_c_1389_n 5.45313e-19 $X=11.525 $Y=1.765
+ $X2=0 $Y2=0
cc_794 N_A_1814_48#_c_1133_n N_VPWR_c_1389_n 0.0158803f $X=11.975 $Y=1.765 $X2=0
+ $Y2=0
cc_795 N_A_1814_48#_c_1129_n N_VPWR_c_1395_n 0.00421101f $X=9.165 $Y=2.305 $X2=0
+ $Y2=0
cc_796 N_A_1814_48#_c_1132_n N_VPWR_c_1396_n 0.00413917f $X=11.525 $Y=1.765
+ $X2=0 $Y2=0
cc_797 N_A_1814_48#_c_1133_n N_VPWR_c_1396_n 0.00413917f $X=11.975 $Y=1.765
+ $X2=0 $Y2=0
cc_798 N_A_1814_48#_c_1129_n N_VPWR_c_1380_n 0.00450151f $X=9.165 $Y=2.305 $X2=0
+ $Y2=0
cc_799 N_A_1814_48#_c_1130_n N_VPWR_c_1380_n 0.00862615f $X=10.625 $Y=1.765
+ $X2=0 $Y2=0
cc_800 N_A_1814_48#_c_1131_n N_VPWR_c_1380_n 0.00857589f $X=11.075 $Y=1.765
+ $X2=0 $Y2=0
cc_801 N_A_1814_48#_c_1132_n N_VPWR_c_1380_n 0.00817726f $X=11.525 $Y=1.765
+ $X2=0 $Y2=0
cc_802 N_A_1814_48#_c_1133_n N_VPWR_c_1380_n 0.00817726f $X=11.975 $Y=1.765
+ $X2=0 $Y2=0
cc_803 N_A_1814_48#_c_1134_n N_VPWR_c_1380_n 0.0132771f $X=9.895 $Y=2.135 $X2=0
+ $Y2=0
cc_804 N_A_1814_48#_c_1130_n N_Q_c_1666_n 0.0116217f $X=10.625 $Y=1.765 $X2=0
+ $Y2=0
cc_805 N_A_1814_48#_c_1131_n N_Q_c_1666_n 0.0127044f $X=11.075 $Y=1.765 $X2=0
+ $Y2=0
cc_806 N_A_1814_48#_c_1132_n N_Q_c_1666_n 7.68479e-19 $X=11.525 $Y=1.765 $X2=0
+ $Y2=0
cc_807 N_A_1814_48#_M1003_g N_Q_c_1660_n 0.00635169f $X=10.61 $Y=0.74 $X2=0
+ $Y2=0
cc_808 N_A_1814_48#_c_1125_n N_Q_c_1660_n 0.0210846f $X=11.38 $Y=1.465 $X2=0
+ $Y2=0
cc_809 N_A_1814_48#_c_1127_n N_Q_c_1660_n 0.0043097f $X=11.975 $Y=1.532 $X2=0
+ $Y2=0
cc_810 N_A_1814_48#_M1003_g N_Q_c_1661_n 0.00486666f $X=10.61 $Y=0.74 $X2=0
+ $Y2=0
cc_811 N_A_1814_48#_M1013_g N_Q_c_1661_n 4.84228e-19 $X=11.125 $Y=0.74 $X2=0
+ $Y2=0
cc_812 N_A_1814_48#_M1013_g N_Q_c_1662_n 0.0146564f $X=11.125 $Y=0.74 $X2=0
+ $Y2=0
cc_813 N_A_1814_48#_M1015_g N_Q_c_1662_n 0.0158223f $X=11.555 $Y=0.74 $X2=0
+ $Y2=0
cc_814 N_A_1814_48#_c_1125_n N_Q_c_1662_n 0.0417005f $X=11.38 $Y=1.465 $X2=0
+ $Y2=0
cc_815 N_A_1814_48#_c_1127_n N_Q_c_1662_n 0.00226244f $X=11.975 $Y=1.532 $X2=0
+ $Y2=0
cc_816 N_A_1814_48#_c_1131_n N_Q_c_1667_n 0.0120074f $X=11.075 $Y=1.765 $X2=0
+ $Y2=0
cc_817 N_A_1814_48#_c_1132_n N_Q_c_1667_n 0.0139944f $X=11.525 $Y=1.765 $X2=0
+ $Y2=0
cc_818 N_A_1814_48#_c_1125_n N_Q_c_1667_n 0.0389377f $X=11.38 $Y=1.465 $X2=0
+ $Y2=0
cc_819 N_A_1814_48#_c_1127_n N_Q_c_1667_n 0.0097652f $X=11.975 $Y=1.532 $X2=0
+ $Y2=0
cc_820 N_A_1814_48#_c_1130_n N_Q_c_1668_n 0.00347745f $X=10.625 $Y=1.765 $X2=0
+ $Y2=0
cc_821 N_A_1814_48#_c_1131_n N_Q_c_1668_n 9.3899e-19 $X=11.075 $Y=1.765 $X2=0
+ $Y2=0
cc_822 N_A_1814_48#_c_1125_n N_Q_c_1668_n 0.0276943f $X=11.38 $Y=1.465 $X2=0
+ $Y2=0
cc_823 N_A_1814_48#_c_1135_n N_Q_c_1668_n 0.00404023f $X=9.932 $Y=1.97 $X2=0
+ $Y2=0
cc_824 N_A_1814_48#_c_1127_n N_Q_c_1668_n 0.00758706f $X=11.975 $Y=1.532 $X2=0
+ $Y2=0
cc_825 N_A_1814_48#_c_1132_n N_Q_c_1669_n 0.00410179f $X=11.525 $Y=1.765 $X2=0
+ $Y2=0
cc_826 N_A_1814_48#_c_1133_n N_Q_c_1669_n 3.7781e-19 $X=11.975 $Y=1.765 $X2=0
+ $Y2=0
cc_827 N_A_1814_48#_M1015_g N_Q_c_1663_n 3.99083e-19 $X=11.555 $Y=0.74 $X2=0
+ $Y2=0
cc_828 N_A_1814_48#_M1028_g N_Q_c_1663_n 3.99083e-19 $X=11.985 $Y=0.74 $X2=0
+ $Y2=0
cc_829 N_A_1814_48#_c_1133_n N_Q_c_1670_n 0.0150686f $X=11.975 $Y=1.765 $X2=0
+ $Y2=0
cc_830 N_A_1814_48#_c_1127_n N_Q_c_1670_n 0.00308272f $X=11.975 $Y=1.532 $X2=0
+ $Y2=0
cc_831 N_A_1814_48#_M1028_g N_Q_c_1664_n 0.0153204f $X=11.985 $Y=0.74 $X2=0
+ $Y2=0
cc_832 N_A_1814_48#_c_1127_n N_Q_c_1664_n 0.0012066f $X=11.975 $Y=1.532 $X2=0
+ $Y2=0
cc_833 N_A_1814_48#_c_1132_n Q 9.17756e-19 $X=11.525 $Y=1.765 $X2=0 $Y2=0
cc_834 N_A_1814_48#_M1015_g Q 0.00469124f $X=11.555 $Y=0.74 $X2=0 $Y2=0
cc_835 N_A_1814_48#_c_1133_n Q 0.00138329f $X=11.975 $Y=1.765 $X2=0 $Y2=0
cc_836 N_A_1814_48#_M1028_g Q 0.00698119f $X=11.985 $Y=0.74 $X2=0 $Y2=0
cc_837 N_A_1814_48#_c_1125_n Q 0.0226429f $X=11.38 $Y=1.465 $X2=0 $Y2=0
cc_838 N_A_1814_48#_c_1127_n Q 0.0360424f $X=11.975 $Y=1.532 $X2=0 $Y2=0
cc_839 N_A_1814_48#_c_1114_n N_VGND_c_1737_n 0.0130582f $X=9.145 $Y=0.9 $X2=0
+ $Y2=0
cc_840 N_A_1814_48#_c_1121_n N_VGND_c_1737_n 0.00473839f $X=9.07 $Y=0.9 $X2=0
+ $Y2=0
cc_841 N_A_1814_48#_c_1123_n N_VGND_c_1737_n 0.0193366f $X=9.92 $Y=0.515 $X2=0
+ $Y2=0
cc_842 N_A_1814_48#_c_1124_n N_VGND_c_1737_n 0.0142497f $X=10.135 $Y=1.465 $X2=0
+ $Y2=0
cc_843 N_A_1814_48#_c_1126_n N_VGND_c_1737_n 0.00133759f $X=9.5 $Y=1.065 $X2=0
+ $Y2=0
cc_844 N_A_1814_48#_M1003_g N_VGND_c_1738_n 0.00193914f $X=10.61 $Y=0.74 $X2=0
+ $Y2=0
cc_845 N_A_1814_48#_c_1123_n N_VGND_c_1738_n 0.0225498f $X=9.92 $Y=0.515 $X2=0
+ $Y2=0
cc_846 N_A_1814_48#_c_1125_n N_VGND_c_1738_n 0.0146017f $X=11.38 $Y=1.465 $X2=0
+ $Y2=0
cc_847 N_A_1814_48#_M1003_g N_VGND_c_1739_n 4.31406e-19 $X=10.61 $Y=0.74 $X2=0
+ $Y2=0
cc_848 N_A_1814_48#_M1013_g N_VGND_c_1739_n 0.00831568f $X=11.125 $Y=0.74 $X2=0
+ $Y2=0
cc_849 N_A_1814_48#_M1015_g N_VGND_c_1739_n 0.00791319f $X=11.555 $Y=0.74 $X2=0
+ $Y2=0
cc_850 N_A_1814_48#_M1028_g N_VGND_c_1739_n 4.27258e-19 $X=11.985 $Y=0.74 $X2=0
+ $Y2=0
cc_851 N_A_1814_48#_M1015_g N_VGND_c_1741_n 4.27258e-19 $X=11.555 $Y=0.74 $X2=0
+ $Y2=0
cc_852 N_A_1814_48#_M1028_g N_VGND_c_1741_n 0.00909727f $X=11.985 $Y=0.74 $X2=0
+ $Y2=0
cc_853 N_A_1814_48#_c_1114_n N_VGND_c_1748_n 0.00383152f $X=9.145 $Y=0.9 $X2=0
+ $Y2=0
cc_854 N_A_1814_48#_c_1123_n N_VGND_c_1749_n 0.00749631f $X=9.92 $Y=0.515 $X2=0
+ $Y2=0
cc_855 N_A_1814_48#_M1003_g N_VGND_c_1750_n 0.00461464f $X=10.61 $Y=0.74 $X2=0
+ $Y2=0
cc_856 N_A_1814_48#_M1013_g N_VGND_c_1750_n 0.00383152f $X=11.125 $Y=0.74 $X2=0
+ $Y2=0
cc_857 N_A_1814_48#_M1015_g N_VGND_c_1751_n 0.00383152f $X=11.555 $Y=0.74 $X2=0
+ $Y2=0
cc_858 N_A_1814_48#_M1028_g N_VGND_c_1751_n 0.00383152f $X=11.985 $Y=0.74 $X2=0
+ $Y2=0
cc_859 N_A_1814_48#_c_1114_n N_VGND_c_1756_n 0.0075725f $X=9.145 $Y=0.9 $X2=0
+ $Y2=0
cc_860 N_A_1814_48#_M1003_g N_VGND_c_1756_n 0.00908838f $X=10.61 $Y=0.74 $X2=0
+ $Y2=0
cc_861 N_A_1814_48#_M1013_g N_VGND_c_1756_n 0.00758328f $X=11.125 $Y=0.74 $X2=0
+ $Y2=0
cc_862 N_A_1814_48#_M1015_g N_VGND_c_1756_n 0.0075754f $X=11.555 $Y=0.74 $X2=0
+ $Y2=0
cc_863 N_A_1814_48#_M1028_g N_VGND_c_1756_n 0.0075754f $X=11.985 $Y=0.74 $X2=0
+ $Y2=0
cc_864 N_A_1814_48#_c_1123_n N_VGND_c_1756_n 0.0062048f $X=9.92 $Y=0.515 $X2=0
+ $Y2=0
cc_865 N_A_1587_74#_c_1267_n N_VPWR_c_1383_n 0.00718629f $X=9.67 $Y=1.885 $X2=0
+ $Y2=0
cc_866 N_A_1587_74#_c_1281_n N_VPWR_c_1383_n 0.012797f $X=8.435 $Y=2.26 $X2=0
+ $Y2=0
cc_867 N_A_1587_74#_c_1276_n N_VPWR_c_1383_n 0.011372f $X=9.63 $Y=1.635 $X2=0
+ $Y2=0
cc_868 N_A_1587_74#_c_1267_n N_VPWR_c_1384_n 0.00458031f $X=9.67 $Y=1.885 $X2=0
+ $Y2=0
cc_869 N_A_1587_74#_c_1280_n N_VPWR_c_1384_n 0.00398926f $X=10.12 $Y=1.885 $X2=0
+ $Y2=0
cc_870 N_A_1587_74#_c_1280_n N_VPWR_c_1385_n 0.00565056f $X=10.12 $Y=1.885 $X2=0
+ $Y2=0
cc_871 N_A_1587_74#_c_1281_n N_VPWR_c_1395_n 0.00780759f $X=8.435 $Y=2.26 $X2=0
+ $Y2=0
cc_872 N_A_1587_74#_c_1267_n N_VPWR_c_1380_n 0.0049649f $X=9.67 $Y=1.885 $X2=0
+ $Y2=0
cc_873 N_A_1587_74#_c_1280_n N_VPWR_c_1380_n 0.0049649f $X=10.12 $Y=1.885 $X2=0
+ $Y2=0
cc_874 N_A_1587_74#_c_1281_n N_VPWR_c_1380_n 0.0108373f $X=8.435 $Y=2.26 $X2=0
+ $Y2=0
cc_875 N_A_1587_74#_c_1280_n N_Q_c_1668_n 4.27663e-19 $X=10.12 $Y=1.885 $X2=0
+ $Y2=0
cc_876 N_A_1587_74#_M1027_g N_VGND_c_1737_n 0.00258825f $X=10.135 $Y=0.74 $X2=0
+ $Y2=0
cc_877 N_A_1587_74#_c_1272_n N_VGND_c_1737_n 0.0055977f $X=8.46 $Y=0.615 $X2=0
+ $Y2=0
cc_878 N_A_1587_74#_M1027_g N_VGND_c_1738_n 0.011506f $X=10.135 $Y=0.74 $X2=0
+ $Y2=0
cc_879 N_A_1587_74#_c_1272_n N_VGND_c_1748_n 0.0146971f $X=8.46 $Y=0.615 $X2=0
+ $Y2=0
cc_880 N_A_1587_74#_M1027_g N_VGND_c_1749_n 0.00383152f $X=10.135 $Y=0.74 $X2=0
+ $Y2=0
cc_881 N_A_1587_74#_M1027_g N_VGND_c_1756_n 0.00762539f $X=10.135 $Y=0.74 $X2=0
+ $Y2=0
cc_882 N_A_1587_74#_c_1272_n N_VGND_c_1756_n 0.012138f $X=8.46 $Y=0.615 $X2=0
+ $Y2=0
cc_883 N_VPWR_M1029_d N_A_301_74#_c_1541_n 0.0119505f $X=2.6 $Y=2.32 $X2=0 $Y2=0
cc_884 N_VPWR_c_1397_n N_A_301_74#_c_1541_n 0.0229891f $X=2.895 $Y=2.815 $X2=0
+ $Y2=0
cc_885 N_VPWR_c_1380_n N_A_301_74#_c_1541_n 0.0235529f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_886 N_VPWR_M1029_d N_A_301_74#_c_1530_n 0.0152167f $X=2.6 $Y=2.32 $X2=0 $Y2=0
cc_887 N_VPWR_M1029_d N_A_301_74#_c_1535_n 0.00131155f $X=2.6 $Y=2.32 $X2=0
+ $Y2=0
cc_888 N_VPWR_M1017_s N_A_301_74#_c_1535_n 0.0185716f $X=3.905 $Y=1.84 $X2=0
+ $Y2=0
cc_889 N_VPWR_c_1397_n N_A_301_74#_c_1535_n 0.0032171f $X=2.895 $Y=2.815 $X2=0
+ $Y2=0
cc_890 N_VPWR_c_1398_n N_A_301_74#_c_1535_n 0.0355337f $X=4.18 $Y=2.815 $X2=0
+ $Y2=0
cc_891 N_VPWR_c_1380_n N_A_301_74#_c_1535_n 0.0260298f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_892 N_VPWR_M1017_s N_A_301_74#_c_1531_n 0.0168186f $X=3.905 $Y=1.84 $X2=0
+ $Y2=0
cc_893 N_VPWR_c_1394_n N_A_301_74#_c_1537_n 0.00632494f $X=6.68 $Y=3.33 $X2=0
+ $Y2=0
cc_894 N_VPWR_c_1380_n N_A_301_74#_c_1537_n 0.00982281f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_895 N_VPWR_M1017_s N_A_301_74#_c_1592_n 7.26784e-19 $X=3.905 $Y=1.84 $X2=0
+ $Y2=0
cc_896 N_VPWR_c_1394_n N_A_301_74#_c_1592_n 0.00302042f $X=6.68 $Y=3.33 $X2=0
+ $Y2=0
cc_897 N_VPWR_c_1398_n N_A_301_74#_c_1592_n 0.00704814f $X=4.18 $Y=2.815 $X2=0
+ $Y2=0
cc_898 N_VPWR_c_1380_n N_A_301_74#_c_1592_n 0.0110509f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_899 N_VPWR_c_1381_n N_A_301_74#_c_1538_n 0.019773f $X=0.89 $Y=2.465 $X2=0
+ $Y2=0
cc_900 N_VPWR_c_1392_n N_A_301_74#_c_1538_n 0.0145363f $X=2.585 $Y=3.33 $X2=0
+ $Y2=0
cc_901 N_VPWR_c_1397_n N_A_301_74#_c_1538_n 0.0063504f $X=2.895 $Y=2.815 $X2=0
+ $Y2=0
cc_902 N_VPWR_c_1380_n N_A_301_74#_c_1538_n 0.011973f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_903 N_VPWR_M1029_d N_A_301_74#_c_1644_n 0.0025281f $X=2.6 $Y=2.32 $X2=0 $Y2=0
cc_904 N_VPWR_c_1397_n N_A_301_74#_c_1644_n 0.0147701f $X=2.895 $Y=2.815 $X2=0
+ $Y2=0
cc_905 N_VPWR_c_1380_n N_A_301_74#_c_1644_n 6.84279e-19 $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_906 N_VPWR_c_1394_n N_A_301_74#_c_1539_n 0.0102952f $X=6.68 $Y=3.33 $X2=0
+ $Y2=0
cc_907 N_VPWR_c_1380_n N_A_301_74#_c_1539_n 0.00896485f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_908 N_VPWR_c_1385_n N_Q_c_1666_n 0.0633647f $X=10.39 $Y=2.105 $X2=0 $Y2=0
cc_909 N_VPWR_c_1386_n N_Q_c_1666_n 0.014552f $X=11.215 $Y=3.33 $X2=0 $Y2=0
cc_910 N_VPWR_c_1387_n N_Q_c_1666_n 0.0563525f $X=11.3 $Y=2.305 $X2=0 $Y2=0
cc_911 N_VPWR_c_1380_n N_Q_c_1666_n 0.0119791f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_912 N_VPWR_M1006_d N_Q_c_1667_n 0.00222494f $X=11.15 $Y=1.84 $X2=0 $Y2=0
cc_913 N_VPWR_c_1387_n N_Q_c_1667_n 0.0154248f $X=11.3 $Y=2.305 $X2=0 $Y2=0
cc_914 N_VPWR_c_1385_n N_Q_c_1668_n 0.00200112f $X=10.39 $Y=2.105 $X2=0 $Y2=0
cc_915 N_VPWR_c_1387_n N_Q_c_1669_n 0.0540451f $X=11.3 $Y=2.305 $X2=0 $Y2=0
cc_916 N_VPWR_c_1389_n N_Q_c_1669_n 0.0291921f $X=12.2 $Y=2.27 $X2=0 $Y2=0
cc_917 N_VPWR_c_1396_n N_Q_c_1669_n 0.00838873f $X=12.035 $Y=3.33 $X2=0 $Y2=0
cc_918 N_VPWR_c_1380_n N_Q_c_1669_n 0.00694347f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_919 N_VPWR_M1033_d N_Q_c_1670_n 0.00366051f $X=12.05 $Y=1.84 $X2=0 $Y2=0
cc_920 N_VPWR_c_1389_n N_Q_c_1670_n 0.0234914f $X=12.2 $Y=2.27 $X2=0 $Y2=0
cc_921 N_A_301_74#_c_1541_n A_412_464# 0.0138302f $X=2.935 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_922 N_A_301_74#_c_1540_n N_VGND_c_1733_n 0.00833256f $X=2.365 $Y=0.515 $X2=0
+ $Y2=0
cc_923 N_A_301_74#_c_1527_n N_VGND_c_1734_n 0.00648541f $X=2.45 $Y=1.18 $X2=0
+ $Y2=0
cc_924 N_A_301_74#_c_1528_n N_VGND_c_1734_n 0.0116171f $X=2.935 $Y=1.265 $X2=0
+ $Y2=0
cc_925 N_A_301_74#_c_1540_n N_VGND_c_1742_n 0.0332162f $X=2.365 $Y=0.515 $X2=0
+ $Y2=0
cc_926 N_A_301_74#_c_1540_n N_VGND_c_1756_n 0.035888f $X=2.365 $Y=0.515 $X2=0
+ $Y2=0
cc_927 N_A_301_74#_c_1540_n A_452_74# 0.00345571f $X=2.365 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_928 N_A_301_74#_c_1527_n A_452_74# 0.00166604f $X=2.45 $Y=1.18 $X2=-0.19
+ $Y2=-0.245
cc_929 N_Q_c_1662_n N_VGND_M1013_d 0.00178571f $X=11.675 $Y=1.005 $X2=0 $Y2=0
cc_930 N_Q_c_1664_n N_VGND_M1028_d 0.00385981f $X=11.77 $Y=0.965 $X2=0 $Y2=0
cc_931 N_Q_c_1661_n N_VGND_c_1738_n 0.0169482f $X=10.91 $Y=0.515 $X2=0 $Y2=0
cc_932 N_Q_c_1661_n N_VGND_c_1739_n 0.0136308f $X=10.91 $Y=0.515 $X2=0 $Y2=0
cc_933 N_Q_c_1662_n N_VGND_c_1739_n 0.0175375f $X=11.675 $Y=1.005 $X2=0 $Y2=0
cc_934 N_Q_c_1663_n N_VGND_c_1739_n 0.0142351f $X=11.77 $Y=0.515 $X2=0 $Y2=0
cc_935 N_Q_c_1663_n N_VGND_c_1741_n 0.0142351f $X=11.77 $Y=0.515 $X2=0 $Y2=0
cc_936 N_Q_c_1664_n N_VGND_c_1741_n 0.0234832f $X=11.77 $Y=0.965 $X2=0 $Y2=0
cc_937 N_Q_c_1661_n N_VGND_c_1750_n 0.011066f $X=10.91 $Y=0.515 $X2=0 $Y2=0
cc_938 N_Q_c_1663_n N_VGND_c_1751_n 0.00838873f $X=11.77 $Y=0.515 $X2=0 $Y2=0
cc_939 N_Q_c_1661_n N_VGND_c_1756_n 0.00915947f $X=10.91 $Y=0.515 $X2=0 $Y2=0
cc_940 N_Q_c_1663_n N_VGND_c_1756_n 0.00694347f $X=11.77 $Y=0.515 $X2=0 $Y2=0
