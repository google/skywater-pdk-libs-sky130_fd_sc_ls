* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__or4b_2 A B C D_N VGND VNB VPB VPWR X
M1000 VPWR a_190_48# X VPB phighvt w=1.12e+06u l=150000u
+  ad=9.828e+11p pd=6.34e+06u as=3.36e+11p ps=2.84e+06u
M1001 a_190_48# a_27_368# a_638_392# VPB phighvt w=1e+06u l=150000u
+  ad=4.45e+11p pd=2.89e+06u as=3.9e+11p ps=2.78e+06u
M1002 a_190_48# C VGND VNB nshort w=640000u l=150000u
+  ad=4.896e+11p pd=4.09e+06u as=1.10645e+12p ps=8.83e+06u
M1003 a_190_48# A VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_190_48# VGND VNB nshort w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1005 VPWR D_N a_27_368# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1006 VGND B a_190_48# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_536_392# B a_452_392# VPB phighvt w=1e+06u l=150000u
+  ad=3.6e+11p pd=2.72e+06u as=2.7e+11p ps=2.54e+06u
M1008 a_638_392# C a_536_392# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND D_N a_27_368# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1010 VGND a_27_368# a_190_48# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_190_48# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_452_392# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_190_48# X VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
