# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__sedfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__sedfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.32000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.060000 0.835000 1.780000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.450000 2.085000 1.780000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.845000 0.620000 15.015000 1.820000 ;
        RECT 14.845000 1.820000 15.240000 2.980000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.860000 1.820000 16.235000 2.980000 ;
        RECT 15.875000 0.370000 16.235000 1.150000 ;
        RECT 16.065000 1.150000 16.235000 1.820000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.075000 1.180000 5.635000 1.510000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475000 1.450000 4.865000 1.780000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.575000 1.180000 7.075000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 16.320000 0.085000 ;
        RECT  1.150000  0.085000  1.480000 0.890000 ;
        RECT  2.210000  0.085000  2.540000 1.005000 ;
        RECT  4.910000  0.085000  5.240000 1.010000 ;
        RECT  6.380000  0.085000  6.550000 1.010000 ;
        RECT  7.290000  0.085000  7.620000 0.670000 ;
        RECT 10.065000  0.085000 10.390000 0.680000 ;
        RECT 11.580000  0.085000 11.830000 0.680000 ;
        RECT 13.190000  0.085000 14.035000 0.600000 ;
        RECT 15.525000  0.085000 15.695000 1.150000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
        RECT 15.995000 -0.085000 16.165000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 16.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 16.320000 3.415000 ;
        RECT  0.955000 2.630000  1.205000 3.245000 ;
        RECT  2.395000 2.650000  2.645000 3.245000 ;
        RECT  4.955000 2.630000  5.205000 3.245000 ;
        RECT  6.275000 2.650000  6.605000 3.245000 ;
        RECT  7.665000 2.650000  7.995000 3.245000 ;
        RECT 10.080000 2.730000 10.410000 3.245000 ;
        RECT 11.175000 2.730000 11.505000 3.245000 ;
        RECT 13.640000 2.650000 14.230000 3.245000 ;
        RECT 15.440000 1.820000 15.690000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
        RECT 15.035000 3.245000 15.205000 3.415000 ;
        RECT 15.515000 3.245000 15.685000 3.415000 ;
        RECT 15.995000 3.245000 16.165000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 16.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 0.480000  0.660000 0.810000 ;
      RECT  0.115000 0.810000  0.285000 2.290000 ;
      RECT  0.115000 2.290000  1.545000 2.460000 ;
      RECT  0.115000 2.460000  0.445000 2.980000 ;
      RECT  1.025000 1.110000  2.040000 1.280000 ;
      RECT  1.025000 1.280000  1.355000 1.950000 ;
      RECT  1.025000 1.950000  2.665000 2.120000 ;
      RECT  1.375000 2.460000  1.545000 2.905000 ;
      RECT  1.375000 2.905000  2.225000 3.075000 ;
      RECT  1.710000 0.545000  2.040000 1.110000 ;
      RECT  1.715000 2.120000  1.885000 2.735000 ;
      RECT  2.055000 2.310000  3.545000 2.480000 ;
      RECT  2.055000 2.480000  2.225000 2.905000 ;
      RECT  2.335000 1.525000  2.665000 1.950000 ;
      RECT  2.875000 1.525000  3.205000 2.140000 ;
      RECT  3.030000 0.545000  3.360000 1.175000 ;
      RECT  3.030000 1.175000  3.545000 1.345000 ;
      RECT  3.185000 2.480000  3.545000 2.980000 ;
      RECT  3.375000 1.345000  3.545000 2.310000 ;
      RECT  3.530000 0.545000  3.885000 1.005000 ;
      RECT  3.715000 1.005000  3.885000 2.300000 ;
      RECT  3.715000 2.300000  3.965000 2.905000 ;
      RECT  3.715000 2.905000  4.785000 3.075000 ;
      RECT  4.055000 0.410000  4.305000 0.605000 ;
      RECT  4.055000 0.605000  4.740000 1.065000 ;
      RECT  4.055000 1.065000  4.305000 1.950000 ;
      RECT  4.055000 1.950000  5.870000 2.120000 ;
      RECT  4.135000 2.120000  4.305000 2.290000 ;
      RECT  4.135000 2.290000  4.445000 2.735000 ;
      RECT  4.615000 2.290000  6.210000 2.310000 ;
      RECT  4.615000 2.310000  8.335000 2.460000 ;
      RECT  4.615000 2.460000  4.785000 2.905000 ;
      RECT  5.565000 1.790000  5.870000 1.950000 ;
      RECT  5.715000 2.460000  8.335000 2.480000 ;
      RECT  5.715000 2.480000  6.045000 2.970000 ;
      RECT  5.740000 0.605000  6.210000 1.010000 ;
      RECT  6.040000 1.010000  6.210000 2.290000 ;
      RECT  6.725000 1.820000  7.525000 2.140000 ;
      RECT  6.730000 0.350000  7.060000 0.840000 ;
      RECT  6.730000 0.840000  7.525000 1.010000 ;
      RECT  7.055000 1.810000  7.525000 1.820000 ;
      RECT  7.355000 1.010000  7.525000 1.810000 ;
      RECT  7.775000 1.480000  8.530000 1.650000 ;
      RECT  7.775000 1.650000  7.945000 2.310000 ;
      RECT  7.800000 0.255000  9.690000 0.425000 ;
      RECT  7.800000 0.425000  8.050000 1.130000 ;
      RECT  8.115000 1.820000  8.870000 2.140000 ;
      RECT  8.165000 2.480000  8.335000 2.730000 ;
      RECT  8.165000 2.730000  9.020000 2.980000 ;
      RECT  8.280000 0.595000  8.530000 1.480000 ;
      RECT  8.585000 2.140000  8.870000 2.380000 ;
      RECT  8.700000 0.425000  8.870000 1.820000 ;
      RECT  9.040000 0.620000  9.320000 0.950000 ;
      RECT  9.040000 0.950000  9.210000 1.620000 ;
      RECT  9.040000 1.620000 10.730000 1.790000 ;
      RECT  9.040000 1.790000  9.210000 2.390000 ;
      RECT  9.040000 2.390000  9.520000 2.560000 ;
      RECT  9.190000 2.560000  9.520000 2.980000 ;
      RECT  9.380000 1.120000  9.690000 1.450000 ;
      RECT  9.380000 1.960000  9.860000 2.220000 ;
      RECT  9.490000 0.425000  9.690000 0.850000 ;
      RECT  9.490000 0.850000 10.730000 1.020000 ;
      RECT  9.490000 1.020000  9.690000 1.120000 ;
      RECT  9.690000 2.220000  9.860000 2.390000 ;
      RECT  9.690000 2.390000 12.595000 2.560000 ;
      RECT  9.860000 1.190000 11.740000 1.360000 ;
      RECT  9.860000 1.360000 10.190000 1.450000 ;
      RECT 10.400000 1.530000 10.730000 1.620000 ;
      RECT 10.400000 1.790000 10.730000 1.830000 ;
      RECT 10.560000 0.255000 11.410000 0.425000 ;
      RECT 10.560000 0.425000 10.730000 0.850000 ;
      RECT 10.615000 2.050000 11.070000 2.220000 ;
      RECT 10.900000 0.595000 11.070000 1.190000 ;
      RECT 10.900000 1.360000 11.740000 1.520000 ;
      RECT 10.900000 1.520000 11.070000 2.050000 ;
      RECT 11.240000 0.425000 11.410000 0.850000 ;
      RECT 11.240000 0.850000 12.120000 1.020000 ;
      RECT 11.950000 1.020000 12.120000 1.130000 ;
      RECT 11.950000 1.130000 13.395000 1.300000 ;
      RECT 11.950000 1.300000 12.255000 1.800000 ;
      RECT 12.290000 0.350000 12.620000 0.770000 ;
      RECT 12.290000 0.770000 13.875000 0.940000 ;
      RECT 12.425000 1.470000 12.855000 1.800000 ;
      RECT 12.425000 1.800000 12.595000 2.390000 ;
      RECT 12.765000 2.520000 13.195000 2.980000 ;
      RECT 13.025000 1.715000 13.875000 1.885000 ;
      RECT 13.025000 1.885000 13.195000 2.520000 ;
      RECT 13.065000 1.300000 13.395000 1.545000 ;
      RECT 13.460000 2.055000 14.600000 2.380000 ;
      RECT 13.705000 0.940000 13.875000 1.200000 ;
      RECT 13.705000 1.200000 14.260000 1.530000 ;
      RECT 13.705000 1.530000 13.875000 1.715000 ;
      RECT 14.045000 1.920000 14.600000 2.055000 ;
      RECT 14.205000 0.255000 15.355000 0.425000 ;
      RECT 14.205000 0.425000 14.600000 1.030000 ;
      RECT 14.430000 1.030000 14.600000 1.920000 ;
      RECT 14.430000 2.380000 14.600000 2.980000 ;
      RECT 15.185000 0.425000 15.355000 1.320000 ;
      RECT 15.185000 1.320000 15.895000 1.650000 ;
    LAYER mcon ;
      RECT  3.035000 1.950000  3.205000 2.120000 ;
      RECT 14.075000 1.950000 14.245000 2.120000 ;
    LAYER met1 ;
      RECT  2.975000 1.920000  3.265000 1.965000 ;
      RECT  2.975000 1.965000 14.305000 2.105000 ;
      RECT  2.975000 2.105000  3.265000 2.150000 ;
      RECT 14.015000 1.920000 14.305000 1.965000 ;
      RECT 14.015000 2.105000 14.305000 2.150000 ;
  END
END sky130_fd_sc_ls__sedfxbp_1
