* File: sky130_fd_sc_ls__conb_1.pex.spice
* Created: Wed Sep  2 10:59:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__CONB_1%HI 1 2 3 4 5 12 14 15 19
r18 19 33 2.97405 $w=3.08e-07 $l=8e-08 $layer=LI1_cond $X=0.24 $Y=0.925 $X2=0.24
+ $Y2=0.845
r19 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.45
+ $Y=0.34 $X2=0.45 $Y2=0.34
r20 12 14 116.448 $w=5.1e-07 $l=1.11e-06 $layer=POLY_cond $X=0.36 $Y=1.45
+ $X2=0.36 $Y2=0.34
r21 4 5 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.665 $X2=0.24
+ $Y2=2.035
r22 3 4 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295 $X2=0.24
+ $Y2=1.665
r23 2 33 2.11141 $w=5.28e-07 $l=3e-09 $layer=LI1_cond $X=0.35 $Y=0.842 $X2=0.35
+ $Y2=0.845
r24 2 3 13.6806 $w=3.08e-07 $l=3.68e-07 $layer=LI1_cond $X=0.24 $Y=0.927
+ $X2=0.24 $Y2=1.295
r25 2 19 0.0743512 $w=3.08e-07 $l=2e-09 $layer=LI1_cond $X=0.24 $Y=0.927
+ $X2=0.24 $Y2=0.925
r26 1 2 6.47688 $w=5.28e-07 $l=2.87e-07 $layer=LI1_cond $X=0.35 $Y=0.555
+ $X2=0.35 $Y2=0.842
r27 1 15 4.85202 $w=5.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.35 $Y=0.555
+ $X2=0.35 $Y2=0.34
.ends

.subckt PM_SKY130_FD_SC_LS__CONB_1%VPWR 3 4 7 8 9 11 18 19
r19 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r20 15 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r21 9 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33 $X2=1.2
+ $Y2=3.33
r22 9 16 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r23 7 15 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=0.285 $Y=3.33 $X2=0.24
+ $Y2=3.33
r24 7 8 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.285 $Y=3.33 $X2=0.45
+ $Y2=3.33
r25 6 18 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.2 $Y2=3.33
r26 6 8 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33 $X2=0.45
+ $Y2=3.33
r27 4 11 116.448 $w=5.1e-07 $l=1.11e-06 $layer=POLY_cond $X=0.36 $Y=2.605
+ $X2=0.36 $Y2=1.495
r28 3 4 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.45 $Y=2.605
+ $X2=0.45 $Y2=2.605
r29 1 8 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.45 $Y=3.245 $X2=0.45
+ $Y2=3.33
r30 1 3 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=0.45 $Y=3.245 $X2=0.45
+ $Y2=2.605
.ends

.subckt PM_SKY130_FD_SC_LS__CONB_1%VGND 3 4 6 7 8 9 11 20
r17 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r18 9 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r19 9 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r20 7 15 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=0.825 $Y=0 $X2=0.72
+ $Y2=0
r21 7 8 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.825 $Y=0 $X2=0.99
+ $Y2=0
r22 6 19 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.2
+ $Y2=0
r23 6 8 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=0.99
+ $Y2=0
r24 4 11 118.546 $w=5.1e-07 $l=1.13e-06 $layer=POLY_cond $X=1.08 $Y=0.32
+ $X2=1.08 $Y2=1.45
r25 3 4 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.99 $Y=0.32
+ $X2=0.99 $Y2=0.32
r26 1 8 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=0.085 $X2=0.99
+ $Y2=0
r27 1 3 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.99 $Y=0.085
+ $X2=0.99 $Y2=0.32
.ends

.subckt PM_SKY130_FD_SC_LS__CONB_1%LO 1 2 3 4 5 12 14 27
r19 27 29 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=1.205 $Y=2.405
+ $X2=1.205 $Y2=2.485
r20 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.99
+ $Y=2.605 $X2=0.99 $Y2=2.605
r21 12 14 116.448 $w=5.1e-07 $l=1.11e-06 $layer=POLY_cond $X=1.08 $Y=1.495
+ $X2=1.08 $Y2=2.605
r22 5 15 3.83648 $w=5.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.09 $Y=2.775
+ $X2=1.09 $Y2=2.605
r23 4 15 2.66297 $w=5.28e-07 $l=1.18e-07 $layer=LI1_cond $X=1.09 $Y=2.487
+ $X2=1.09 $Y2=2.605
r24 4 29 2.27911 $w=5.28e-07 $l=2e-09 $layer=LI1_cond $X=1.09 $Y=2.487 $X2=1.09
+ $Y2=2.485
r25 4 27 0.115244 $w=2.98e-07 $l=3e-09 $layer=LI1_cond $X=1.205 $Y=2.402
+ $X2=1.205 $Y2=2.405
r26 3 4 14.0982 $w=2.98e-07 $l=3.67e-07 $layer=LI1_cond $X=1.205 $Y=2.035
+ $X2=1.205 $Y2=2.402
r27 2 3 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.205 $Y=1.665
+ $X2=1.205 $Y2=2.035
r28 1 2 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.205 $Y=1.295
+ $X2=1.205 $Y2=1.665
.ends

