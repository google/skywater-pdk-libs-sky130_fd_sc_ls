* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_30_368# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 a_27_74# B1 a_834_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 a_30_368# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 a_834_74# C1 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X6 Y A2 a_30_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 Y C1 a_834_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X9 a_30_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X10 a_834_74# B1 a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X11 a_834_74# C1 Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X12 a_834_74# B1 a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X13 Y A2 a_30_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X14 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X15 a_30_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X16 Y C1 a_834_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X18 a_27_74# B1 a_834_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X19 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X20 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X21 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X23 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X24 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X25 VPWR A1 a_30_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X26 VPWR A1 a_30_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X27 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends
