* File: sky130_fd_sc_ls__xor2_2.pex.spice
* Created: Wed Sep  2 11:31:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__XOR2_2%A 2 3 5 8 12 14 16 19 21 23 26 28 29 31 32 39
+ 40 46
c105 29 0 1.24099e-19 $X=2.35 $Y=1.515
c106 28 0 7.27408e-20 $X=2.35 $Y=1.515
c107 14 0 9.04372e-20 $X=1.935 $Y=1.765
c108 12 0 3.01101e-20 $X=1.92 $Y=0.74
r109 42 43 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=1.92 $Y=1.557
+ $X2=1.935 $Y2=1.557
r110 38 40 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.75 $Y=1.33 $X2=0.84
+ $Y2=1.33
r111 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.33 $X2=0.75 $Y2=1.33
r112 35 38 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=0.505 $Y=1.33
+ $X2=0.75 $Y2=1.33
r113 32 46 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=1.705
+ $X2=0.75 $Y2=1.62
r114 32 46 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=0.75 $Y=1.6 $X2=0.75
+ $Y2=1.62
r115 32 39 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=0.75 $Y=1.6
+ $X2=0.75 $Y2=1.33
r116 29 45 10.9253 $w=3.75e-07 $l=8.5e-08 $layer=POLY_cond $X=2.35 $Y=1.557
+ $X2=2.435 $Y2=1.557
r117 29 43 53.3413 $w=3.75e-07 $l=4.15e-07 $layer=POLY_cond $X=2.35 $Y=1.557
+ $X2=1.935 $Y2=1.557
r118 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.35
+ $Y=1.515 $X2=2.35 $Y2=1.515
r119 26 31 10.2759 $w=4.38e-07 $l=2.2e-07 $layer=LI1_cond $X=2.065 $Y=1.57
+ $X2=1.845 $Y2=1.57
r120 26 28 7.46469 $w=4.38e-07 $l=2.85e-07 $layer=LI1_cond $X=2.065 $Y=1.57
+ $X2=2.35 $Y2=1.57
r121 25 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=1.705
+ $X2=0.75 $Y2=1.705
r122 25 31 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=0.915 $Y=1.705
+ $X2=1.845 $Y2=1.705
r123 21 45 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.435 $Y=1.765
+ $X2=2.435 $Y2=1.557
r124 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.435 $Y=1.765
+ $X2=2.435 $Y2=2.4
r125 17 29 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=1.35
+ $X2=2.35 $Y2=1.557
r126 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.35 $Y=1.35
+ $X2=2.35 $Y2=0.74
r127 14 43 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.935 $Y=1.765
+ $X2=1.935 $Y2=1.557
r128 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.935 $Y=1.765
+ $X2=1.935 $Y2=2.4
r129 10 42 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.92 $Y=1.35
+ $X2=1.92 $Y2=1.557
r130 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.92 $Y=1.35
+ $X2=1.92 $Y2=0.74
r131 6 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.165
+ $X2=0.84 $Y2=1.33
r132 6 8 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=0.84 $Y=1.165
+ $X2=0.84 $Y2=0.69
r133 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.46
r134 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.795
+ $X2=0.505 $Y2=1.885
r135 1 35 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.495
+ $X2=0.505 $Y2=1.33
r136 1 2 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=0.505 $Y=1.495
+ $X2=0.505 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_2%B 1 3 4 5 7 10 11 13 14 16 17 19 20 22 25 29
+ 31 34 40 41 44
c118 34 0 3.01111e-20 $X=1.32 $Y=1.12
c119 25 0 1.24099e-19 $X=1.32 $Y=1.095
r120 41 42 2.23148 $w=4.32e-07 $l=2e-08 $layer=POLY_cond $X=4.285 $Y=1.492
+ $X2=4.305 $Y2=1.492
r121 39 41 34.0301 $w=4.32e-07 $l=3.05e-07 $layer=POLY_cond $X=3.98 $Y=1.492
+ $X2=4.285 $Y2=1.492
r122 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.98
+ $Y=1.385 $X2=3.98 $Y2=1.385
r123 37 39 21.7569 $w=4.32e-07 $l=1.95e-07 $layer=POLY_cond $X=3.785 $Y=1.492
+ $X2=3.98 $Y2=1.492
r124 36 37 8.36806 $w=4.32e-07 $l=7.5e-08 $layer=POLY_cond $X=3.71 $Y=1.492
+ $X2=3.785 $Y2=1.492
r125 31 40 8.41685 $w=5.38e-07 $l=3.8e-07 $layer=LI1_cond $X=3.6 $Y=1.28
+ $X2=3.98 $Y2=1.28
r126 31 44 8.66048 $w=5.38e-07 $l=1.15e-07 $layer=LI1_cond $X=3.6 $Y=1.28
+ $X2=3.485 $Y2=1.28
r127 29 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.32 $Y=1.285
+ $X2=1.32 $Y2=1.45
r128 29 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.32 $Y=1.285
+ $X2=1.32 $Y2=1.12
r129 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.32
+ $Y=1.285 $X2=1.32 $Y2=1.285
r130 25 28 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.32 $Y=1.095
+ $X2=1.32 $Y2=1.285
r131 24 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=1.095
+ $X2=1.32 $Y2=1.095
r132 24 44 130.481 $w=1.68e-07 $l=2e-06 $layer=LI1_cond $X=1.485 $Y=1.095
+ $X2=3.485 $Y2=1.095
r133 20 42 27.7542 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.305 $Y=1.22
+ $X2=4.305 $Y2=1.492
r134 20 22 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.305 $Y=1.22
+ $X2=4.305 $Y2=0.74
r135 17 41 27.7542 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.285 $Y=1.765
+ $X2=4.285 $Y2=1.492
r136 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.285 $Y=1.765
+ $X2=4.285 $Y2=2.4
r137 14 37 27.7542 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.785 $Y=1.765
+ $X2=3.785 $Y2=1.492
r138 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.785 $Y=1.765
+ $X2=3.785 $Y2=2.4
r139 11 36 27.7542 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.71 $Y=1.22
+ $X2=3.71 $Y2=1.492
r140 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.71 $Y=1.22
+ $X2=3.71 $Y2=0.74
r141 10 34 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.27 $Y=0.69
+ $X2=1.27 $Y2=1.12
r142 7 35 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.23 $Y=1.735
+ $X2=1.23 $Y2=1.45
r143 4 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.155 $Y=1.81
+ $X2=1.23 $Y2=1.735
r144 4 5 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.155 $Y=1.81 $X2=1
+ $Y2=1.81
r145 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.925 $Y=1.885
+ $X2=1 $Y2=1.81
r146 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.925 $Y=1.885
+ $X2=0.925 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_2%A_183_74# 1 2 7 9 12 14 16 18 19 20 21 22 25
+ 27 30 32 37 41 46
c113 19 0 3.01111e-20 $X=0.89 $Y=0.755
c114 7 0 7.27408e-20 $X=2.885 $Y=1.765
r115 46 47 7.01323 $w=3.78e-07 $l=5.5e-08 $layer=POLY_cond $X=3.28 $Y=1.557
+ $X2=3.335 $Y2=1.557
r116 42 46 40.8042 $w=3.78e-07 $l=3.2e-07 $layer=POLY_cond $X=2.96 $Y=1.557
+ $X2=3.28 $Y2=1.557
r117 42 44 9.56349 $w=3.78e-07 $l=7.5e-08 $layer=POLY_cond $X=2.96 $Y=1.557
+ $X2=2.885 $Y2=1.557
r118 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.96
+ $Y=1.515 $X2=2.96 $Y2=1.515
r119 38 41 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.77 $Y=1.515
+ $X2=2.96 $Y2=1.515
r120 32 34 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.055 $Y=0.595
+ $X2=1.055 $Y2=0.755
r121 29 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.77 $Y=1.68
+ $X2=2.77 $Y2=1.515
r122 29 30 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.77 $Y=1.68
+ $X2=2.77 $Y2=1.96
r123 28 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.315 $Y=2.045
+ $X2=1.19 $Y2=2.045
r124 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.685 $Y=2.045
+ $X2=2.77 $Y2=1.96
r125 27 28 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=2.685 $Y=2.045
+ $X2=1.315 $Y2=2.045
r126 23 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=2.13
+ $X2=1.19 $Y2=2.045
r127 23 25 31.5769 $w=2.48e-07 $l=6.85e-07 $layer=LI1_cond $X=1.19 $Y=2.13
+ $X2=1.19 $Y2=2.815
r128 21 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.065 $Y=2.045
+ $X2=1.19 $Y2=2.045
r129 21 22 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.065 $Y=2.045
+ $X2=0.415 $Y2=2.045
r130 19 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=0.755
+ $X2=1.055 $Y2=0.755
r131 19 20 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=0.89 $Y=0.755
+ $X2=0.415 $Y2=0.755
r132 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.33 $Y=1.96
+ $X2=0.415 $Y2=2.045
r133 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.33 $Y=0.84
+ $X2=0.415 $Y2=0.755
r134 17 18 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=0.33 $Y=0.84
+ $X2=0.33 $Y2=1.96
r135 14 47 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.335 $Y=1.765
+ $X2=3.335 $Y2=1.557
r136 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.335 $Y=1.765
+ $X2=3.335 $Y2=2.4
r137 10 46 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.28 $Y=1.35
+ $X2=3.28 $Y2=1.557
r138 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.28 $Y=1.35
+ $X2=3.28 $Y2=0.74
r139 7 44 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.885 $Y=1.765
+ $X2=2.885 $Y2=1.557
r140 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.885 $Y=1.765
+ $X2=2.885 $Y2=2.4
r141 2 37 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=1 $Y=1.96
+ $X2=1.15 $Y2=2.125
r142 2 25 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=1.96 $X2=1.15 $Y2=2.815
r143 1 32 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=0.915
+ $Y=0.37 $X2=1.055 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_2%VPWR 1 2 3 10 12 16 20 22 24 32 42 43 49 52
r59 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r61 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r62 43 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r63 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r64 40 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.175 $Y=3.33
+ $X2=4.01 $Y2=3.33
r65 40 42 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.175 $Y=3.33
+ $X2=4.56 $Y2=3.33
r66 39 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r67 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r68 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r69 35 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r70 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r71 33 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.16 $Y2=3.33
r72 33 35 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.64 $Y2=3.33
r73 32 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.845 $Y=3.33
+ $X2=4.01 $Y2=3.33
r74 32 38 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.845 $Y=3.33
+ $X2=3.6 $Y2=3.33
r75 31 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r76 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r77 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r78 28 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r79 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r80 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r81 25 46 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r82 25 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r83 24 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.16 $Y2=3.33
r84 24 30 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r85 22 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r86 22 50 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r87 18 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.01 $Y=3.245
+ $X2=4.01 $Y2=3.33
r88 18 20 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=4.01 $Y=3.245 $X2=4.01
+ $Y2=2.645
r89 14 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=3.245
+ $X2=2.16 $Y2=3.33
r90 14 16 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.16 $Y=3.245
+ $X2=2.16 $Y2=2.81
r91 10 46 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r92 10 12 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.465
r93 3 20 600 $w=1.7e-07 $l=8.76798e-07 $layer=licon1_PDIFF $count=1 $X=3.86
+ $Y=1.84 $X2=4.01 $Y2=2.645
r94 2 16 600 $w=1.7e-07 $l=1.04231e-06 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.84 $X2=2.16 $Y2=2.81
r95 1 12 300 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_2%A_313_368# 1 2 3 4 15 17 18 19 20 21 24 25 30
+ 36
c60 20 0 9.04372e-20 $X=2.825 $Y=2.99
c61 4 0 5.47968e-20 $X=4.36 $Y=1.84
r62 26 34 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.675 $Y=2.275
+ $X2=3.535 $Y2=2.275
r63 25 36 5.2341 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.345 $Y=2.275
+ $X2=4.515 $Y2=2.275
r64 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.345 $Y=2.275
+ $X2=3.675 $Y2=2.275
r65 22 24 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=3.535 $Y=2.905
+ $X2=3.535 $Y2=2.815
r66 21 34 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=2.36
+ $X2=3.535 $Y2=2.275
r67 21 24 18.7272 $w=2.78e-07 $l=4.55e-07 $layer=LI1_cond $X=3.535 $Y=2.36
+ $X2=3.535 $Y2=2.815
r68 19 22 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.395 $Y=2.99
+ $X2=3.535 $Y2=2.905
r69 19 20 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.395 $Y=2.99
+ $X2=2.825 $Y2=2.99
r70 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.66 $Y=2.905
+ $X2=2.825 $Y2=2.99
r71 17 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=2.47 $X2=2.66
+ $Y2=2.385
r72 17 18 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.66 $Y=2.47
+ $X2=2.66 $Y2=2.905
r73 16 30 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.795 $Y=2.385
+ $X2=1.67 $Y2=2.385
r74 15 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.495 $Y=2.385
+ $X2=2.66 $Y2=2.385
r75 15 16 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.495 $Y=2.385
+ $X2=1.795 $Y2=2.385
r76 4 36 300 $w=1.7e-07 $l=5.06606e-07 $layer=licon1_PDIFF $count=2 $X=4.36
+ $Y=1.84 $X2=4.515 $Y2=2.275
r77 3 34 600 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=1.84 $X2=3.56 $Y2=2.275
r78 3 24 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=1.84 $X2=3.56 $Y2=2.815
r79 2 32 300 $w=1.7e-07 $l=6.95971e-07 $layer=licon1_PDIFF $count=2 $X=2.51
+ $Y=1.84 $X2=2.66 $Y2=2.465
r80 1 30 300 $w=1.7e-07 $l=6.93722e-07 $layer=licon1_PDIFF $count=2 $X=1.565
+ $Y=1.84 $X2=1.71 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_2%X 1 2 3 12 14 17 21 23 24 25 26
c55 24 0 5.47968e-20 $X=4.56 $Y=0.925
r56 25 26 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.52 $Y=1.295
+ $X2=4.52 $Y2=1.665
r57 24 25 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.52 $Y=0.925
+ $X2=4.52 $Y2=1.295
r58 23 24 4.31269 $w=5e-07 $l=2.64244e-07 $layer=LI1_cond $X=4.52 $Y=0.595
+ $X2=4.56 $Y2=0.84
r59 22 26 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.52 $Y=1.85
+ $X2=4.52 $Y2=1.665
r60 19 21 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=3.495 $Y=0.717
+ $X2=3.66 $Y2=0.717
r61 14 23 4.91798 $w=1.7e-07 $l=2.31571e-07 $layer=LI1_cond $X=4.355 $Y=0.755
+ $X2=4.52 $Y2=0.595
r62 14 21 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.355 $Y=0.755
+ $X2=3.66 $Y2=0.755
r63 13 17 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.195 $Y=1.935
+ $X2=3.11 $Y2=1.935
r64 12 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.355 $Y=1.935
+ $X2=4.52 $Y2=1.85
r65 12 13 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=4.355 $Y=1.935
+ $X2=3.195 $Y2=1.935
r66 3 17 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=2.96
+ $Y=1.84 $X2=3.11 $Y2=2.015
r67 2 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.38
+ $Y=0.37 $X2=4.52 $Y2=0.515
r68 1 19 182 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=1 $X=3.355
+ $Y=0.37 $X2=3.495 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_2%VGND 1 2 3 12 16 19 20 21 23 27 36 37 45
r67 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r68 40 43 4.01161 $w=5.17e-07 $l=1.7e-07 $layer=LI1_cond $X=0.24 $Y=0.207
+ $X2=0.41 $Y2=0.207
r69 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r70 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r71 34 37 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r72 34 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r73 33 36 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r74 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r75 31 45 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.82 $Y=0 $X2=2.65
+ $Y2=0
r76 31 33 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.82 $Y=0 $X2=3.12
+ $Y2=0
r77 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r78 27 45 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.48 $Y=0 $X2=2.65
+ $Y2=0
r79 27 29 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.48 $Y=0 $X2=2.16
+ $Y2=0
r80 26 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r81 26 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r82 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r83 23 43 13.0006 $w=5.17e-07 $l=3.9e-07 $layer=LI1_cond $X=0.71 $Y=0 $X2=0.41
+ $Y2=0.207
r84 23 25 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=0.71 $Y=0 $X2=1.2
+ $Y2=0
r85 21 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r86 21 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r87 19 25 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.39 $Y=0 $X2=1.2
+ $Y2=0
r88 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=0 $X2=1.555
+ $Y2=0
r89 18 29 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.72 $Y=0 $X2=2.16
+ $Y2=0
r90 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=0 $X2=1.555
+ $Y2=0
r91 14 45 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=0.085
+ $X2=2.65 $Y2=0
r92 14 16 8.47385 $w=3.38e-07 $l=2.5e-07 $layer=LI1_cond $X=2.65 $Y=0.085
+ $X2=2.65 $Y2=0.335
r93 10 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=0.085
+ $X2=1.555 $Y2=0
r94 10 12 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.555 $Y=0.085
+ $X2=1.555 $Y2=0.595
r95 3 16 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.37 $X2=2.65 $Y2=0.335
r96 2 12 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=1.345
+ $Y=0.37 $X2=1.555 $Y2=0.595
r97 1 43 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.19 $X2=0.41 $Y2=0.335
.ends

.subckt PM_SKY130_FD_SC_LS__XOR2_2%A_399_74# 1 2 7 10 12 14 19 20
c39 7 0 3.01101e-20 $X=2.99 $Y=0.755
r40 19 20 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=4.005 $Y=0.377
+ $X2=3.84 $Y2=0.377
r41 14 16 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.135 $Y=0.595
+ $X2=2.135 $Y2=0.755
r42 12 20 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.16 $Y=0.34
+ $X2=3.84 $Y2=0.34
r43 9 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.075 $Y=0.425
+ $X2=3.16 $Y2=0.34
r44 9 10 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.075 $Y=0.425
+ $X2=3.075 $Y2=0.67
r45 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.3 $Y=0.755
+ $X2=2.135 $Y2=0.755
r46 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.99 $Y=0.755
+ $X2=3.075 $Y2=0.67
r47 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.99 $Y=0.755 $X2=2.3
+ $Y2=0.755
r48 2 19 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=3.785
+ $Y=0.37 $X2=4.005 $Y2=0.415
r49 1 14 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=1.995
+ $Y=0.37 $X2=2.135 $Y2=0.595
.ends

