* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_258_392# A2_N a_257_126# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_605_126# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 a_530_392# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 X a_93_264# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 a_93_264# a_257_126# a_530_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VPWR A1_N a_258_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND A1_N a_257_126# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X7 VGND a_257_126# a_93_264# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 a_257_126# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X9 VPWR B1 a_530_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_93_264# B2 a_605_126# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 X a_93_264# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
.ends
