# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__nor2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ls__nor2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.755000 1.780000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.530000 1.470000 0.860000 1.800000 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  0.824400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 0.350000 1.815000 0.960000 ;
        RECT 1.645000 0.960000 2.745000 1.010000 ;
        RECT 1.645000 1.010000 3.235000 1.180000 ;
        RECT 1.645000 1.180000 1.820000 2.735000 ;
        RECT 2.495000 0.350000 2.745000 0.960000 ;
        RECT 3.005000 1.180000 3.235000 1.410000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.110000  0.450000 0.780000 1.130000 ;
      RECT 0.110000  1.130000 1.475000 1.300000 ;
      RECT 0.110000  1.300000 0.360000 2.980000 ;
      RECT 0.560000  1.970000 0.890000 3.245000 ;
      RECT 0.985000  0.085000 1.315000 0.960000 ;
      RECT 1.120000  1.820000 1.450000 2.905000 ;
      RECT 1.120000  2.905000 2.350000 3.075000 ;
      RECT 1.145000  1.300000 1.475000 1.550000 ;
      RECT 1.985000  0.085000 2.315000 0.790000 ;
      RECT 2.020000  1.950000 3.250000 2.120000 ;
      RECT 2.020000  2.120000 2.350000 2.905000 ;
      RECT 2.550000  2.290000 2.800000 3.245000 ;
      RECT 2.915000  0.085000 3.245000 0.840000 ;
      RECT 3.000000  1.820000 3.250000 1.950000 ;
      RECT 3.000000  2.120000 3.250000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_ls__nor2b_2
END LIBRARY
