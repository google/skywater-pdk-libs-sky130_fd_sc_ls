* File: sky130_fd_sc_ls__xnor3_2.spice
* Created: Wed Sep  2 11:30:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ls__xnor3_2.pex.spice"
.subckt sky130_fd_sc_ls__xnor3_2  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_83_247#_M1009_g N_A_27_373#_M1009_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1152 AS=0.1824 PD=1 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1007 N_A_83_247#_M1007_d N_A_M1007_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.64
+ AD=0.12 AS=0.1152 PD=1.015 PS=1 NRD=0 NRS=14.988 M=1 R=4.26667 SA=75000.7
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1018 N_A_329_81#_M1018_d N_B_M1018_g N_A_83_247#_M1007_d VNB NSHORT L=0.15
+ W=0.64 AD=0.144664 AS=0.12 PD=1.44906 PS=1.015 NRD=0 NRS=17.808 M=1 R=4.26667
+ SA=75001.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1002 N_A_27_373#_M1002_d N_A_397_21#_M1002_g N_A_329_81#_M1018_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0817019 AS=0.0949358 PD=0.792453 PS=0.950943 NRD=0
+ NRS=48.864 M=1 R=2.8 SA=75000.9 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1001 N_A_332_373#_M1001_d N_B_M1001_g N_A_27_373#_M1002_d VNB NSHORT L=0.15
+ W=0.64 AD=0.112 AS=0.124498 PD=0.99 PS=1.20755 NRD=2.808 NRS=14.988 M=1
+ R=4.26667 SA=75001 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1000 N_A_83_247#_M1000_d N_A_397_21#_M1000_g N_A_332_373#_M1001_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.3525 AS=0.112 PD=2.83 PS=0.99 NRD=92.952 NRS=10.308 M=1
+ R=4.26667 SA=75001.5 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1014 N_VGND_M1014_d N_B_M1014_g N_A_397_21#_M1014_s VNB NSHORT L=0.15 W=0.74
+ AD=0.3368 AS=0.2109 PD=2.67 PS=2.05 NRD=64.884 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1023 N_A_1057_74#_M1023_d N_A_1027_48#_M1023_g N_A_329_81#_M1023_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1019 N_A_332_373#_M1019_d N_C_M1019_g N_A_1057_74#_M1023_d VNB NSHORT L=0.15
+ W=0.64 AD=0.2272 AS=0.112 PD=1.99 PS=0.99 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1010 N_VGND_M1010_d N_C_M1010_g N_A_1027_48#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.276711 AS=0.1197 PD=1.33603 PS=1.41 NRD=172.524 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_1057_74#_M1006_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.487539 PD=1.02 PS=2.35397 NRD=0 NRS=17.016 M=1 R=4.93333
+ SA=75000.9 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1015 N_X_M1006_d N_A_1057_74#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_A_83_247#_M1008_g N_A_27_373#_M1008_s VPB PHIGHVT L=0.15
+ W=1 AD=0.195 AS=0.295 PD=1.39 PS=2.59 NRD=4.9053 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1011 N_A_83_247#_M1011_d N_A_M1011_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.202826 AS=0.195 PD=1.51087 PS=1.39 NRD=3.9203 NRS=16.7253 M=1 R=6.66667
+ SA=75000.8 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1005 N_A_332_373#_M1005_d N_B_M1005_g N_A_83_247#_M1011_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.197741 AS=0.170374 PD=1.47568 PS=1.26913 NRD=39.8531 NRS=21.6897
+ M=1 R=5.6 SA=75001.3 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1004 N_A_27_373#_M1004_d N_A_397_21#_M1004_g N_A_332_373#_M1005_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1024 AS=0.150659 PD=0.96 PS=1.12432 NRD=9.2196 NRS=3.0732
+ M=1 R=4.26667 SA=75001.9 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1003 N_A_329_81#_M1003_d N_B_M1003_g N_A_27_373#_M1004_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.133449 AS=0.1024 PD=1.06378 PS=0.96 NRD=31.5397 NRS=3.0732 M=1
+ R=4.26667 SA=75002.4 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1012 N_A_83_247#_M1012_d N_A_397_21#_M1012_g N_A_329_81#_M1003_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.3766 AS=0.175151 PD=2.89 PS=1.39622 NRD=92.2354 NRS=2.3443
+ M=1 R=5.6 SA=75002.3 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1020 N_VPWR_M1020_d N_B_M1020_g N_A_397_21#_M1020_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.4382 AS=0.3248 PD=3.15 PS=2.82 NRD=16.7056 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.3 A=0.168 P=2.54 MULT=1
MM1021 N_A_1057_74#_M1021_d N_A_1027_48#_M1021_g N_A_332_373#_M1021_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.213825 AS=0.2436 PD=1.435 PS=2.26 NRD=22.261
+ NRS=2.3443 M=1 R=5.6 SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1016 N_A_329_81#_M1016_d N_C_M1016_g N_A_1057_74#_M1021_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2436 AS=0.213825 PD=2.26 PS=1.435 NRD=2.3443 NRS=23.443 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1017 N_VPWR_M1017_d N_C_M1017_g N_A_1027_48#_M1017_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.174836 AS=0.1856 PD=1.2 PS=1.86 NRD=75.4116 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1013 N_X_M1013_d N_A_1057_74#_M1013_g N_VPWR_M1017_d VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.305964 PD=1.42 PS=2.1 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1022 N_X_M1013_d N_A_1057_74#_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1.12
+ AD=0.168 AS=0.3248 PD=1.42 PS=2.82 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX24_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_ls__xnor3_2.pxi.spice"
*
.ends
*
*
