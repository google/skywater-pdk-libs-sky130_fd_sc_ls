* File: sky130_fd_sc_ls__dfxtp_1.pxi.spice
* Created: Wed Sep  2 11:02:18 2020
* 
x_PM_SKY130_FD_SC_LS__DFXTP_1%CLK N_CLK_M1022_g N_CLK_c_183_n N_CLK_M1014_g CLK
+ N_CLK_c_184_n PM_SKY130_FD_SC_LS__DFXTP_1%CLK
x_PM_SKY130_FD_SC_LS__DFXTP_1%A_27_74# N_A_27_74#_M1022_s N_A_27_74#_M1014_s
+ N_A_27_74#_c_215_n N_A_27_74#_M1015_g N_A_27_74#_c_216_n N_A_27_74#_M1001_g
+ N_A_27_74#_M1017_g N_A_27_74#_c_240_n N_A_27_74#_c_241_n N_A_27_74#_M1013_g
+ N_A_27_74#_c_242_n N_A_27_74#_M1019_g N_A_27_74#_c_243_n N_A_27_74#_M1023_g
+ N_A_27_74#_c_245_n N_A_27_74#_c_219_n N_A_27_74#_c_246_n N_A_27_74#_c_247_n
+ N_A_27_74#_c_220_n N_A_27_74#_c_221_n N_A_27_74#_c_265_n N_A_27_74#_c_222_n
+ N_A_27_74#_c_223_n N_A_27_74#_c_224_n N_A_27_74#_c_225_n N_A_27_74#_c_226_n
+ N_A_27_74#_c_227_n N_A_27_74#_c_228_n N_A_27_74#_c_229_n N_A_27_74#_c_230_n
+ N_A_27_74#_c_249_n N_A_27_74#_c_250_n N_A_27_74#_c_231_n N_A_27_74#_c_232_n
+ N_A_27_74#_c_347_p N_A_27_74#_c_300_p N_A_27_74#_c_233_n N_A_27_74#_c_234_n
+ N_A_27_74#_c_272_n N_A_27_74#_c_298_p N_A_27_74#_c_235_n N_A_27_74#_c_236_n
+ N_A_27_74#_c_237_n PM_SKY130_FD_SC_LS__DFXTP_1%A_27_74#
x_PM_SKY130_FD_SC_LS__DFXTP_1%D N_D_c_496_n N_D_M1012_g N_D_c_493_n N_D_M1006_g
+ D N_D_c_494_n N_D_c_495_n D PM_SKY130_FD_SC_LS__DFXTP_1%D
x_PM_SKY130_FD_SC_LS__DFXTP_1%A_206_368# N_A_206_368#_M1001_d
+ N_A_206_368#_M1015_d N_A_206_368#_c_540_n N_A_206_368#_c_541_n
+ N_A_206_368#_c_553_n N_A_206_368#_c_554_n N_A_206_368#_c_555_n
+ N_A_206_368#_M1021_g N_A_206_368#_M1016_g N_A_206_368#_c_543_n
+ N_A_206_368#_M1005_g N_A_206_368#_c_556_n N_A_206_368#_M1002_g
+ N_A_206_368#_c_557_n N_A_206_368#_c_544_n N_A_206_368#_c_558_n
+ N_A_206_368#_c_559_n N_A_206_368#_c_606_n N_A_206_368#_c_545_n
+ N_A_206_368#_c_546_n N_A_206_368#_c_547_n N_A_206_368#_c_561_n
+ N_A_206_368#_c_562_n N_A_206_368#_c_563_n N_A_206_368#_c_564_n
+ N_A_206_368#_c_548_n N_A_206_368#_c_549_n N_A_206_368#_c_567_n
+ N_A_206_368#_c_568_n N_A_206_368#_c_569_n N_A_206_368#_c_550_n
+ N_A_206_368#_c_551_n N_A_206_368#_c_552_n
+ PM_SKY130_FD_SC_LS__DFXTP_1%A_206_368#
x_PM_SKY130_FD_SC_LS__DFXTP_1%A_713_458# N_A_713_458#_M1004_d
+ N_A_713_458#_M1018_d N_A_713_458#_M1000_g N_A_713_458#_M1011_g
+ N_A_713_458#_c_776_n N_A_713_458#_c_784_n N_A_713_458#_c_777_n
+ N_A_713_458#_c_778_n N_A_713_458#_c_803_n N_A_713_458#_c_779_n
+ N_A_713_458#_c_824_n N_A_713_458#_c_780_n N_A_713_458#_c_781_n
+ N_A_713_458#_c_782_n PM_SKY130_FD_SC_LS__DFXTP_1%A_713_458#
x_PM_SKY130_FD_SC_LS__DFXTP_1%A_561_463# N_A_561_463#_M1017_d
+ N_A_561_463#_M1021_d N_A_561_463#_c_880_n N_A_561_463#_M1018_g
+ N_A_561_463#_c_871_n N_A_561_463#_M1004_g N_A_561_463#_c_873_n
+ N_A_561_463#_c_874_n N_A_561_463#_c_875_n N_A_561_463#_c_876_n
+ N_A_561_463#_c_882_n N_A_561_463#_c_877_n N_A_561_463#_c_883_n
+ N_A_561_463#_c_884_n N_A_561_463#_c_878_n N_A_561_463#_c_879_n
+ PM_SKY130_FD_SC_LS__DFXTP_1%A_561_463#
x_PM_SKY130_FD_SC_LS__DFXTP_1%A_1210_314# N_A_1210_314#_M1007_s
+ N_A_1210_314#_M1008_s N_A_1210_314#_c_1001_n N_A_1210_314#_M1003_g
+ N_A_1210_314#_M1020_g N_A_1210_314#_c_992_n N_A_1210_314#_M1010_g
+ N_A_1210_314#_M1009_g N_A_1210_314#_c_1003_n N_A_1210_314#_c_1004_n
+ N_A_1210_314#_c_1005_n N_A_1210_314#_c_994_n N_A_1210_314#_c_1006_n
+ N_A_1210_314#_c_995_n N_A_1210_314#_c_996_n N_A_1210_314#_c_997_n
+ N_A_1210_314#_c_998_n N_A_1210_314#_c_1009_n N_A_1210_314#_c_999_n
+ N_A_1210_314#_c_1000_n PM_SKY130_FD_SC_LS__DFXTP_1%A_1210_314#
x_PM_SKY130_FD_SC_LS__DFXTP_1%A_1011_424# N_A_1011_424#_M1005_d
+ N_A_1011_424#_M1019_d N_A_1011_424#_c_1107_n N_A_1011_424#_c_1108_n
+ N_A_1011_424#_c_1116_n N_A_1011_424#_M1008_g N_A_1011_424#_M1007_g
+ N_A_1011_424#_c_1117_n N_A_1011_424#_c_1123_n N_A_1011_424#_c_1118_n
+ N_A_1011_424#_c_1119_n N_A_1011_424#_c_1110_n N_A_1011_424#_c_1111_n
+ N_A_1011_424#_c_1112_n N_A_1011_424#_c_1113_n N_A_1011_424#_c_1114_n
+ PM_SKY130_FD_SC_LS__DFXTP_1%A_1011_424#
x_PM_SKY130_FD_SC_LS__DFXTP_1%VPWR N_VPWR_M1014_d N_VPWR_M1012_s N_VPWR_M1000_d
+ N_VPWR_M1003_d N_VPWR_M1008_d N_VPWR_c_1210_n N_VPWR_c_1211_n N_VPWR_c_1212_n
+ N_VPWR_c_1213_n N_VPWR_c_1214_n VPWR N_VPWR_c_1215_n N_VPWR_c_1216_n
+ N_VPWR_c_1217_n N_VPWR_c_1218_n N_VPWR_c_1209_n N_VPWR_c_1220_n
+ N_VPWR_c_1221_n N_VPWR_c_1222_n N_VPWR_c_1223_n
+ PM_SKY130_FD_SC_LS__DFXTP_1%VPWR
x_PM_SKY130_FD_SC_LS__DFXTP_1%A_454_503# N_A_454_503#_M1006_d
+ N_A_454_503#_M1012_d N_A_454_503#_c_1308_n N_A_454_503#_c_1309_n
+ N_A_454_503#_c_1310_n PM_SKY130_FD_SC_LS__DFXTP_1%A_454_503#
x_PM_SKY130_FD_SC_LS__DFXTP_1%Q N_Q_M1009_d N_Q_M1010_d N_Q_c_1346_n
+ N_Q_c_1347_n N_Q_c_1343_n Q Q Q PM_SKY130_FD_SC_LS__DFXTP_1%Q
x_PM_SKY130_FD_SC_LS__DFXTP_1%VGND N_VGND_M1022_d N_VGND_M1006_s N_VGND_M1011_d
+ N_VGND_M1020_d N_VGND_M1007_d N_VGND_c_1369_n N_VGND_c_1370_n N_VGND_c_1371_n
+ N_VGND_c_1372_n N_VGND_c_1373_n N_VGND_c_1374_n N_VGND_c_1375_n VGND
+ N_VGND_c_1376_n N_VGND_c_1377_n N_VGND_c_1378_n N_VGND_c_1379_n
+ N_VGND_c_1380_n N_VGND_c_1381_n N_VGND_c_1382_n N_VGND_c_1383_n
+ N_VGND_c_1384_n N_VGND_c_1385_n PM_SKY130_FD_SC_LS__DFXTP_1%VGND
cc_1 VNB N_CLK_M1022_g 0.0305265f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_CLK_c_183_n 0.0463134f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_CLK_c_184_n 0.0163904f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_4 VNB N_A_27_74#_c_215_n 0.0427448f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_5 VNB N_A_27_74#_c_216_n 0.0185203f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.465
cc_6 VNB N_A_27_74#_M1017_g 0.0495777f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.665
cc_7 VNB N_A_27_74#_M1023_g 0.0374125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_219_n 0.0247745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_220_n 0.00335275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_221_n 0.00891132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_222_n 0.00152612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_223_n 0.00741633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_224_n 0.00134302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_225_n 0.00296184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_226_n 0.0079485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_227_n 0.00222565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_228_n 0.00300069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_229_n 0.0239223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_230_n 0.00245548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_231_n 4.22754e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_232_n 0.00684074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_233_n 0.00151705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_74#_c_234_n 0.00509724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_235_n 0.00404212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_236_n 0.0462362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_74#_c_237_n 0.0130783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_D_c_493_n 0.0184239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_D_c_494_n 0.0469166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_D_c_495_n 0.00642682f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.665
cc_30 VNB N_A_206_368#_c_540_n 0.13302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_206_368#_c_541_n 0.0124288f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.465
cc_32 VNB N_A_206_368#_M1016_g 0.0271992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_206_368#_c_543_n 0.0181774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_206_368#_c_544_n 0.00421781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_206_368#_c_545_n 0.00479134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_206_368#_c_546_n 0.00437351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_206_368#_c_547_n 0.0030093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_206_368#_c_548_n 0.00444634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_206_368#_c_549_n 0.0279774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_206_368#_c_550_n 0.0053436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_206_368#_c_551_n 0.0393248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_206_368#_c_552_n 0.0655348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_713_458#_M1011_g 0.0212764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_713_458#_c_776_n 0.0155751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_713_458#_c_777_n 0.00387496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_713_458#_c_778_n 0.00790294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_713_458#_c_779_n 0.00580454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_713_458#_c_780_n 0.0040861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_713_458#_c_781_n 9.8498e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_713_458#_c_782_n 0.0574805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_561_463#_c_871_n 0.011518f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_52 VNB N_A_561_463#_M1004_g 0.0345542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_561_463#_c_873_n 0.0125006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_561_463#_c_874_n 0.00148109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_561_463#_c_875_n 0.00864345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_561_463#_c_876_n 0.00334202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_561_463#_c_877_n 0.00360489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_561_463#_c_878_n 0.00203572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_561_463#_c_879_n 0.0138802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1210_314#_M1020_g 0.0472681f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_61 VNB N_A_1210_314#_c_992_n 0.0263455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1210_314#_M1009_g 0.0310216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1210_314#_c_994_n 0.00711261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1210_314#_c_995_n 0.00176879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1210_314#_c_996_n 0.00372926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1210_314#_c_997_n 0.00374187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1210_314#_c_998_n 0.0113192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1210_314#_c_999_n 0.0042334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1210_314#_c_1000_n 0.00376244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1011_424#_c_1107_n 0.0365784f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_71 VNB N_A_1011_424#_c_1108_n 0.0100925f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_72 VNB N_A_1011_424#_M1007_g 0.0321248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1011_424#_c_1110_n 0.00173344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1011_424#_c_1111_n 0.00513905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1011_424#_c_1112_n 0.00104376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1011_424#_c_1113_n 0.00243913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1011_424#_c_1114_n 0.0360822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VPWR_c_1209_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_454_503#_c_1308_n 0.00650149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_454_503#_c_1309_n 6.56034e-19 $X=-0.19 $Y=-0.245 $X2=0.34
+ $Y2=1.465
cc_81 VNB N_A_454_503#_c_1310_n 0.00163418f $X=-0.19 $Y=-0.245 $X2=0.315
+ $Y2=1.465
cc_82 VNB N_Q_c_1343_n 0.0247211f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.665
cc_83 VNB Q 0.0265914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB Q 0.0126022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1369_n 0.00530967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1370_n 0.00615071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1371_n 0.00712015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1372_n 0.0199091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1373_n 0.00575282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1374_n 0.0464757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1375_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1376_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1377_n 0.0278703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1378_n 0.0413632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1379_n 0.0188435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1380_n 0.0192354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1381_n 0.443225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1382_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1383_n 0.0043669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1384_n 0.00477982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1385_n 0.00586939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VPB N_CLK_c_183_n 0.0289619f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_103 VPB N_CLK_c_184_n 0.0073823f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_104 VPB N_A_27_74#_c_215_n 0.0252403f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_105 VPB N_A_27_74#_M1017_g 0.00503294f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=1.665
cc_106 VPB N_A_27_74#_c_240_n 0.0149453f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_27_74#_c_241_n 0.0226066f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_27_74#_c_242_n 0.0165272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_27_74#_c_243_n 0.0458434f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_27_74#_M1023_g 0.00176303f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_27_74#_c_245_n 0.0236601f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_27_74#_c_246_n 0.00758177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_27_74#_c_247_n 0.035396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_27_74#_c_222_n 0.0030872f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_74#_c_249_n 0.00894186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_27_74#_c_250_n 0.0324191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_27_74#_c_232_n 0.00101285f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_D_c_496_n 0.069304f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_119 VPB N_D_c_495_n 0.00456891f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=1.665
cc_120 VPB D 0.00365325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_206_368#_c_553_n 0.0688733f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_122 VPB N_A_206_368#_c_554_n 0.0173431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_206_368#_c_555_n 0.0214269f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=1.665
cc_124 VPB N_A_206_368#_c_556_n 0.0612378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_206_368#_c_557_n 0.0222625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_206_368#_c_558_n 0.00608915f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_206_368#_c_559_n 0.011479f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_206_368#_c_545_n 0.00408019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_206_368#_c_561_n 0.00590845f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_206_368#_c_562_n 0.00379772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_206_368#_c_563_n 0.00973344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_206_368#_c_564_n 0.00160725f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_206_368#_c_548_n 5.28092e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_206_368#_c_549_n 0.0248155f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_206_368#_c_567_n 0.00133504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_206_368#_c_568_n 0.00131318f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_206_368#_c_569_n 0.0022225f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_713_458#_c_776_n 0.029545f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_713_458#_c_784_n 0.0257248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_713_458#_c_780_n 0.00489235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_561_463#_c_880_n 0.0188172f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_142 VPB N_A_561_463#_c_874_n 0.00525969f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_561_463#_c_882_n 0.0136116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_561_463#_c_883_n 0.00234446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_561_463#_c_884_n 0.00559867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_561_463#_c_878_n 7.67418e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_561_463#_c_879_n 0.0500183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_1210_314#_c_1001_n 0.0191465f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_149 VPB N_A_1210_314#_c_992_n 0.031255f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_1210_314#_c_1003_n 0.0668874f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_1210_314#_c_1004_n 0.0158383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_1210_314#_c_1005_n 0.01231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_1210_314#_c_1006_n 0.00261305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_1210_314#_c_997_n 0.00361628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_1210_314#_c_998_n 0.00515132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_1210_314#_c_1009_n 0.00279611f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_1210_314#_c_999_n 0.00129348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_1011_424#_c_1108_n 9.33079e-19 $X=-0.19 $Y=1.66 $X2=0.155
+ $Y2=1.58
cc_159 VPB N_A_1011_424#_c_1116_n 0.0227322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_1011_424#_c_1117_n 0.00823029f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_1011_424#_c_1118_n 0.00757102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_1011_424#_c_1119_n 2.36604e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_1011_424#_c_1111_n 0.00103061f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_1210_n 0.00799246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_1211_n 0.0229599f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1212_n 0.0186927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_1213_n 0.0518589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1214_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_1215_n 0.0203276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1216_n 0.0469022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1217_n 0.0204602f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1218_n 0.0190763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1209_n 0.11565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1220_n 0.0233502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1221_n 0.0152649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1222_n 0.0145986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1223_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_454_503#_c_1308_n 0.00839922f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_Q_c_1346_n 0.0333962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_Q_c_1347_n 0.00710642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_Q_c_1343_n 0.0154743f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=1.665
cc_182 N_CLK_M1022_g N_A_27_74#_c_215_n 0.0040435f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_183 N_CLK_c_183_n N_A_27_74#_c_215_n 0.0455528f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_184 N_CLK_c_184_n N_A_27_74#_c_215_n 2.10791e-19 $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_185 N_CLK_M1022_g N_A_27_74#_c_216_n 0.0163593f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_186 N_CLK_M1022_g N_A_27_74#_c_219_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_187 N_CLK_c_183_n N_A_27_74#_c_246_n 0.0016558f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_188 N_CLK_c_184_n N_A_27_74#_c_246_n 0.0258609f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_189 N_CLK_c_183_n N_A_27_74#_c_247_n 0.0104891f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_190 N_CLK_M1022_g N_A_27_74#_c_220_n 0.0143116f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_191 N_CLK_c_183_n N_A_27_74#_c_220_n 0.00138858f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_192 N_CLK_c_184_n N_A_27_74#_c_220_n 0.010454f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_193 N_CLK_c_183_n N_A_27_74#_c_221_n 0.0015038f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_194 N_CLK_c_184_n N_A_27_74#_c_221_n 0.0209983f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_195 N_CLK_c_183_n N_A_27_74#_c_265_n 0.0139121f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_196 N_CLK_c_184_n N_A_27_74#_c_265_n 0.00433199f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_197 N_CLK_c_183_n N_A_27_74#_c_222_n 0.00397589f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_198 N_CLK_M1022_g N_A_27_74#_c_224_n 4.27363e-19 $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_199 N_CLK_M1022_g N_A_27_74#_c_234_n 0.00515282f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_200 N_CLK_c_183_n N_A_27_74#_c_234_n 0.00330504f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_201 N_CLK_c_184_n N_A_27_74#_c_234_n 0.0379192f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_202 N_CLK_M1022_g N_A_27_74#_c_272_n 0.0018749f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_203 N_CLK_c_183_n N_A_206_368#_c_557_n 5.38656e-19 $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_204 N_CLK_c_183_n N_VPWR_c_1210_n 0.00486623f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_205 N_CLK_c_183_n N_VPWR_c_1209_n 0.00861168f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_206 N_CLK_c_183_n N_VPWR_c_1220_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_207 N_CLK_M1022_g N_VGND_c_1369_n 0.0122115f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_208 N_CLK_M1022_g N_VGND_c_1376_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_209 N_CLK_M1022_g N_VGND_c_1381_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A_27_74#_M1017_g N_D_c_493_n 0.0147551f $X=3.105 $Y=0.835 $X2=0 $Y2=0
cc_211 N_A_27_74#_c_225_n N_D_c_493_n 0.00129456f $X=1.73 $Y=0.73 $X2=0 $Y2=0
cc_212 N_A_27_74#_c_226_n N_D_c_493_n 0.0131377f $X=2.485 $Y=0.815 $X2=0 $Y2=0
cc_213 N_A_27_74#_c_228_n N_D_c_493_n 0.00837729f $X=2.57 $Y=0.73 $X2=0 $Y2=0
cc_214 N_A_27_74#_c_226_n N_D_c_494_n 0.00498006f $X=2.485 $Y=0.815 $X2=0 $Y2=0
cc_215 N_A_27_74#_c_226_n N_D_c_495_n 0.0176307f $X=2.485 $Y=0.815 $X2=0 $Y2=0
cc_216 N_A_27_74#_c_223_n N_A_206_368#_M1001_d 0.00654387f $X=1.645 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_217 N_A_27_74#_M1017_g N_A_206_368#_c_540_n 0.00736788f $X=3.105 $Y=0.835
+ $X2=0 $Y2=0
cc_218 N_A_27_74#_c_223_n N_A_206_368#_c_540_n 4.6256e-19 $X=1.645 $Y=0.34 $X2=0
+ $Y2=0
cc_219 N_A_27_74#_c_226_n N_A_206_368#_c_540_n 0.00369117f $X=2.485 $Y=0.815
+ $X2=0 $Y2=0
cc_220 N_A_27_74#_c_229_n N_A_206_368#_c_540_n 0.015252f $X=3.59 $Y=0.36 $X2=0
+ $Y2=0
cc_221 N_A_27_74#_c_230_n N_A_206_368#_c_540_n 0.0035717f $X=2.655 $Y=0.36 $X2=0
+ $Y2=0
cc_222 N_A_27_74#_c_216_n N_A_206_368#_c_541_n 0.0119162f $X=1.115 $Y=1.22 $X2=0
+ $Y2=0
cc_223 N_A_27_74#_c_223_n N_A_206_368#_c_541_n 9.85082e-19 $X=1.645 $Y=0.34
+ $X2=0 $Y2=0
cc_224 N_A_27_74#_M1017_g N_A_206_368#_c_553_n 0.0127641f $X=3.105 $Y=0.835
+ $X2=0 $Y2=0
cc_225 N_A_27_74#_c_249_n N_A_206_368#_c_553_n 2.94693e-19 $X=3.59 $Y=1.915
+ $X2=0 $Y2=0
cc_226 N_A_27_74#_c_240_n N_A_206_368#_c_554_n 0.00479623f $X=3.265 $Y=2.35
+ $X2=0 $Y2=0
cc_227 N_A_27_74#_c_250_n N_A_206_368#_c_554_n 0.0127641f $X=3.235 $Y=1.915
+ $X2=0 $Y2=0
cc_228 N_A_27_74#_c_240_n N_A_206_368#_c_555_n 0.0041237f $X=3.265 $Y=2.35 $X2=0
+ $Y2=0
cc_229 N_A_27_74#_c_241_n N_A_206_368#_c_555_n 0.00926866f $X=3.265 $Y=2.44
+ $X2=0 $Y2=0
cc_230 N_A_27_74#_M1017_g N_A_206_368#_M1016_g 0.00749916f $X=3.105 $Y=0.835
+ $X2=0 $Y2=0
cc_231 N_A_27_74#_c_229_n N_A_206_368#_M1016_g 0.0133538f $X=3.59 $Y=0.36 $X2=0
+ $Y2=0
cc_232 N_A_27_74#_c_249_n N_A_206_368#_M1016_g 0.0021868f $X=3.59 $Y=1.915 $X2=0
+ $Y2=0
cc_233 N_A_27_74#_c_231_n N_A_206_368#_M1016_g 0.00667594f $X=3.675 $Y=0.69
+ $X2=0 $Y2=0
cc_234 N_A_27_74#_c_232_n N_A_206_368#_M1016_g 0.00426708f $X=3.675 $Y=1.75
+ $X2=0 $Y2=0
cc_235 N_A_27_74#_c_298_p N_A_206_368#_M1016_g 0.00373495f $X=3.675 $Y=0.775
+ $X2=0 $Y2=0
cc_236 N_A_27_74#_M1023_g N_A_206_368#_c_543_n 0.0139309f $X=5.765 $Y=0.83 $X2=0
+ $Y2=0
cc_237 N_A_27_74#_c_300_p N_A_206_368#_c_543_n 9.72585e-19 $X=4.575 $Y=0.69
+ $X2=0 $Y2=0
cc_238 N_A_27_74#_c_235_n N_A_206_368#_c_543_n 4.97101e-19 $X=5.73 $Y=0.345
+ $X2=0 $Y2=0
cc_239 N_A_27_74#_c_236_n N_A_206_368#_c_543_n 0.00468991f $X=5.73 $Y=0.345
+ $X2=0 $Y2=0
cc_240 N_A_27_74#_c_237_n N_A_206_368#_c_543_n 0.0118082f $X=5.565 $Y=0.382
+ $X2=0 $Y2=0
cc_241 N_A_27_74#_c_242_n N_A_206_368#_c_556_n 0.0221559f $X=4.98 $Y=2.045 $X2=0
+ $Y2=0
cc_242 N_A_27_74#_c_243_n N_A_206_368#_c_556_n 0.0270049f $X=5.69 $Y=1.765 $X2=0
+ $Y2=0
cc_243 N_A_27_74#_c_215_n N_A_206_368#_c_557_n 0.0121876f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_244 N_A_27_74#_c_247_n N_A_206_368#_c_557_n 0.00481788f $X=0.28 $Y=2.815
+ $X2=0 $Y2=0
cc_245 N_A_27_74#_c_216_n N_A_206_368#_c_544_n 0.0060011f $X=1.115 $Y=1.22 $X2=0
+ $Y2=0
cc_246 N_A_27_74#_c_223_n N_A_206_368#_c_544_n 0.012787f $X=1.645 $Y=0.34 $X2=0
+ $Y2=0
cc_247 N_A_27_74#_c_225_n N_A_206_368#_c_544_n 0.00944376f $X=1.73 $Y=0.73 $X2=0
+ $Y2=0
cc_248 N_A_27_74#_c_227_n N_A_206_368#_c_544_n 0.0133618f $X=1.815 $Y=0.815
+ $X2=0 $Y2=0
cc_249 N_A_27_74#_c_272_n N_A_206_368#_c_544_n 0.0554258f $X=0.905 $Y=0.96 $X2=0
+ $Y2=0
cc_250 N_A_27_74#_c_241_n N_A_206_368#_c_559_n 0.00849081f $X=3.265 $Y=2.44
+ $X2=0 $Y2=0
cc_251 N_A_27_74#_c_242_n N_A_206_368#_c_606_n 3.68762e-19 $X=4.98 $Y=2.045
+ $X2=0 $Y2=0
cc_252 N_A_27_74#_c_242_n N_A_206_368#_c_545_n 0.0134889f $X=4.98 $Y=2.045 $X2=0
+ $Y2=0
cc_253 N_A_27_74#_c_245_n N_A_206_368#_c_545_n 0.0113102f $X=4.98 $Y=1.765 $X2=0
+ $Y2=0
cc_254 N_A_27_74#_c_245_n N_A_206_368#_c_546_n 0.00601497f $X=4.98 $Y=1.765
+ $X2=0 $Y2=0
cc_255 N_A_27_74#_c_242_n N_A_206_368#_c_561_n 0.00985245f $X=4.98 $Y=2.045
+ $X2=0 $Y2=0
cc_256 N_A_27_74#_c_242_n N_A_206_368#_c_562_n 7.86426e-19 $X=4.98 $Y=2.045
+ $X2=0 $Y2=0
cc_257 N_A_27_74#_c_243_n N_A_206_368#_c_562_n 4.51027e-19 $X=5.69 $Y=1.765
+ $X2=0 $Y2=0
cc_258 N_A_27_74#_c_215_n N_A_206_368#_c_563_n 0.00641904f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_259 N_A_27_74#_c_222_n N_A_206_368#_c_563_n 0.00584697f $X=0.76 $Y=1.95 $X2=0
+ $Y2=0
cc_260 N_A_27_74#_c_234_n N_A_206_368#_c_563_n 0.00736457f $X=0.905 $Y=1.045
+ $X2=0 $Y2=0
cc_261 N_A_27_74#_c_215_n N_A_206_368#_c_564_n 0.00120435f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_262 N_A_27_74#_c_222_n N_A_206_368#_c_564_n 0.0052471f $X=0.76 $Y=1.95 $X2=0
+ $Y2=0
cc_263 N_A_27_74#_c_215_n N_A_206_368#_c_548_n 0.00263834f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_264 N_A_27_74#_c_222_n N_A_206_368#_c_548_n 0.00523409f $X=0.76 $Y=1.95 $X2=0
+ $Y2=0
cc_265 N_A_27_74#_c_227_n N_A_206_368#_c_548_n 0.00414227f $X=1.815 $Y=0.815
+ $X2=0 $Y2=0
cc_266 N_A_27_74#_c_234_n N_A_206_368#_c_548_n 0.016628f $X=0.905 $Y=1.045 $X2=0
+ $Y2=0
cc_267 N_A_27_74#_c_215_n N_A_206_368#_c_549_n 0.0176835f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_268 N_A_27_74#_c_241_n N_A_206_368#_c_568_n 0.00789803f $X=3.265 $Y=2.44
+ $X2=0 $Y2=0
cc_269 N_A_27_74#_c_242_n N_A_206_368#_c_569_n 0.0113526f $X=4.98 $Y=2.045 $X2=0
+ $Y2=0
cc_270 N_A_27_74#_c_243_n N_A_206_368#_c_550_n 0.00167373f $X=5.69 $Y=1.765
+ $X2=0 $Y2=0
cc_271 N_A_27_74#_M1023_g N_A_206_368#_c_550_n 7.90155e-19 $X=5.765 $Y=0.83
+ $X2=0 $Y2=0
cc_272 N_A_27_74#_M1023_g N_A_206_368#_c_551_n 0.020918f $X=5.765 $Y=0.83 $X2=0
+ $Y2=0
cc_273 N_A_27_74#_c_245_n N_A_206_368#_c_551_n 0.0251563f $X=4.98 $Y=1.765 $X2=0
+ $Y2=0
cc_274 N_A_27_74#_c_215_n N_A_206_368#_c_552_n 0.0119162f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_275 N_A_27_74#_c_223_n N_A_206_368#_c_552_n 0.00806761f $X=1.645 $Y=0.34
+ $X2=0 $Y2=0
cc_276 N_A_27_74#_c_225_n N_A_206_368#_c_552_n 0.00952884f $X=1.73 $Y=0.73 $X2=0
+ $Y2=0
cc_277 N_A_27_74#_c_227_n N_A_206_368#_c_552_n 0.00894445f $X=1.815 $Y=0.815
+ $X2=0 $Y2=0
cc_278 N_A_27_74#_c_272_n N_A_206_368#_c_552_n 7.55802e-19 $X=0.905 $Y=0.96
+ $X2=0 $Y2=0
cc_279 N_A_27_74#_c_237_n N_A_713_458#_M1004_d 0.00277152f $X=5.565 $Y=0.382
+ $X2=-0.19 $Y2=-0.245
cc_280 N_A_27_74#_M1017_g N_A_713_458#_M1011_g 0.00207737f $X=3.105 $Y=0.835
+ $X2=0 $Y2=0
cc_281 N_A_27_74#_c_229_n N_A_713_458#_M1011_g 6.23789e-19 $X=3.59 $Y=0.36 $X2=0
+ $Y2=0
cc_282 N_A_27_74#_c_231_n N_A_713_458#_M1011_g 0.00418052f $X=3.675 $Y=0.69
+ $X2=0 $Y2=0
cc_283 N_A_27_74#_c_232_n N_A_713_458#_M1011_g 0.00631548f $X=3.675 $Y=1.75
+ $X2=0 $Y2=0
cc_284 N_A_27_74#_c_347_p N_A_713_458#_M1011_g 0.0141002f $X=4.49 $Y=0.775 $X2=0
+ $Y2=0
cc_285 N_A_27_74#_c_240_n N_A_713_458#_c_776_n 0.0105386f $X=3.265 $Y=2.35 $X2=0
+ $Y2=0
cc_286 N_A_27_74#_c_249_n N_A_713_458#_c_776_n 0.0102386f $X=3.59 $Y=1.915 $X2=0
+ $Y2=0
cc_287 N_A_27_74#_c_250_n N_A_713_458#_c_776_n 0.0213493f $X=3.235 $Y=1.915
+ $X2=0 $Y2=0
cc_288 N_A_27_74#_c_232_n N_A_713_458#_c_776_n 0.0151009f $X=3.675 $Y=1.75 $X2=0
+ $Y2=0
cc_289 N_A_27_74#_c_240_n N_A_713_458#_c_784_n 0.00964421f $X=3.265 $Y=2.35
+ $X2=0 $Y2=0
cc_290 N_A_27_74#_c_241_n N_A_713_458#_c_784_n 0.0330974f $X=3.265 $Y=2.44 $X2=0
+ $Y2=0
cc_291 N_A_27_74#_c_249_n N_A_713_458#_c_784_n 3.22945e-19 $X=3.59 $Y=1.915
+ $X2=0 $Y2=0
cc_292 N_A_27_74#_c_347_p N_A_713_458#_c_777_n 0.0132764f $X=4.49 $Y=0.775 $X2=0
+ $Y2=0
cc_293 N_A_27_74#_c_245_n N_A_713_458#_c_778_n 3.29975e-19 $X=4.98 $Y=1.765
+ $X2=0 $Y2=0
cc_294 N_A_27_74#_c_347_p N_A_713_458#_c_778_n 0.00373759f $X=4.49 $Y=0.775
+ $X2=0 $Y2=0
cc_295 N_A_27_74#_c_237_n N_A_713_458#_c_778_n 0.00391108f $X=5.565 $Y=0.382
+ $X2=0 $Y2=0
cc_296 N_A_27_74#_c_347_p N_A_713_458#_c_803_n 0.0133618f $X=4.49 $Y=0.775 $X2=0
+ $Y2=0
cc_297 N_A_27_74#_c_300_p N_A_713_458#_c_803_n 0.00663557f $X=4.575 $Y=0.69
+ $X2=0 $Y2=0
cc_298 N_A_27_74#_c_237_n N_A_713_458#_c_803_n 0.0127055f $X=5.565 $Y=0.382
+ $X2=0 $Y2=0
cc_299 N_A_27_74#_c_232_n N_A_713_458#_c_779_n 0.0283347f $X=3.675 $Y=1.75 $X2=0
+ $Y2=0
cc_300 N_A_27_74#_c_347_p N_A_713_458#_c_779_n 0.0233764f $X=4.49 $Y=0.775 $X2=0
+ $Y2=0
cc_301 N_A_27_74#_c_242_n N_A_713_458#_c_780_n 0.00123273f $X=4.98 $Y=2.045
+ $X2=0 $Y2=0
cc_302 N_A_27_74#_c_245_n N_A_713_458#_c_780_n 8.61424e-19 $X=4.98 $Y=1.765
+ $X2=0 $Y2=0
cc_303 N_A_27_74#_c_347_p N_A_713_458#_c_781_n 0.012114f $X=4.49 $Y=0.775 $X2=0
+ $Y2=0
cc_304 N_A_27_74#_M1017_g N_A_713_458#_c_782_n 0.0117921f $X=3.105 $Y=0.835
+ $X2=0 $Y2=0
cc_305 N_A_27_74#_c_232_n N_A_713_458#_c_782_n 0.00816607f $X=3.675 $Y=1.75
+ $X2=0 $Y2=0
cc_306 N_A_27_74#_c_347_p N_A_713_458#_c_782_n 0.00338734f $X=4.49 $Y=0.775
+ $X2=0 $Y2=0
cc_307 N_A_27_74#_c_242_n N_A_561_463#_c_880_n 0.0135356f $X=4.98 $Y=2.045 $X2=0
+ $Y2=0
cc_308 N_A_27_74#_c_347_p N_A_561_463#_M1004_g 0.0075113f $X=4.49 $Y=0.775 $X2=0
+ $Y2=0
cc_309 N_A_27_74#_c_300_p N_A_561_463#_M1004_g 0.00821107f $X=4.575 $Y=0.69
+ $X2=0 $Y2=0
cc_310 N_A_27_74#_c_233_n N_A_561_463#_M1004_g 0.00466043f $X=4.66 $Y=0.34 $X2=0
+ $Y2=0
cc_311 N_A_27_74#_c_237_n N_A_561_463#_M1004_g 0.00504908f $X=5.565 $Y=0.382
+ $X2=0 $Y2=0
cc_312 N_A_27_74#_M1017_g N_A_561_463#_c_874_n 0.00521584f $X=3.105 $Y=0.835
+ $X2=0 $Y2=0
cc_313 N_A_27_74#_c_240_n N_A_561_463#_c_874_n 0.00404517f $X=3.265 $Y=2.35
+ $X2=0 $Y2=0
cc_314 N_A_27_74#_c_249_n N_A_561_463#_c_874_n 0.0261475f $X=3.59 $Y=1.915 $X2=0
+ $Y2=0
cc_315 N_A_27_74#_c_232_n N_A_561_463#_c_874_n 0.00487749f $X=3.675 $Y=1.75
+ $X2=0 $Y2=0
cc_316 N_A_27_74#_M1017_g N_A_561_463#_c_875_n 0.0172767f $X=3.105 $Y=0.835
+ $X2=0 $Y2=0
cc_317 N_A_27_74#_c_249_n N_A_561_463#_c_875_n 0.026212f $X=3.59 $Y=1.915 $X2=0
+ $Y2=0
cc_318 N_A_27_74#_c_250_n N_A_561_463#_c_875_n 0.00580943f $X=3.235 $Y=1.915
+ $X2=0 $Y2=0
cc_319 N_A_27_74#_c_232_n N_A_561_463#_c_875_n 0.0143195f $X=3.675 $Y=1.75 $X2=0
+ $Y2=0
cc_320 N_A_27_74#_c_240_n N_A_561_463#_c_882_n 0.00523114f $X=3.265 $Y=2.35
+ $X2=0 $Y2=0
cc_321 N_A_27_74#_c_241_n N_A_561_463#_c_882_n 0.00724124f $X=3.265 $Y=2.44
+ $X2=0 $Y2=0
cc_322 N_A_27_74#_c_249_n N_A_561_463#_c_882_n 0.0112019f $X=3.59 $Y=1.915 $X2=0
+ $Y2=0
cc_323 N_A_27_74#_c_250_n N_A_561_463#_c_882_n 9.85964e-19 $X=3.235 $Y=1.915
+ $X2=0 $Y2=0
cc_324 N_A_27_74#_M1017_g N_A_561_463#_c_877_n 0.0200862f $X=3.105 $Y=0.835
+ $X2=0 $Y2=0
cc_325 N_A_27_74#_c_226_n N_A_561_463#_c_877_n 0.00598289f $X=2.485 $Y=0.815
+ $X2=0 $Y2=0
cc_326 N_A_27_74#_c_228_n N_A_561_463#_c_877_n 0.00359183f $X=2.57 $Y=0.73 $X2=0
+ $Y2=0
cc_327 N_A_27_74#_c_229_n N_A_561_463#_c_877_n 0.0205117f $X=3.59 $Y=0.36 $X2=0
+ $Y2=0
cc_328 N_A_27_74#_c_231_n N_A_561_463#_c_877_n 0.00541862f $X=3.675 $Y=0.69
+ $X2=0 $Y2=0
cc_329 N_A_27_74#_c_232_n N_A_561_463#_c_877_n 0.0417773f $X=3.675 $Y=1.75 $X2=0
+ $Y2=0
cc_330 N_A_27_74#_c_298_p N_A_561_463#_c_877_n 0.0137879f $X=3.675 $Y=0.775
+ $X2=0 $Y2=0
cc_331 N_A_27_74#_c_241_n N_A_561_463#_c_884_n 0.00480202f $X=3.265 $Y=2.44
+ $X2=0 $Y2=0
cc_332 N_A_27_74#_c_249_n N_A_561_463#_c_884_n 0.0321162f $X=3.59 $Y=1.915 $X2=0
+ $Y2=0
cc_333 N_A_27_74#_c_250_n N_A_561_463#_c_884_n 0.00493382f $X=3.235 $Y=1.915
+ $X2=0 $Y2=0
cc_334 N_A_27_74#_c_249_n N_A_561_463#_c_878_n 0.0221387f $X=3.59 $Y=1.915 $X2=0
+ $Y2=0
cc_335 N_A_27_74#_c_232_n N_A_561_463#_c_878_n 0.00745226f $X=3.675 $Y=1.75
+ $X2=0 $Y2=0
cc_336 N_A_27_74#_c_245_n N_A_561_463#_c_879_n 0.00910348f $X=4.98 $Y=1.765
+ $X2=0 $Y2=0
cc_337 N_A_27_74#_c_249_n N_A_561_463#_c_879_n 7.47084e-19 $X=3.59 $Y=1.915
+ $X2=0 $Y2=0
cc_338 N_A_27_74#_c_232_n N_A_561_463#_c_879_n 4.99875e-19 $X=3.675 $Y=1.75
+ $X2=0 $Y2=0
cc_339 N_A_27_74#_M1023_g N_A_1210_314#_M1020_g 0.0487323f $X=5.765 $Y=0.83
+ $X2=0 $Y2=0
cc_340 N_A_27_74#_c_236_n N_A_1210_314#_M1020_g 0.00120024f $X=5.73 $Y=0.345
+ $X2=0 $Y2=0
cc_341 N_A_27_74#_c_243_n N_A_1210_314#_c_1003_n 0.00854279f $X=5.69 $Y=1.765
+ $X2=0 $Y2=0
cc_342 N_A_27_74#_M1023_g N_A_1210_314#_c_997_n 9.78231e-19 $X=5.765 $Y=0.83
+ $X2=0 $Y2=0
cc_343 N_A_27_74#_M1023_g N_A_1210_314#_c_998_n 0.00854279f $X=5.765 $Y=0.83
+ $X2=0 $Y2=0
cc_344 N_A_27_74#_c_242_n N_A_1011_424#_c_1117_n 0.00351148f $X=4.98 $Y=2.045
+ $X2=0 $Y2=0
cc_345 N_A_27_74#_c_245_n N_A_1011_424#_c_1117_n 0.00377355f $X=4.98 $Y=1.765
+ $X2=0 $Y2=0
cc_346 N_A_27_74#_M1023_g N_A_1011_424#_c_1123_n 0.0117759f $X=5.765 $Y=0.83
+ $X2=0 $Y2=0
cc_347 N_A_27_74#_c_235_n N_A_1011_424#_c_1123_n 0.0132333f $X=5.73 $Y=0.345
+ $X2=0 $Y2=0
cc_348 N_A_27_74#_c_236_n N_A_1011_424#_c_1123_n 0.00181648f $X=5.73 $Y=0.345
+ $X2=0 $Y2=0
cc_349 N_A_27_74#_c_237_n N_A_1011_424#_c_1123_n 0.0144503f $X=5.565 $Y=0.382
+ $X2=0 $Y2=0
cc_350 N_A_27_74#_c_243_n N_A_1011_424#_c_1118_n 0.0173146f $X=5.69 $Y=1.765
+ $X2=0 $Y2=0
cc_351 N_A_27_74#_c_243_n N_A_1011_424#_c_1119_n 0.00882584f $X=5.69 $Y=1.765
+ $X2=0 $Y2=0
cc_352 N_A_27_74#_c_245_n N_A_1011_424#_c_1119_n 9.59081e-19 $X=4.98 $Y=1.765
+ $X2=0 $Y2=0
cc_353 N_A_27_74#_M1023_g N_A_1011_424#_c_1110_n 0.00756063f $X=5.765 $Y=0.83
+ $X2=0 $Y2=0
cc_354 N_A_27_74#_c_243_n N_A_1011_424#_c_1111_n 0.00217196f $X=5.69 $Y=1.765
+ $X2=0 $Y2=0
cc_355 N_A_27_74#_M1023_g N_A_1011_424#_c_1111_n 0.0096767f $X=5.765 $Y=0.83
+ $X2=0 $Y2=0
cc_356 N_A_27_74#_M1023_g N_A_1011_424#_c_1112_n 0.00250438f $X=5.765 $Y=0.83
+ $X2=0 $Y2=0
cc_357 N_A_27_74#_M1023_g N_A_1011_424#_c_1114_n 0.00342707f $X=5.765 $Y=0.83
+ $X2=0 $Y2=0
cc_358 N_A_27_74#_c_265_n N_VPWR_M1014_d 0.00457874f $X=0.675 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_359 N_A_27_74#_c_222_n N_VPWR_M1014_d 0.0015936f $X=0.76 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_360 N_A_27_74#_c_215_n N_VPWR_c_1210_n 0.00486117f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_361 N_A_27_74#_c_247_n N_VPWR_c_1210_n 0.0449718f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_362 N_A_27_74#_c_265_n N_VPWR_c_1210_n 0.0148103f $X=0.675 $Y=2.035 $X2=0
+ $Y2=0
cc_363 N_A_27_74#_c_242_n N_VPWR_c_1213_n 0.0027945f $X=4.98 $Y=2.045 $X2=0
+ $Y2=0
cc_364 N_A_27_74#_c_215_n N_VPWR_c_1215_n 0.00444469f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_365 N_A_27_74#_c_241_n N_VPWR_c_1216_n 0.00399296f $X=3.265 $Y=2.44 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_c_215_n N_VPWR_c_1209_n 0.00858806f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_367 N_A_27_74#_c_241_n N_VPWR_c_1209_n 0.00537853f $X=3.265 $Y=2.44 $X2=0
+ $Y2=0
cc_368 N_A_27_74#_c_242_n N_VPWR_c_1209_n 0.00355626f $X=4.98 $Y=2.045 $X2=0
+ $Y2=0
cc_369 N_A_27_74#_c_247_n N_VPWR_c_1209_n 0.0120466f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_370 N_A_27_74#_c_247_n N_VPWR_c_1220_n 0.0145938f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_371 N_A_27_74#_c_215_n N_VPWR_c_1221_n 0.00276925f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_372 N_A_27_74#_c_226_n N_A_454_503#_M1006_d 0.00342102f $X=2.485 $Y=0.815
+ $X2=-0.19 $Y2=-0.245
cc_373 N_A_27_74#_c_228_n N_A_454_503#_M1006_d 0.00192055f $X=2.57 $Y=0.73
+ $X2=-0.19 $Y2=-0.245
cc_374 N_A_27_74#_M1017_g N_A_454_503#_c_1308_n 0.00328909f $X=3.105 $Y=0.835
+ $X2=0 $Y2=0
cc_375 N_A_27_74#_c_226_n N_A_454_503#_c_1309_n 0.0116776f $X=2.485 $Y=0.815
+ $X2=0 $Y2=0
cc_376 N_A_27_74#_M1017_g N_A_454_503#_c_1310_n 0.00181634f $X=3.105 $Y=0.835
+ $X2=0 $Y2=0
cc_377 N_A_27_74#_c_226_n N_A_454_503#_c_1310_n 0.00517656f $X=2.485 $Y=0.815
+ $X2=0 $Y2=0
cc_378 N_A_27_74#_c_229_n N_A_454_503#_c_1310_n 0.00926147f $X=3.59 $Y=0.36
+ $X2=0 $Y2=0
cc_379 N_A_27_74#_c_220_n N_VGND_M1022_d 8.95418e-19 $X=0.675 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_380 N_A_27_74#_c_224_n N_VGND_M1022_d 5.22721e-19 $X=1.135 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_381 N_A_27_74#_c_234_n N_VGND_M1022_d 0.0097696f $X=0.905 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_382 N_A_27_74#_c_272_n N_VGND_M1022_d 0.00582661f $X=0.905 $Y=0.96 $X2=-0.19
+ $Y2=-0.245
cc_383 N_A_27_74#_c_226_n N_VGND_M1006_s 0.00763168f $X=2.485 $Y=0.815 $X2=0
+ $Y2=0
cc_384 N_A_27_74#_c_347_p N_VGND_M1011_d 0.0112581f $X=4.49 $Y=0.775 $X2=0 $Y2=0
cc_385 N_A_27_74#_c_216_n N_VGND_c_1369_n 0.00202754f $X=1.115 $Y=1.22 $X2=0
+ $Y2=0
cc_386 N_A_27_74#_c_219_n N_VGND_c_1369_n 0.0158413f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_387 N_A_27_74#_c_220_n N_VGND_c_1369_n 0.00573342f $X=0.675 $Y=1.045 $X2=0
+ $Y2=0
cc_388 N_A_27_74#_c_224_n N_VGND_c_1369_n 0.0145677f $X=1.135 $Y=0.34 $X2=0
+ $Y2=0
cc_389 N_A_27_74#_c_234_n N_VGND_c_1369_n 0.0106391f $X=0.905 $Y=1.045 $X2=0
+ $Y2=0
cc_390 N_A_27_74#_c_272_n N_VGND_c_1369_n 0.0272627f $X=0.905 $Y=0.96 $X2=0
+ $Y2=0
cc_391 N_A_27_74#_c_223_n N_VGND_c_1370_n 0.0150375f $X=1.645 $Y=0.34 $X2=0
+ $Y2=0
cc_392 N_A_27_74#_c_225_n N_VGND_c_1370_n 0.0106642f $X=1.73 $Y=0.73 $X2=0 $Y2=0
cc_393 N_A_27_74#_c_226_n N_VGND_c_1370_n 0.0257465f $X=2.485 $Y=0.815 $X2=0
+ $Y2=0
cc_394 N_A_27_74#_c_228_n N_VGND_c_1370_n 0.00872018f $X=2.57 $Y=0.73 $X2=0
+ $Y2=0
cc_395 N_A_27_74#_c_230_n N_VGND_c_1370_n 0.0150385f $X=2.655 $Y=0.36 $X2=0
+ $Y2=0
cc_396 N_A_27_74#_c_229_n N_VGND_c_1371_n 0.0096942f $X=3.59 $Y=0.36 $X2=0 $Y2=0
cc_397 N_A_27_74#_c_231_n N_VGND_c_1371_n 0.00335995f $X=3.675 $Y=0.69 $X2=0
+ $Y2=0
cc_398 N_A_27_74#_c_347_p N_VGND_c_1371_n 0.0191408f $X=4.49 $Y=0.775 $X2=0
+ $Y2=0
cc_399 N_A_27_74#_c_233_n N_VGND_c_1371_n 0.0121213f $X=4.66 $Y=0.34 $X2=0 $Y2=0
cc_400 N_A_27_74#_M1023_g N_VGND_c_1372_n 0.00198934f $X=5.765 $Y=0.83 $X2=0
+ $Y2=0
cc_401 N_A_27_74#_c_235_n N_VGND_c_1372_n 0.0124765f $X=5.73 $Y=0.345 $X2=0
+ $Y2=0
cc_402 N_A_27_74#_c_236_n N_VGND_c_1372_n 0.00337434f $X=5.73 $Y=0.345 $X2=0
+ $Y2=0
cc_403 N_A_27_74#_c_347_p N_VGND_c_1374_n 0.00261614f $X=4.49 $Y=0.775 $X2=0
+ $Y2=0
cc_404 N_A_27_74#_c_233_n N_VGND_c_1374_n 0.0116816f $X=4.66 $Y=0.34 $X2=0 $Y2=0
cc_405 N_A_27_74#_c_236_n N_VGND_c_1374_n 0.00653686f $X=5.73 $Y=0.345 $X2=0
+ $Y2=0
cc_406 N_A_27_74#_c_237_n N_VGND_c_1374_n 0.0789953f $X=5.565 $Y=0.382 $X2=0
+ $Y2=0
cc_407 N_A_27_74#_c_219_n N_VGND_c_1376_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_408 N_A_27_74#_c_216_n N_VGND_c_1377_n 0.00278179f $X=1.115 $Y=1.22 $X2=0
+ $Y2=0
cc_409 N_A_27_74#_c_223_n N_VGND_c_1377_n 0.0440512f $X=1.645 $Y=0.34 $X2=0
+ $Y2=0
cc_410 N_A_27_74#_c_224_n N_VGND_c_1377_n 0.0118529f $X=1.135 $Y=0.34 $X2=0
+ $Y2=0
cc_411 N_A_27_74#_c_226_n N_VGND_c_1377_n 0.00254217f $X=2.485 $Y=0.815 $X2=0
+ $Y2=0
cc_412 N_A_27_74#_c_226_n N_VGND_c_1378_n 0.00192775f $X=2.485 $Y=0.815 $X2=0
+ $Y2=0
cc_413 N_A_27_74#_c_229_n N_VGND_c_1378_n 0.0638335f $X=3.59 $Y=0.36 $X2=0 $Y2=0
cc_414 N_A_27_74#_c_230_n N_VGND_c_1378_n 0.0107439f $X=2.655 $Y=0.36 $X2=0
+ $Y2=0
cc_415 N_A_27_74#_c_347_p N_VGND_c_1378_n 0.00384226f $X=4.49 $Y=0.775 $X2=0
+ $Y2=0
cc_416 N_A_27_74#_c_216_n N_VGND_c_1381_n 0.00356272f $X=1.115 $Y=1.22 $X2=0
+ $Y2=0
cc_417 N_A_27_74#_c_219_n N_VGND_c_1381_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_418 N_A_27_74#_c_223_n N_VGND_c_1381_n 0.0245464f $X=1.645 $Y=0.34 $X2=0
+ $Y2=0
cc_419 N_A_27_74#_c_224_n N_VGND_c_1381_n 0.00617452f $X=1.135 $Y=0.34 $X2=0
+ $Y2=0
cc_420 N_A_27_74#_c_226_n N_VGND_c_1381_n 0.00888428f $X=2.485 $Y=0.815 $X2=0
+ $Y2=0
cc_421 N_A_27_74#_c_229_n N_VGND_c_1381_n 0.0371527f $X=3.59 $Y=0.36 $X2=0 $Y2=0
cc_422 N_A_27_74#_c_230_n N_VGND_c_1381_n 0.00585125f $X=2.655 $Y=0.36 $X2=0
+ $Y2=0
cc_423 N_A_27_74#_c_347_p N_VGND_c_1381_n 0.0140465f $X=4.49 $Y=0.775 $X2=0
+ $Y2=0
cc_424 N_A_27_74#_c_233_n N_VGND_c_1381_n 0.00606295f $X=4.66 $Y=0.34 $X2=0
+ $Y2=0
cc_425 N_A_27_74#_c_236_n N_VGND_c_1381_n 0.0102677f $X=5.73 $Y=0.345 $X2=0
+ $Y2=0
cc_426 N_A_27_74#_c_237_n N_VGND_c_1381_n 0.0448715f $X=5.565 $Y=0.382 $X2=0
+ $Y2=0
cc_427 N_A_27_74#_c_231_n A_731_101# 0.00204684f $X=3.675 $Y=0.69 $X2=-0.19
+ $Y2=-0.245
cc_428 N_A_27_74#_c_232_n A_731_101# 7.15614e-19 $X=3.675 $Y=1.75 $X2=-0.19
+ $Y2=-0.245
cc_429 N_A_27_74#_c_347_p A_731_101# 0.00153437f $X=4.49 $Y=0.775 $X2=-0.19
+ $Y2=-0.245
cc_430 N_D_c_493_n N_A_206_368#_c_540_n 0.00966037f $X=2.445 $Y=1.125 $X2=0
+ $Y2=0
cc_431 N_D_c_496_n N_A_206_368#_c_553_n 0.0266665f $X=2.195 $Y=2.44 $X2=0 $Y2=0
cc_432 N_D_c_494_n N_A_206_368#_c_553_n 0.0292902f $X=2.135 $Y=1.29 $X2=0 $Y2=0
cc_433 N_D_c_495_n N_A_206_368#_c_553_n 0.0146252f $X=2.135 $Y=1.29 $X2=0 $Y2=0
cc_434 D N_A_206_368#_c_553_n 6.61663e-19 $X=2.16 $Y=2.035 $X2=0 $Y2=0
cc_435 N_D_c_496_n N_A_206_368#_c_554_n 0.00587014f $X=2.195 $Y=2.44 $X2=0 $Y2=0
cc_436 N_D_c_496_n N_A_206_368#_c_555_n 0.0126627f $X=2.195 $Y=2.44 $X2=0 $Y2=0
cc_437 N_D_c_496_n N_A_206_368#_c_557_n 0.00643962f $X=2.195 $Y=2.44 $X2=0 $Y2=0
cc_438 N_D_c_495_n N_A_206_368#_c_544_n 0.00745251f $X=2.135 $Y=1.29 $X2=0 $Y2=0
cc_439 N_D_c_496_n N_A_206_368#_c_558_n 0.00129002f $X=2.195 $Y=2.44 $X2=0 $Y2=0
cc_440 D N_A_206_368#_c_558_n 0.0107463f $X=2.16 $Y=2.035 $X2=0 $Y2=0
cc_441 N_D_c_496_n N_A_206_368#_c_559_n 0.00534435f $X=2.195 $Y=2.44 $X2=0 $Y2=0
cc_442 N_D_c_496_n N_A_206_368#_c_563_n 0.00681776f $X=2.195 $Y=2.44 $X2=0 $Y2=0
cc_443 D N_A_206_368#_c_563_n 0.0144543f $X=2.16 $Y=2.035 $X2=0 $Y2=0
cc_444 N_D_c_495_n N_A_206_368#_c_564_n 0.0123923f $X=2.135 $Y=1.29 $X2=0 $Y2=0
cc_445 N_D_c_494_n N_A_206_368#_c_548_n 3.62223e-19 $X=2.135 $Y=1.29 $X2=0 $Y2=0
cc_446 N_D_c_495_n N_A_206_368#_c_548_n 0.0220028f $X=2.135 $Y=1.29 $X2=0 $Y2=0
cc_447 N_D_c_495_n N_A_206_368#_c_549_n 9.76154e-19 $X=2.135 $Y=1.29 $X2=0 $Y2=0
cc_448 N_D_c_496_n N_A_206_368#_c_567_n 0.0157162f $X=2.195 $Y=2.44 $X2=0 $Y2=0
cc_449 D N_A_206_368#_c_567_n 0.00827903f $X=2.16 $Y=2.035 $X2=0 $Y2=0
cc_450 N_D_c_493_n N_A_206_368#_c_552_n 0.011002f $X=2.445 $Y=1.125 $X2=0 $Y2=0
cc_451 N_D_c_494_n N_A_206_368#_c_552_n 0.0206359f $X=2.135 $Y=1.29 $X2=0 $Y2=0
cc_452 N_D_c_495_n N_A_206_368#_c_552_n 8.43694e-19 $X=2.135 $Y=1.29 $X2=0 $Y2=0
cc_453 N_D_c_493_n N_A_561_463#_c_877_n 0.00113547f $X=2.445 $Y=1.125 $X2=0
+ $Y2=0
cc_454 N_D_c_496_n N_VPWR_c_1216_n 0.00399229f $X=2.195 $Y=2.44 $X2=0 $Y2=0
cc_455 N_D_c_496_n N_VPWR_c_1209_n 0.00537853f $X=2.195 $Y=2.44 $X2=0 $Y2=0
cc_456 N_D_c_496_n N_VPWR_c_1221_n 0.00355987f $X=2.195 $Y=2.44 $X2=0 $Y2=0
cc_457 N_D_c_496_n N_A_454_503#_c_1308_n 0.0086914f $X=2.195 $Y=2.44 $X2=0 $Y2=0
cc_458 N_D_c_494_n N_A_454_503#_c_1308_n 0.00690033f $X=2.135 $Y=1.29 $X2=0
+ $Y2=0
cc_459 N_D_c_495_n N_A_454_503#_c_1308_n 0.0842118f $X=2.135 $Y=1.29 $X2=0 $Y2=0
cc_460 N_D_c_493_n N_A_454_503#_c_1309_n 0.00392055f $X=2.445 $Y=1.125 $X2=0
+ $Y2=0
cc_461 N_D_c_494_n N_A_454_503#_c_1309_n 0.00458046f $X=2.135 $Y=1.29 $X2=0
+ $Y2=0
cc_462 N_D_c_495_n N_A_454_503#_c_1309_n 0.00892592f $X=2.135 $Y=1.29 $X2=0
+ $Y2=0
cc_463 N_D_c_493_n N_VGND_c_1370_n 0.0010673f $X=2.445 $Y=1.125 $X2=0 $Y2=0
cc_464 N_D_c_493_n N_VGND_c_1381_n 7.22543e-19 $X=2.445 $Y=1.125 $X2=0 $Y2=0
cc_465 N_A_206_368#_c_606_n N_A_713_458#_M1018_d 0.0166057f $X=4.78 $Y=2.71
+ $X2=0 $Y2=0
cc_466 N_A_206_368#_c_545_n N_A_713_458#_M1018_d 0.00554389f $X=4.865 $Y=2.625
+ $X2=0 $Y2=0
cc_467 N_A_206_368#_c_569_n N_A_713_458#_M1018_d 0.00284573f $X=4.865 $Y=2.71
+ $X2=0 $Y2=0
cc_468 N_A_206_368#_M1016_g N_A_713_458#_M1011_g 0.040722f $X=3.58 $Y=0.715
+ $X2=0 $Y2=0
cc_469 N_A_206_368#_c_606_n N_A_713_458#_c_784_n 0.01086f $X=4.78 $Y=2.71 $X2=0
+ $Y2=0
cc_470 N_A_206_368#_c_568_n N_A_713_458#_c_784_n 0.00386441f $X=3.375 $Y=2.71
+ $X2=0 $Y2=0
cc_471 N_A_206_368#_c_543_n N_A_713_458#_c_778_n 0.0024606f $X=5.13 $Y=1.15
+ $X2=0 $Y2=0
cc_472 N_A_206_368#_c_546_n N_A_713_458#_c_778_n 0.00414536f $X=5.17 $Y=1.455
+ $X2=0 $Y2=0
cc_473 N_A_206_368#_c_547_n N_A_713_458#_c_778_n 0.0153318f $X=4.95 $Y=1.455
+ $X2=0 $Y2=0
cc_474 N_A_206_368#_c_550_n N_A_713_458#_c_778_n 0.00419808f $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_475 N_A_206_368#_c_606_n N_A_713_458#_c_824_n 0.0172511f $X=4.78 $Y=2.71
+ $X2=0 $Y2=0
cc_476 N_A_206_368#_c_545_n N_A_713_458#_c_780_n 0.0679022f $X=4.865 $Y=2.625
+ $X2=0 $Y2=0
cc_477 N_A_206_368#_c_547_n N_A_713_458#_c_780_n 0.0130528f $X=4.95 $Y=1.455
+ $X2=0 $Y2=0
cc_478 N_A_206_368#_c_550_n N_A_713_458#_c_780_n 0.0045377f $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_479 N_A_206_368#_c_551_n N_A_713_458#_c_780_n 7.59146e-19 $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_480 N_A_206_368#_M1016_g N_A_713_458#_c_782_n 0.00294341f $X=3.58 $Y=0.715
+ $X2=0 $Y2=0
cc_481 N_A_206_368#_c_559_n N_A_561_463#_M1021_d 0.00241932f $X=3.29 $Y=2.88
+ $X2=0 $Y2=0
cc_482 N_A_206_368#_c_606_n N_A_561_463#_c_880_n 0.0159167f $X=4.78 $Y=2.71
+ $X2=0 $Y2=0
cc_483 N_A_206_368#_c_545_n N_A_561_463#_c_880_n 0.00277241f $X=4.865 $Y=2.625
+ $X2=0 $Y2=0
cc_484 N_A_206_368#_c_569_n N_A_561_463#_c_880_n 0.00393225f $X=4.865 $Y=2.71
+ $X2=0 $Y2=0
cc_485 N_A_206_368#_c_545_n N_A_561_463#_c_871_n 0.0040355f $X=4.865 $Y=2.625
+ $X2=0 $Y2=0
cc_486 N_A_206_368#_c_547_n N_A_561_463#_c_871_n 0.00146346f $X=4.95 $Y=1.455
+ $X2=0 $Y2=0
cc_487 N_A_206_368#_c_551_n N_A_561_463#_c_871_n 7.0989e-19 $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_488 N_A_206_368#_c_543_n N_A_561_463#_M1004_g 0.0132876f $X=5.13 $Y=1.15
+ $X2=0 $Y2=0
cc_489 N_A_206_368#_c_550_n N_A_561_463#_M1004_g 5.7185e-19 $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_490 N_A_206_368#_c_547_n N_A_561_463#_c_873_n 6.71581e-19 $X=4.95 $Y=1.455
+ $X2=0 $Y2=0
cc_491 N_A_206_368#_c_551_n N_A_561_463#_c_873_n 0.0132876f $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_492 N_A_206_368#_c_553_n N_A_561_463#_c_874_n 0.00472003f $X=2.64 $Y=1.74
+ $X2=0 $Y2=0
cc_493 N_A_206_368#_c_554_n N_A_561_463#_c_874_n 0.00633941f $X=2.73 $Y=2.15
+ $X2=0 $Y2=0
cc_494 N_A_206_368#_c_555_n N_A_561_463#_c_874_n 0.00319034f $X=2.73 $Y=2.24
+ $X2=0 $Y2=0
cc_495 N_A_206_368#_c_559_n N_A_561_463#_c_882_n 0.00578093f $X=3.29 $Y=2.88
+ $X2=0 $Y2=0
cc_496 N_A_206_368#_c_606_n N_A_561_463#_c_882_n 0.0463133f $X=4.78 $Y=2.71
+ $X2=0 $Y2=0
cc_497 N_A_206_368#_c_568_n N_A_561_463#_c_882_n 0.0105359f $X=3.375 $Y=2.71
+ $X2=0 $Y2=0
cc_498 N_A_206_368#_M1016_g N_A_561_463#_c_877_n 0.00185496f $X=3.58 $Y=0.715
+ $X2=0 $Y2=0
cc_499 N_A_206_368#_c_555_n N_A_561_463#_c_884_n 0.00523332f $X=2.73 $Y=2.24
+ $X2=0 $Y2=0
cc_500 N_A_206_368#_c_559_n N_A_561_463#_c_884_n 0.0241581f $X=3.29 $Y=2.88
+ $X2=0 $Y2=0
cc_501 N_A_206_368#_c_606_n N_A_561_463#_c_878_n 0.00232465f $X=4.78 $Y=2.71
+ $X2=0 $Y2=0
cc_502 N_A_206_368#_c_606_n N_A_561_463#_c_879_n 5.30241e-19 $X=4.78 $Y=2.71
+ $X2=0 $Y2=0
cc_503 N_A_206_368#_c_556_n N_A_1210_314#_c_1001_n 0.0119305f $X=5.515 $Y=2.465
+ $X2=0 $Y2=0
cc_504 N_A_206_368#_c_561_n N_A_1210_314#_c_1001_n 0.001726f $X=5.51 $Y=2.99
+ $X2=0 $Y2=0
cc_505 N_A_206_368#_c_562_n N_A_1210_314#_c_1001_n 0.00486501f $X=5.675 $Y=2.215
+ $X2=0 $Y2=0
cc_506 N_A_206_368#_c_556_n N_A_1210_314#_c_1003_n 0.0228354f $X=5.515 $Y=2.465
+ $X2=0 $Y2=0
cc_507 N_A_206_368#_c_562_n N_A_1210_314#_c_1003_n 0.00366101f $X=5.675 $Y=2.215
+ $X2=0 $Y2=0
cc_508 N_A_206_368#_c_556_n N_A_1210_314#_c_997_n 6.90151e-19 $X=5.515 $Y=2.465
+ $X2=0 $Y2=0
cc_509 N_A_206_368#_c_562_n N_A_1210_314#_c_997_n 0.0120093f $X=5.675 $Y=2.215
+ $X2=0 $Y2=0
cc_510 N_A_206_368#_c_561_n N_A_1011_424#_M1019_d 0.00579062f $X=5.51 $Y=2.99
+ $X2=0 $Y2=0
cc_511 N_A_206_368#_c_556_n N_A_1011_424#_c_1117_n 0.00555548f $X=5.515 $Y=2.465
+ $X2=0 $Y2=0
cc_512 N_A_206_368#_c_545_n N_A_1011_424#_c_1117_n 0.0602335f $X=4.865 $Y=2.625
+ $X2=0 $Y2=0
cc_513 N_A_206_368#_c_561_n N_A_1011_424#_c_1117_n 0.012787f $X=5.51 $Y=2.99
+ $X2=0 $Y2=0
cc_514 N_A_206_368#_c_562_n N_A_1011_424#_c_1117_n 0.0415397f $X=5.675 $Y=2.215
+ $X2=0 $Y2=0
cc_515 N_A_206_368#_c_550_n N_A_1011_424#_c_1123_n 0.0184109f $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_516 N_A_206_368#_c_551_n N_A_1011_424#_c_1123_n 0.00177816f $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_517 N_A_206_368#_c_556_n N_A_1011_424#_c_1118_n 0.00284269f $X=5.515 $Y=2.465
+ $X2=0 $Y2=0
cc_518 N_A_206_368#_c_562_n N_A_1011_424#_c_1118_n 0.0261799f $X=5.675 $Y=2.215
+ $X2=0 $Y2=0
cc_519 N_A_206_368#_c_550_n N_A_1011_424#_c_1118_n 0.014508f $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_520 N_A_206_368#_c_551_n N_A_1011_424#_c_1118_n 2.02945e-19 $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_521 N_A_206_368#_c_545_n N_A_1011_424#_c_1119_n 0.013162f $X=4.865 $Y=2.625
+ $X2=0 $Y2=0
cc_522 N_A_206_368#_c_546_n N_A_1011_424#_c_1119_n 0.00399569f $X=5.17 $Y=1.455
+ $X2=0 $Y2=0
cc_523 N_A_206_368#_c_550_n N_A_1011_424#_c_1119_n 0.0101622f $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_524 N_A_206_368#_c_543_n N_A_1011_424#_c_1110_n 0.00102454f $X=5.13 $Y=1.15
+ $X2=0 $Y2=0
cc_525 N_A_206_368#_c_550_n N_A_1011_424#_c_1110_n 0.00594629f $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_526 N_A_206_368#_c_551_n N_A_1011_424#_c_1110_n 4.343e-19 $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_527 N_A_206_368#_c_550_n N_A_1011_424#_c_1111_n 0.0106791f $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_528 N_A_206_368#_c_551_n N_A_1011_424#_c_1111_n 4.343e-19 $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_529 N_A_206_368#_c_550_n N_A_1011_424#_c_1112_n 0.0142756f $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_530 N_A_206_368#_c_551_n N_A_1011_424#_c_1112_n 0.0010737f $X=5.315 $Y=1.315
+ $X2=0 $Y2=0
cc_531 N_A_206_368#_c_562_n N_A_1011_424#_c_1114_n 4.59501e-19 $X=5.675 $Y=2.215
+ $X2=0 $Y2=0
cc_532 N_A_206_368#_c_558_n N_VPWR_M1012_s 0.0212312f $X=2.08 $Y=2.71 $X2=0
+ $Y2=0
cc_533 N_A_206_368#_c_606_n N_VPWR_M1000_d 0.00824604f $X=4.78 $Y=2.71 $X2=0
+ $Y2=0
cc_534 N_A_206_368#_c_557_n N_VPWR_c_1210_n 0.046267f $X=1.245 $Y=2.625 $X2=0
+ $Y2=0
cc_535 N_A_206_368#_c_556_n N_VPWR_c_1211_n 5.11441e-19 $X=5.515 $Y=2.465 $X2=0
+ $Y2=0
cc_536 N_A_206_368#_c_561_n N_VPWR_c_1211_n 0.00809786f $X=5.51 $Y=2.99 $X2=0
+ $Y2=0
cc_537 N_A_206_368#_c_562_n N_VPWR_c_1211_n 0.0168084f $X=5.675 $Y=2.215 $X2=0
+ $Y2=0
cc_538 N_A_206_368#_c_556_n N_VPWR_c_1213_n 0.00278193f $X=5.515 $Y=2.465 $X2=0
+ $Y2=0
cc_539 N_A_206_368#_c_606_n N_VPWR_c_1213_n 0.0131309f $X=4.78 $Y=2.71 $X2=0
+ $Y2=0
cc_540 N_A_206_368#_c_561_n N_VPWR_c_1213_n 0.0588814f $X=5.51 $Y=2.99 $X2=0
+ $Y2=0
cc_541 N_A_206_368#_c_569_n N_VPWR_c_1213_n 0.0118887f $X=4.865 $Y=2.71 $X2=0
+ $Y2=0
cc_542 N_A_206_368#_c_557_n N_VPWR_c_1215_n 0.0179726f $X=1.245 $Y=2.625 $X2=0
+ $Y2=0
cc_543 N_A_206_368#_c_558_n N_VPWR_c_1215_n 0.00228036f $X=2.08 $Y=2.71 $X2=0
+ $Y2=0
cc_544 N_A_206_368#_c_555_n N_VPWR_c_1216_n 6.57382e-19 $X=2.73 $Y=2.24 $X2=0
+ $Y2=0
cc_545 N_A_206_368#_c_558_n N_VPWR_c_1216_n 0.00360091f $X=2.08 $Y=2.71 $X2=0
+ $Y2=0
cc_546 N_A_206_368#_c_559_n N_VPWR_c_1216_n 0.039311f $X=3.29 $Y=2.88 $X2=0
+ $Y2=0
cc_547 N_A_206_368#_c_606_n N_VPWR_c_1216_n 0.00627628f $X=4.78 $Y=2.71 $X2=0
+ $Y2=0
cc_548 N_A_206_368#_c_567_n N_VPWR_c_1216_n 0.00638941f $X=2.165 $Y=2.71 $X2=0
+ $Y2=0
cc_549 N_A_206_368#_c_568_n N_VPWR_c_1216_n 0.00660141f $X=3.375 $Y=2.71 $X2=0
+ $Y2=0
cc_550 N_A_206_368#_c_556_n N_VPWR_c_1209_n 0.00356044f $X=5.515 $Y=2.465 $X2=0
+ $Y2=0
cc_551 N_A_206_368#_c_557_n N_VPWR_c_1209_n 0.0163583f $X=1.245 $Y=2.625 $X2=0
+ $Y2=0
cc_552 N_A_206_368#_c_558_n N_VPWR_c_1209_n 0.0102379f $X=2.08 $Y=2.71 $X2=0
+ $Y2=0
cc_553 N_A_206_368#_c_559_n N_VPWR_c_1209_n 0.0363011f $X=3.29 $Y=2.88 $X2=0
+ $Y2=0
cc_554 N_A_206_368#_c_606_n N_VPWR_c_1209_n 0.0315431f $X=4.78 $Y=2.71 $X2=0
+ $Y2=0
cc_555 N_A_206_368#_c_561_n N_VPWR_c_1209_n 0.0327139f $X=5.51 $Y=2.99 $X2=0
+ $Y2=0
cc_556 N_A_206_368#_c_567_n N_VPWR_c_1209_n 0.0059026f $X=2.165 $Y=2.71 $X2=0
+ $Y2=0
cc_557 N_A_206_368#_c_568_n N_VPWR_c_1209_n 0.00596797f $X=3.375 $Y=2.71 $X2=0
+ $Y2=0
cc_558 N_A_206_368#_c_569_n N_VPWR_c_1209_n 0.00633012f $X=4.865 $Y=2.71 $X2=0
+ $Y2=0
cc_559 N_A_206_368#_c_557_n N_VPWR_c_1221_n 0.00101596f $X=1.245 $Y=2.625 $X2=0
+ $Y2=0
cc_560 N_A_206_368#_c_558_n N_VPWR_c_1221_n 0.0245924f $X=2.08 $Y=2.71 $X2=0
+ $Y2=0
cc_561 N_A_206_368#_c_606_n N_VPWR_c_1222_n 0.0242026f $X=4.78 $Y=2.71 $X2=0
+ $Y2=0
cc_562 N_A_206_368#_c_569_n N_VPWR_c_1222_n 0.00338029f $X=4.865 $Y=2.71 $X2=0
+ $Y2=0
cc_563 N_A_206_368#_c_559_n N_A_454_503#_M1012_d 0.00499081f $X=3.29 $Y=2.88
+ $X2=0 $Y2=0
cc_564 N_A_206_368#_c_553_n N_A_454_503#_c_1308_n 0.0135006f $X=2.64 $Y=1.74
+ $X2=0 $Y2=0
cc_565 N_A_206_368#_c_554_n N_A_454_503#_c_1308_n 0.00655506f $X=2.73 $Y=2.15
+ $X2=0 $Y2=0
cc_566 N_A_206_368#_c_555_n N_A_454_503#_c_1308_n 0.00146414f $X=2.73 $Y=2.24
+ $X2=0 $Y2=0
cc_567 N_A_206_368#_c_559_n N_A_454_503#_c_1308_n 0.0131313f $X=3.29 $Y=2.88
+ $X2=0 $Y2=0
cc_568 N_A_206_368#_c_552_n N_A_454_503#_c_1309_n 2.66553e-19 $X=1.595 $Y=1.35
+ $X2=0 $Y2=0
cc_569 N_A_206_368#_c_553_n N_A_454_503#_c_1310_n 0.00532338f $X=2.64 $Y=1.74
+ $X2=0 $Y2=0
cc_570 N_A_206_368#_c_606_n A_668_503# 0.00203787f $X=4.78 $Y=2.71 $X2=-0.19
+ $Y2=-0.245
cc_571 N_A_206_368#_c_568_n A_668_503# 0.00262938f $X=3.375 $Y=2.71 $X2=-0.19
+ $Y2=-0.245
cc_572 N_A_206_368#_c_561_n A_1118_508# 8.83155e-19 $X=5.51 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_573 N_A_206_368#_c_562_n A_1118_508# 0.00558111f $X=5.675 $Y=2.215 $X2=-0.19
+ $Y2=-0.245
cc_574 N_A_206_368#_c_540_n N_VGND_c_1370_n 0.0246014f $X=3.505 $Y=0.18 $X2=0
+ $Y2=0
cc_575 N_A_206_368#_c_552_n N_VGND_c_1370_n 0.00115203f $X=1.595 $Y=1.35 $X2=0
+ $Y2=0
cc_576 N_A_206_368#_c_540_n N_VGND_c_1371_n 0.00365801f $X=3.505 $Y=0.18 $X2=0
+ $Y2=0
cc_577 N_A_206_368#_M1016_g N_VGND_c_1371_n 5.83992e-19 $X=3.58 $Y=0.715 $X2=0
+ $Y2=0
cc_578 N_A_206_368#_c_543_n N_VGND_c_1374_n 7.26245e-19 $X=5.13 $Y=1.15 $X2=0
+ $Y2=0
cc_579 N_A_206_368#_c_541_n N_VGND_c_1377_n 0.00932626f $X=1.76 $Y=0.18 $X2=0
+ $Y2=0
cc_580 N_A_206_368#_c_540_n N_VGND_c_1378_n 0.0290765f $X=3.505 $Y=0.18 $X2=0
+ $Y2=0
cc_581 N_A_206_368#_c_540_n N_VGND_c_1381_n 0.0403312f $X=3.505 $Y=0.18 $X2=0
+ $Y2=0
cc_582 N_A_206_368#_c_541_n N_VGND_c_1381_n 0.00600554f $X=1.76 $Y=0.18 $X2=0
+ $Y2=0
cc_583 N_A_713_458#_c_776_n N_A_561_463#_c_880_n 0.00766958f $X=3.662 $Y=2.29
+ $X2=0 $Y2=0
cc_584 N_A_713_458#_c_784_n N_A_561_463#_c_880_n 0.0163093f $X=3.662 $Y=2.44
+ $X2=0 $Y2=0
cc_585 N_A_713_458#_c_824_n N_A_561_463#_c_880_n 0.00413011f $X=4.51 $Y=2.29
+ $X2=0 $Y2=0
cc_586 N_A_713_458#_c_780_n N_A_561_463#_c_880_n 8.53938e-19 $X=4.472 $Y=2.125
+ $X2=0 $Y2=0
cc_587 N_A_713_458#_c_780_n N_A_561_463#_c_871_n 0.00545385f $X=4.472 $Y=2.125
+ $X2=0 $Y2=0
cc_588 N_A_713_458#_M1011_g N_A_561_463#_M1004_g 0.0138258f $X=3.94 $Y=0.715
+ $X2=0 $Y2=0
cc_589 N_A_713_458#_c_778_n N_A_561_463#_M1004_g 0.00843882f $X=4.83 $Y=1.115
+ $X2=0 $Y2=0
cc_590 N_A_713_458#_c_803_n N_A_561_463#_M1004_g 0.00560514f $X=4.915 $Y=0.825
+ $X2=0 $Y2=0
cc_591 N_A_713_458#_c_779_n N_A_561_463#_M1004_g 2.6853e-19 $X=4.095 $Y=1.115
+ $X2=0 $Y2=0
cc_592 N_A_713_458#_c_780_n N_A_561_463#_M1004_g 0.00268861f $X=4.472 $Y=2.125
+ $X2=0 $Y2=0
cc_593 N_A_713_458#_c_781_n N_A_561_463#_M1004_g 0.00412415f $X=4.525 $Y=1.115
+ $X2=0 $Y2=0
cc_594 N_A_713_458#_c_782_n N_A_561_463#_M1004_g 0.00937479f $X=3.94 $Y=1.25
+ $X2=0 $Y2=0
cc_595 N_A_713_458#_c_780_n N_A_561_463#_c_873_n 0.00501148f $X=4.472 $Y=2.125
+ $X2=0 $Y2=0
cc_596 N_A_713_458#_c_782_n N_A_561_463#_c_873_n 0.00636638f $X=3.94 $Y=1.25
+ $X2=0 $Y2=0
cc_597 N_A_713_458#_c_782_n N_A_561_463#_c_875_n 7.10477e-19 $X=3.94 $Y=1.25
+ $X2=0 $Y2=0
cc_598 N_A_713_458#_c_776_n N_A_561_463#_c_882_n 0.00228592f $X=3.662 $Y=2.29
+ $X2=0 $Y2=0
cc_599 N_A_713_458#_c_784_n N_A_561_463#_c_882_n 0.0101435f $X=3.662 $Y=2.44
+ $X2=0 $Y2=0
cc_600 N_A_713_458#_c_824_n N_A_561_463#_c_882_n 0.0124674f $X=4.51 $Y=2.29
+ $X2=0 $Y2=0
cc_601 N_A_713_458#_M1011_g N_A_561_463#_c_877_n 3.06794e-19 $X=3.94 $Y=0.715
+ $X2=0 $Y2=0
cc_602 N_A_713_458#_c_782_n N_A_561_463#_c_877_n 5.19731e-19 $X=3.94 $Y=1.25
+ $X2=0 $Y2=0
cc_603 N_A_713_458#_c_776_n N_A_561_463#_c_883_n 0.00478354f $X=3.662 $Y=2.29
+ $X2=0 $Y2=0
cc_604 N_A_713_458#_c_824_n N_A_561_463#_c_883_n 0.0104458f $X=4.51 $Y=2.29
+ $X2=0 $Y2=0
cc_605 N_A_713_458#_c_780_n N_A_561_463#_c_883_n 0.00854771f $X=4.472 $Y=2.125
+ $X2=0 $Y2=0
cc_606 N_A_713_458#_c_776_n N_A_561_463#_c_878_n 6.38789e-19 $X=3.662 $Y=2.29
+ $X2=0 $Y2=0
cc_607 N_A_713_458#_c_777_n N_A_561_463#_c_878_n 3.4162e-19 $X=4.44 $Y=1.115
+ $X2=0 $Y2=0
cc_608 N_A_713_458#_c_779_n N_A_561_463#_c_878_n 0.0192551f $X=4.095 $Y=1.115
+ $X2=0 $Y2=0
cc_609 N_A_713_458#_c_780_n N_A_561_463#_c_878_n 0.0240591f $X=4.472 $Y=2.125
+ $X2=0 $Y2=0
cc_610 N_A_713_458#_c_782_n N_A_561_463#_c_878_n 3.61728e-19 $X=3.94 $Y=1.25
+ $X2=0 $Y2=0
cc_611 N_A_713_458#_c_776_n N_A_561_463#_c_879_n 0.0227048f $X=3.662 $Y=2.29
+ $X2=0 $Y2=0
cc_612 N_A_713_458#_c_777_n N_A_561_463#_c_879_n 0.00501112f $X=4.44 $Y=1.115
+ $X2=0 $Y2=0
cc_613 N_A_713_458#_c_779_n N_A_561_463#_c_879_n 3.62853e-19 $X=4.095 $Y=1.115
+ $X2=0 $Y2=0
cc_614 N_A_713_458#_c_824_n N_A_561_463#_c_879_n 0.00159933f $X=4.51 $Y=2.29
+ $X2=0 $Y2=0
cc_615 N_A_713_458#_c_780_n N_A_561_463#_c_879_n 0.0136537f $X=4.472 $Y=2.125
+ $X2=0 $Y2=0
cc_616 N_A_713_458#_c_782_n N_A_561_463#_c_879_n 0.0188551f $X=3.94 $Y=1.25
+ $X2=0 $Y2=0
cc_617 N_A_713_458#_c_778_n N_A_1011_424#_c_1110_n 0.00355585f $X=4.83 $Y=1.115
+ $X2=0 $Y2=0
cc_618 N_A_713_458#_c_784_n N_VPWR_c_1216_n 0.00418282f $X=3.662 $Y=2.44 $X2=0
+ $Y2=0
cc_619 N_A_713_458#_c_784_n N_VPWR_c_1209_n 0.00537853f $X=3.662 $Y=2.44 $X2=0
+ $Y2=0
cc_620 N_A_713_458#_c_784_n N_VPWR_c_1222_n 0.00288568f $X=3.662 $Y=2.44 $X2=0
+ $Y2=0
cc_621 N_A_713_458#_M1011_g N_VGND_c_1371_n 0.00170921f $X=3.94 $Y=0.715 $X2=0
+ $Y2=0
cc_622 N_A_713_458#_M1011_g N_VGND_c_1378_n 0.00376447f $X=3.94 $Y=0.715 $X2=0
+ $Y2=0
cc_623 N_A_713_458#_M1011_g N_VGND_c_1381_n 0.00503886f $X=3.94 $Y=0.715 $X2=0
+ $Y2=0
cc_624 N_A_561_463#_c_882_n N_VPWR_M1000_d 0.00685193f $X=3.97 $Y=2.37 $X2=0
+ $Y2=0
cc_625 N_A_561_463#_c_883_n N_VPWR_M1000_d 0.00475776f $X=4.055 $Y=2.285 $X2=0
+ $Y2=0
cc_626 N_A_561_463#_c_880_n N_VPWR_c_1213_n 0.00314961f $X=4.275 $Y=2.045 $X2=0
+ $Y2=0
cc_627 N_A_561_463#_c_880_n N_VPWR_c_1209_n 0.00397076f $X=4.275 $Y=2.045 $X2=0
+ $Y2=0
cc_628 N_A_561_463#_c_880_n N_VPWR_c_1222_n 0.00247808f $X=4.275 $Y=2.045 $X2=0
+ $Y2=0
cc_629 N_A_561_463#_c_874_n N_A_454_503#_c_1308_n 0.0500398f $X=2.845 $Y=2.285
+ $X2=0 $Y2=0
cc_630 N_A_561_463#_c_876_n N_A_454_503#_c_1308_n 0.0143225f $X=2.93 $Y=1.495
+ $X2=0 $Y2=0
cc_631 N_A_561_463#_c_877_n N_A_454_503#_c_1308_n 0.00504133f $X=3.325 $Y=0.78
+ $X2=0 $Y2=0
cc_632 N_A_561_463#_c_884_n N_A_454_503#_c_1308_n 0.0259474f $X=3.12 $Y=2.455
+ $X2=0 $Y2=0
cc_633 N_A_561_463#_c_875_n N_A_454_503#_c_1310_n 0.00331755f $X=3.155 $Y=1.495
+ $X2=0 $Y2=0
cc_634 N_A_561_463#_c_876_n N_A_454_503#_c_1310_n 0.014132f $X=2.93 $Y=1.495
+ $X2=0 $Y2=0
cc_635 N_A_561_463#_c_877_n N_A_454_503#_c_1310_n 0.0131425f $X=3.325 $Y=0.78
+ $X2=0 $Y2=0
cc_636 N_A_561_463#_M1004_g N_VGND_c_1371_n 0.00161104f $X=4.62 $Y=0.65 $X2=0
+ $Y2=0
cc_637 N_A_561_463#_M1004_g N_VGND_c_1374_n 0.00275597f $X=4.62 $Y=0.65 $X2=0
+ $Y2=0
cc_638 N_A_561_463#_M1004_g N_VGND_c_1381_n 0.00544287f $X=4.62 $Y=0.65 $X2=0
+ $Y2=0
cc_639 N_A_1210_314#_M1020_g N_A_1011_424#_c_1107_n 0.00439113f $X=6.18 $Y=0.83
+ $X2=0 $Y2=0
cc_640 N_A_1210_314#_c_992_n N_A_1011_424#_c_1107_n 0.0195388f $X=7.655 $Y=1.765
+ $X2=0 $Y2=0
cc_641 N_A_1210_314#_M1009_g N_A_1011_424#_c_1107_n 2.60463e-19 $X=7.665 $Y=0.74
+ $X2=0 $Y2=0
cc_642 N_A_1210_314#_c_1006_n N_A_1011_424#_c_1107_n 0.00124453f $X=7.375
+ $Y=1.775 $X2=0 $Y2=0
cc_643 N_A_1210_314#_c_995_n N_A_1011_424#_c_1107_n 0.00135071f $X=7.375
+ $Y=0.935 $X2=0 $Y2=0
cc_644 N_A_1210_314#_c_996_n N_A_1011_424#_c_1107_n 0.00383565f $X=7.04 $Y=0.935
+ $X2=0 $Y2=0
cc_645 N_A_1210_314#_c_1009_n N_A_1011_424#_c_1107_n 0.00314491f $X=6.885
+ $Y=1.775 $X2=0 $Y2=0
cc_646 N_A_1210_314#_c_1000_n N_A_1011_424#_c_1107_n 0.00266191f $X=7.555
+ $Y=1.35 $X2=0 $Y2=0
cc_647 N_A_1210_314#_c_997_n N_A_1011_424#_c_1108_n 5.77296e-19 $X=6.215
+ $Y=1.735 $X2=0 $Y2=0
cc_648 N_A_1210_314#_c_998_n N_A_1011_424#_c_1108_n 0.00110332f $X=6.215
+ $Y=1.735 $X2=0 $Y2=0
cc_649 N_A_1210_314#_c_999_n N_A_1011_424#_c_1108_n 0.00266191f $X=7.62 $Y=1.515
+ $X2=0 $Y2=0
cc_650 N_A_1210_314#_c_992_n N_A_1011_424#_c_1116_n 0.0221556f $X=7.655 $Y=1.765
+ $X2=0 $Y2=0
cc_651 N_A_1210_314#_c_1003_n N_A_1011_424#_c_1116_n 0.00434093f $X=6.215
+ $Y=2.075 $X2=0 $Y2=0
cc_652 N_A_1210_314#_c_1005_n N_A_1011_424#_c_1116_n 0.00869272f $X=6.925
+ $Y=1.985 $X2=0 $Y2=0
cc_653 N_A_1210_314#_c_1006_n N_A_1011_424#_c_1116_n 0.0166471f $X=7.375
+ $Y=1.775 $X2=0 $Y2=0
cc_654 N_A_1210_314#_c_999_n N_A_1011_424#_c_1116_n 2.22718e-19 $X=7.62 $Y=1.515
+ $X2=0 $Y2=0
cc_655 N_A_1210_314#_M1009_g N_A_1011_424#_M1007_g 0.022122f $X=7.665 $Y=0.74
+ $X2=0 $Y2=0
cc_656 N_A_1210_314#_c_994_n N_A_1011_424#_M1007_g 0.00216784f $X=6.955 $Y=0.645
+ $X2=0 $Y2=0
cc_657 N_A_1210_314#_c_995_n N_A_1011_424#_M1007_g 0.0136415f $X=7.375 $Y=0.935
+ $X2=0 $Y2=0
cc_658 N_A_1210_314#_c_1000_n N_A_1011_424#_M1007_g 0.00496447f $X=7.555 $Y=1.35
+ $X2=0 $Y2=0
cc_659 N_A_1210_314#_M1020_g N_A_1011_424#_c_1123_n 8.58394e-19 $X=6.18 $Y=0.83
+ $X2=0 $Y2=0
cc_660 N_A_1210_314#_c_1003_n N_A_1011_424#_c_1118_n 6.02883e-19 $X=6.215
+ $Y=2.075 $X2=0 $Y2=0
cc_661 N_A_1210_314#_c_997_n N_A_1011_424#_c_1118_n 0.0113488f $X=6.215 $Y=1.735
+ $X2=0 $Y2=0
cc_662 N_A_1210_314#_M1020_g N_A_1011_424#_c_1110_n 0.00131381f $X=6.18 $Y=0.83
+ $X2=0 $Y2=0
cc_663 N_A_1210_314#_M1020_g N_A_1011_424#_c_1111_n 0.00103566f $X=6.18 $Y=0.83
+ $X2=0 $Y2=0
cc_664 N_A_1210_314#_c_997_n N_A_1011_424#_c_1111_n 0.00789854f $X=6.215
+ $Y=1.735 $X2=0 $Y2=0
cc_665 N_A_1210_314#_M1020_g N_A_1011_424#_c_1113_n 7.77493e-19 $X=6.18 $Y=0.83
+ $X2=0 $Y2=0
cc_666 N_A_1210_314#_c_1006_n N_A_1011_424#_c_1113_n 0.014075f $X=7.375 $Y=1.775
+ $X2=0 $Y2=0
cc_667 N_A_1210_314#_c_995_n N_A_1011_424#_c_1113_n 0.0119514f $X=7.375 $Y=0.935
+ $X2=0 $Y2=0
cc_668 N_A_1210_314#_c_996_n N_A_1011_424#_c_1113_n 0.013898f $X=7.04 $Y=0.935
+ $X2=0 $Y2=0
cc_669 N_A_1210_314#_c_1009_n N_A_1011_424#_c_1113_n 0.011385f $X=6.885 $Y=1.775
+ $X2=0 $Y2=0
cc_670 N_A_1210_314#_c_1000_n N_A_1011_424#_c_1113_n 0.0262494f $X=7.555 $Y=1.35
+ $X2=0 $Y2=0
cc_671 N_A_1210_314#_M1020_g N_A_1011_424#_c_1114_n 0.0154848f $X=6.18 $Y=0.83
+ $X2=0 $Y2=0
cc_672 N_A_1210_314#_c_1004_n N_A_1011_424#_c_1114_n 0.0197016f $X=6.76 $Y=1.775
+ $X2=0 $Y2=0
cc_673 N_A_1210_314#_c_996_n N_A_1011_424#_c_1114_n 0.00614577f $X=7.04 $Y=0.935
+ $X2=0 $Y2=0
cc_674 N_A_1210_314#_c_997_n N_A_1011_424#_c_1114_n 0.02578f $X=6.215 $Y=1.735
+ $X2=0 $Y2=0
cc_675 N_A_1210_314#_c_998_n N_A_1011_424#_c_1114_n 0.00125303f $X=6.215
+ $Y=1.735 $X2=0 $Y2=0
cc_676 N_A_1210_314#_c_1009_n N_A_1011_424#_c_1114_n 0.0066671f $X=6.885
+ $Y=1.775 $X2=0 $Y2=0
cc_677 N_A_1210_314#_c_1006_n N_VPWR_M1008_d 0.00103504f $X=7.375 $Y=1.775 $X2=0
+ $Y2=0
cc_678 N_A_1210_314#_c_999_n N_VPWR_M1008_d 0.0016724f $X=7.62 $Y=1.515 $X2=0
+ $Y2=0
cc_679 N_A_1210_314#_c_1001_n N_VPWR_c_1211_n 0.0124028f $X=6.14 $Y=2.465 $X2=0
+ $Y2=0
cc_680 N_A_1210_314#_c_1003_n N_VPWR_c_1211_n 0.00160209f $X=6.215 $Y=2.075
+ $X2=0 $Y2=0
cc_681 N_A_1210_314#_c_1004_n N_VPWR_c_1211_n 0.004853f $X=6.76 $Y=1.775 $X2=0
+ $Y2=0
cc_682 N_A_1210_314#_c_1005_n N_VPWR_c_1211_n 0.0118856f $X=6.925 $Y=1.985 $X2=0
+ $Y2=0
cc_683 N_A_1210_314#_c_997_n N_VPWR_c_1211_n 0.0108319f $X=6.215 $Y=1.735 $X2=0
+ $Y2=0
cc_684 N_A_1210_314#_c_992_n N_VPWR_c_1212_n 0.0126023f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_685 N_A_1210_314#_c_1005_n N_VPWR_c_1212_n 0.0449538f $X=6.925 $Y=1.985 $X2=0
+ $Y2=0
cc_686 N_A_1210_314#_c_1006_n N_VPWR_c_1212_n 0.00859068f $X=7.375 $Y=1.775
+ $X2=0 $Y2=0
cc_687 N_A_1210_314#_c_999_n N_VPWR_c_1212_n 0.0132538f $X=7.62 $Y=1.515 $X2=0
+ $Y2=0
cc_688 N_A_1210_314#_c_1001_n N_VPWR_c_1213_n 0.00413917f $X=6.14 $Y=2.465 $X2=0
+ $Y2=0
cc_689 N_A_1210_314#_c_1005_n N_VPWR_c_1217_n 0.00507497f $X=6.925 $Y=1.985
+ $X2=0 $Y2=0
cc_690 N_A_1210_314#_c_992_n N_VPWR_c_1218_n 0.00445602f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_691 N_A_1210_314#_c_1001_n N_VPWR_c_1209_n 0.0081916f $X=6.14 $Y=2.465 $X2=0
+ $Y2=0
cc_692 N_A_1210_314#_c_992_n N_VPWR_c_1209_n 0.00865325f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_693 N_A_1210_314#_c_1003_n N_VPWR_c_1209_n 3.7828e-19 $X=6.215 $Y=2.075 $X2=0
+ $Y2=0
cc_694 N_A_1210_314#_c_1005_n N_VPWR_c_1209_n 0.00755367f $X=6.925 $Y=1.985
+ $X2=0 $Y2=0
cc_695 N_A_1210_314#_c_992_n N_Q_c_1346_n 0.00803445f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_696 N_A_1210_314#_c_992_n N_Q_c_1347_n 0.00192604f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_697 N_A_1210_314#_c_999_n N_Q_c_1347_n 0.00111741f $X=7.62 $Y=1.515 $X2=0
+ $Y2=0
cc_698 N_A_1210_314#_c_992_n N_Q_c_1343_n 0.0136308f $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_699 N_A_1210_314#_M1009_g N_Q_c_1343_n 0.00360849f $X=7.665 $Y=0.74 $X2=0
+ $Y2=0
cc_700 N_A_1210_314#_c_999_n N_Q_c_1343_n 0.0380678f $X=7.62 $Y=1.515 $X2=0
+ $Y2=0
cc_701 N_A_1210_314#_c_1000_n N_Q_c_1343_n 0.00756951f $X=7.555 $Y=1.35 $X2=0
+ $Y2=0
cc_702 N_A_1210_314#_M1009_g Q 0.009724f $X=7.665 $Y=0.74 $X2=0 $Y2=0
cc_703 N_A_1210_314#_c_992_n Q 0.00190025f $X=7.655 $Y=1.765 $X2=0 $Y2=0
cc_704 N_A_1210_314#_M1009_g Q 0.00281925f $X=7.665 $Y=0.74 $X2=0 $Y2=0
cc_705 N_A_1210_314#_c_999_n Q 0.00121064f $X=7.62 $Y=1.515 $X2=0 $Y2=0
cc_706 N_A_1210_314#_c_1000_n Q 0.00489765f $X=7.555 $Y=1.35 $X2=0 $Y2=0
cc_707 N_A_1210_314#_c_995_n N_VGND_M1007_d 0.00417906f $X=7.375 $Y=0.935 $X2=0
+ $Y2=0
cc_708 N_A_1210_314#_c_1000_n N_VGND_M1007_d 0.00153963f $X=7.555 $Y=1.35 $X2=0
+ $Y2=0
cc_709 N_A_1210_314#_M1020_g N_VGND_c_1372_n 0.0138099f $X=6.18 $Y=0.83 $X2=0
+ $Y2=0
cc_710 N_A_1210_314#_c_994_n N_VGND_c_1372_n 0.0329832f $X=6.955 $Y=0.645 $X2=0
+ $Y2=0
cc_711 N_A_1210_314#_c_996_n N_VGND_c_1372_n 0.0121616f $X=7.04 $Y=0.935 $X2=0
+ $Y2=0
cc_712 N_A_1210_314#_c_992_n N_VGND_c_1373_n 2.33587e-19 $X=7.655 $Y=1.765 $X2=0
+ $Y2=0
cc_713 N_A_1210_314#_M1009_g N_VGND_c_1373_n 0.00318537f $X=7.665 $Y=0.74 $X2=0
+ $Y2=0
cc_714 N_A_1210_314#_c_994_n N_VGND_c_1373_n 0.0124717f $X=6.955 $Y=0.645 $X2=0
+ $Y2=0
cc_715 N_A_1210_314#_c_995_n N_VGND_c_1373_n 0.0214421f $X=7.375 $Y=0.935 $X2=0
+ $Y2=0
cc_716 N_A_1210_314#_M1020_g N_VGND_c_1374_n 0.00347405f $X=6.18 $Y=0.83 $X2=0
+ $Y2=0
cc_717 N_A_1210_314#_c_994_n N_VGND_c_1379_n 0.011054f $X=6.955 $Y=0.645 $X2=0
+ $Y2=0
cc_718 N_A_1210_314#_M1009_g N_VGND_c_1380_n 0.00434272f $X=7.665 $Y=0.74 $X2=0
+ $Y2=0
cc_719 N_A_1210_314#_M1020_g N_VGND_c_1381_n 0.00395485f $X=6.18 $Y=0.83 $X2=0
+ $Y2=0
cc_720 N_A_1210_314#_M1009_g N_VGND_c_1381_n 0.00824612f $X=7.665 $Y=0.74 $X2=0
+ $Y2=0
cc_721 N_A_1210_314#_c_994_n N_VGND_c_1381_n 0.00915483f $X=6.955 $Y=0.645 $X2=0
+ $Y2=0
cc_722 N_A_1210_314#_c_995_n N_VGND_c_1381_n 0.0067624f $X=7.375 $Y=0.935 $X2=0
+ $Y2=0
cc_723 N_A_1011_424#_c_1116_n N_VPWR_c_1211_n 0.003066f $X=7.15 $Y=1.765 $X2=0
+ $Y2=0
cc_724 N_A_1011_424#_c_1116_n N_VPWR_c_1212_n 0.0141077f $X=7.15 $Y=1.765 $X2=0
+ $Y2=0
cc_725 N_A_1011_424#_c_1116_n N_VPWR_c_1217_n 0.00361294f $X=7.15 $Y=1.765 $X2=0
+ $Y2=0
cc_726 N_A_1011_424#_c_1116_n N_VPWR_c_1209_n 0.00419404f $X=7.15 $Y=1.765 $X2=0
+ $Y2=0
cc_727 N_A_1011_424#_c_1116_n N_Q_c_1347_n 2.44869e-19 $X=7.15 $Y=1.765 $X2=0
+ $Y2=0
cc_728 N_A_1011_424#_M1007_g Q 6.76541e-19 $X=7.17 $Y=0.645 $X2=0 $Y2=0
cc_729 N_A_1011_424#_M1007_g N_VGND_c_1372_n 0.00428687f $X=7.17 $Y=0.645 $X2=0
+ $Y2=0
cc_730 N_A_1011_424#_c_1123_n N_VGND_c_1372_n 0.00968609f $X=5.65 $Y=0.855 $X2=0
+ $Y2=0
cc_731 N_A_1011_424#_c_1110_n N_VGND_c_1372_n 0.00279148f $X=5.735 $Y=1.23 $X2=0
+ $Y2=0
cc_732 N_A_1011_424#_c_1114_n N_VGND_c_1372_n 0.0275041f $X=6.875 $Y=1.355 $X2=0
+ $Y2=0
cc_733 N_A_1011_424#_M1007_g N_VGND_c_1373_n 0.00828491f $X=7.17 $Y=0.645 $X2=0
+ $Y2=0
cc_734 N_A_1011_424#_M1007_g N_VGND_c_1379_n 0.00383152f $X=7.17 $Y=0.645 $X2=0
+ $Y2=0
cc_735 N_A_1011_424#_M1007_g N_VGND_c_1381_n 0.00391057f $X=7.17 $Y=0.645 $X2=0
+ $Y2=0
cc_736 N_VPWR_c_1218_n N_Q_c_1346_n 0.0159324f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_737 N_VPWR_c_1209_n N_Q_c_1346_n 0.0131546f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_738 N_VPWR_c_1212_n N_Q_c_1347_n 0.036031f $X=7.375 $Y=2.135 $X2=0 $Y2=0
cc_739 Q N_VGND_c_1373_n 0.0127401f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_740 Q N_VGND_c_1380_n 0.0159025f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_741 Q N_VGND_c_1381_n 0.0131064f $X=7.835 $Y=0.47 $X2=0 $Y2=0
