# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ls__dlymetal6s2s_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ls__dlymetal6s2s_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.355000 0.555000 1.765000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.835000 1.380000 3.075000 ;
        RECT 1.090000 0.255000 1.380000 1.075000 ;
        RECT 1.210000 1.075000 1.380000 1.315000 ;
        RECT 1.210000 1.315000 1.995000 1.605000 ;
        RECT 1.210000 1.605000 1.380000 1.835000 ;
      LAYER mcon ;
        RECT 1.115000 1.950000 1.285000 2.120000 ;
      LAYER met1 ;
        RECT 0.965000 1.920000 1.345000 2.320000 ;
        RECT 0.965000 2.320000 4.210000 2.490000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.800000 0.085000 ;
        RECT 0.590000  0.085000 0.920000 0.805000 ;
        RECT 2.030000  0.085000 2.360000 0.805000 ;
        RECT 3.470000  0.085000 3.800000 0.805000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 4.800000 3.415000 ;
        RECT 0.590000 2.310000 0.885000 3.245000 ;
        RECT 2.100000 2.310000 2.395000 3.245000 ;
        RECT 3.585000 2.310000 3.880000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.100000 0.700000 0.395000 0.975000 ;
      RECT 0.100000 0.975000 0.895000 1.145000 ;
      RECT 0.100000 1.935000 0.895000 2.140000 ;
      RECT 0.100000 2.140000 0.430000 2.225000 ;
      RECT 0.725000 1.145000 0.895000 1.275000 ;
      RECT 0.725000 1.275000 1.040000 1.605000 ;
      RECT 0.725000 1.605000 0.895000 1.935000 ;
      RECT 1.550000 0.700000 1.835000 0.975000 ;
      RECT 1.550000 0.975000 2.335000 1.145000 ;
      RECT 1.550000 1.895000 2.335000 2.140000 ;
      RECT 1.550000 2.140000 1.870000 2.225000 ;
      RECT 2.165000 1.145000 2.335000 1.275000 ;
      RECT 2.165000 1.275000 2.525000 1.605000 ;
      RECT 2.165000 1.605000 2.335000 1.895000 ;
      RECT 2.505000 1.835000 2.865000 2.160000 ;
      RECT 2.530000 0.255000 2.865000 1.075000 ;
      RECT 2.565000 2.160000 2.865000 3.075000 ;
      RECT 2.695000 1.075000 2.865000 1.315000 ;
      RECT 2.695000 1.315000 3.435000 1.605000 ;
      RECT 2.695000 1.605000 2.865000 1.835000 ;
      RECT 3.060000 0.700000 3.275000 0.975000 ;
      RECT 3.060000 0.975000 3.775000 1.145000 ;
      RECT 3.070000 1.895000 3.805000 2.140000 ;
      RECT 3.070000 2.140000 3.400000 2.225000 ;
      RECT 3.605000 1.145000 3.775000 1.275000 ;
      RECT 3.605000 1.275000 4.010000 1.605000 ;
      RECT 3.605000 1.605000 3.805000 1.895000 ;
      RECT 3.970000 0.255000 4.350000 1.075000 ;
      RECT 3.975000 1.835000 4.350000 2.160000 ;
      RECT 4.050000 2.160000 4.350000 3.075000 ;
      RECT 4.180000 1.075000 4.350000 1.835000 ;
    LAYER mcon ;
      RECT 2.555000 1.950000 2.725000 2.120000 ;
      RECT 3.995000 1.950000 4.165000 2.120000 ;
    LAYER met1 ;
      RECT 2.405000 1.920000 2.785000 2.150000 ;
      RECT 3.845000 1.920000 4.225000 2.150000 ;
  END
END sky130_fd_sc_ls__dlymetal6s2s_1
