* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_409_81# a_27_74# a_512_464# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_512_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_835_98# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_1747_74# a_1034_392# a_1969_489# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR a_1747_74# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X5 a_409_81# a_835_98# a_1234_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_2513_424# a_1747_74# VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X7 VGND a_1234_119# a_1367_93# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 a_2124_74# a_1747_74# a_2008_48# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_312_81# D a_409_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR a_835_98# a_1034_392# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_225_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR a_1234_119# a_1367_93# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_2008_48# a_1747_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 VPWR RESET_B a_1234_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 VGND a_835_98# a_1034_392# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 a_1234_119# a_835_98# a_1332_457# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_225_81# a_27_74# a_312_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_2513_424# a_1747_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X19 a_1969_489# a_2008_48# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VGND RESET_B a_2124_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_338_464# D a_409_81# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 a_1367_93# a_1034_392# a_1747_74# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X23 VGND a_2513_424# Q VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X24 a_1367_93# a_835_98# a_1747_74# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 VGND a_1747_74# Q_N VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X27 VPWR RESET_B a_409_81# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X28 a_1320_119# a_1367_93# a_1397_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_409_81# SCE a_545_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 VPWR a_2513_424# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X32 VPWR RESET_B a_2008_48# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 a_1747_74# a_835_98# a_1966_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_1332_457# a_1367_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X35 a_835_98# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X36 a_1234_119# a_1034_392# a_1320_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 VPWR SCE a_338_464# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X38 a_409_81# a_1034_392# a_1234_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X39 a_545_81# SCD a_225_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 a_1397_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 a_1966_74# a_2008_48# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
