* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfxtp_1 CLK D VGND VNB VPB VPWR Q
M1000 VPWR a_713_458# a_668_503# VPB phighvt w=420000u l=150000u
+  ad=1.50923e+12p pd=1.272e+07u as=1.008e+11p ps=1.32e+06u
M1001 a_206_368# a_27_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.553e+11p pd=2.17e+06u as=1.2645e+12p ps=1.059e+07u
M1002 a_1118_508# a_206_368# a_1011_424# VPB phighvt w=420000u l=150000u
+  ad=1.995e+11p pd=1.79e+06u as=2.856e+11p ps=2.45e+06u
M1003 VPWR a_1210_314# a_1118_508# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_713_458# a_561_463# VGND VNB nshort w=550000u l=150000u
+  ad=2.18125e+11p pd=2.05e+06u as=0p ps=0u
M1005 a_1011_424# a_206_368# a_713_458# VNB nshort w=550000u l=150000u
+  ad=2.362e+11p pd=2.07e+06u as=0p ps=0u
M1006 a_454_503# D VGND VNB nshort w=420000u l=150000u
+  ad=3.1125e+11p pd=2.43e+06u as=0p ps=0u
M1007 VGND a_1011_424# a_1210_314# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1008 VPWR a_1011_424# a_1210_314# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1009 Q a_1210_314# VGND VNB nshort w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1010 Q a_1210_314# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1011 VGND a_713_458# a_731_101# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1012 a_454_503# D VPWR VPB phighvt w=420000u l=150000u
+  ad=1.967e+11p pd=2.01e+06u as=0p ps=0u
M1013 a_668_503# a_27_74# a_561_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.967e+11p ps=2.01e+06u
M1014 VPWR CLK a_27_74# VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1015 a_206_368# a_27_74# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1016 a_731_101# a_206_368# a_561_463# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.575e+11p ps=1.73e+06u
M1017 a_561_463# a_27_74# a_454_503# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_713_458# a_561_463# VPWR VPB phighvt w=840000u l=150000u
+  ad=4.662e+11p pd=2.79e+06u as=0p ps=0u
M1019 a_1011_424# a_27_74# a_713_458# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_1210_314# a_1168_124# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1021 a_561_463# a_206_368# a_454_503# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND CLK a_27_74# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1023 a_1168_124# a_27_74# a_1011_424# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
