* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__einvn_2 A TE_B VGND VNB VPB VPWR Z
X0 Z A a_227_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VPWR TE_B a_227_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 a_231_74# a_115_464# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 VGND a_115_464# a_231_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X4 VPWR TE_B a_115_464# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_231_74# A Z VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 Z A a_231_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X7 a_227_368# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 a_227_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 VGND TE_B a_115_464# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
