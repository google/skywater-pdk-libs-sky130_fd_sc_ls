* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__clkbuf_2 A VGND VNB VPB VPWR X
M1000 a_43_192# A VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.528e+11p pd=2.87e+06u as=6.552e+11p ps=5.65e+06u
M1001 a_43_192# A VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=2.667e+11p ps=2.95e+06u
M1002 X a_43_192# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1003 VPWR a_43_192# X VPB phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_43_192# VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1005 VGND a_43_192# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
