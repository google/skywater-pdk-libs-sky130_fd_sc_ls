* File: sky130_fd_sc_ls__o32a_1.pxi.spice
* Created: Fri Aug 28 13:53:58 2020
* 
x_PM_SKY130_FD_SC_LS__O32A_1%A_83_264# N_A_83_264#_M1002_d N_A_83_264#_M1011_d
+ N_A_83_264#_c_68_n N_A_83_264#_M1007_g N_A_83_264#_M1004_g N_A_83_264#_c_70_n
+ N_A_83_264#_c_80_p N_A_83_264#_c_128_p N_A_83_264#_c_76_n N_A_83_264#_c_97_p
+ N_A_83_264#_c_71_n N_A_83_264#_c_72_n N_A_83_264#_c_73_n N_A_83_264#_c_93_p
+ PM_SKY130_FD_SC_LS__O32A_1%A_83_264#
x_PM_SKY130_FD_SC_LS__O32A_1%A1 N_A1_c_150_n N_A1_M1010_g N_A1_M1009_g A1
+ N_A1_c_152_n PM_SKY130_FD_SC_LS__O32A_1%A1
x_PM_SKY130_FD_SC_LS__O32A_1%A2 N_A2_c_185_n N_A2_M1006_g N_A2_M1001_g A2
+ N_A2_c_187_n PM_SKY130_FD_SC_LS__O32A_1%A2
x_PM_SKY130_FD_SC_LS__O32A_1%A3 N_A3_c_215_n N_A3_M1011_g N_A3_M1005_g A3
+ N_A3_c_217_n PM_SKY130_FD_SC_LS__O32A_1%A3
x_PM_SKY130_FD_SC_LS__O32A_1%B2 N_B2_c_246_n N_B2_M1003_g N_B2_M1002_g B2
+ N_B2_c_248_n PM_SKY130_FD_SC_LS__O32A_1%B2
x_PM_SKY130_FD_SC_LS__O32A_1%B1 N_B1_c_280_n N_B1_c_285_n N_B1_M1008_g
+ N_B1_M1000_g B1 B1 N_B1_c_283_n PM_SKY130_FD_SC_LS__O32A_1%B1
x_PM_SKY130_FD_SC_LS__O32A_1%X N_X_M1004_s N_X_M1007_s N_X_c_315_n N_X_c_316_n
+ N_X_c_312_n X X N_X_c_313_n X PM_SKY130_FD_SC_LS__O32A_1%X
x_PM_SKY130_FD_SC_LS__O32A_1%VPWR N_VPWR_M1007_d N_VPWR_M1008_d N_VPWR_c_340_n
+ N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n N_VPWR_c_344_n VPWR
+ N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n N_VPWR_c_339_n
+ PM_SKY130_FD_SC_LS__O32A_1%VPWR
x_PM_SKY130_FD_SC_LS__O32A_1%VGND N_VGND_M1004_d N_VGND_M1001_d N_VGND_c_383_n
+ N_VGND_c_384_n N_VGND_c_385_n N_VGND_c_386_n N_VGND_c_387_n N_VGND_c_388_n
+ VGND N_VGND_c_389_n N_VGND_c_390_n PM_SKY130_FD_SC_LS__O32A_1%VGND
x_PM_SKY130_FD_SC_LS__O32A_1%A_251_74# N_A_251_74#_M1009_d N_A_251_74#_M1005_d
+ N_A_251_74#_M1000_d N_A_251_74#_c_427_n N_A_251_74#_c_428_n
+ N_A_251_74#_c_429_n N_A_251_74#_c_430_n N_A_251_74#_c_448_n
+ N_A_251_74#_c_431_n N_A_251_74#_c_432_n PM_SKY130_FD_SC_LS__O32A_1%A_251_74#
cc_1 VNB N_A_83_264#_c_68_n 0.0343522f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_A_83_264#_M1004_g 0.03041f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_3 VNB N_A_83_264#_c_70_n 2.45937e-19 $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.95
cc_4 VNB N_A_83_264#_c_71_n 0.00753812f $X=-0.19 $Y=-0.245 $X2=3.15 $Y2=1.18
cc_5 VNB N_A_83_264#_c_72_n 0.0036728f $X=-0.19 $Y=-0.245 $X2=3.15 $Y2=1.95
cc_6 VNB N_A_83_264#_c_73_n 0.0027277f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.485
cc_7 VNB N_A1_c_150_n 0.0243054f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=0.37
cc_8 VNB N_A1_M1009_g 0.0314409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A1_c_152_n 0.00547709f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_10 VNB N_A2_c_185_n 0.0262312f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=0.37
cc_11 VNB N_A2_M1001_g 0.0305392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_187_n 0.00165774f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_13 VNB N_A3_c_215_n 0.0262279f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=0.37
cc_14 VNB N_A3_M1005_g 0.0316956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A3_c_217_n 0.00165645f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_16 VNB N_B2_c_246_n 0.0249237f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=0.37
cc_17 VNB N_B2_M1002_g 0.0326134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B2_c_248_n 0.0051357f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_19 VNB N_B1_c_280_n 0.00797545f $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=1.84
cc_20 VNB N_B1_M1000_g 0.0294724f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_21 VNB B1 0.0119477f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.32
cc_22 VNB N_B1_c_283_n 0.067073f $X=-0.19 $Y=-0.245 $X2=2.4 $Y2=2.12
cc_23 VNB N_X_c_312_n 0.0251021f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.95
cc_24 VNB N_X_c_313_n 0.0283371f $X=-0.19 $Y=-0.245 $X2=2.595 $Y2=2.035
cc_25 VNB X 0.0180876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_339_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_383_n 0.0109103f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_28 VNB N_VGND_c_384_n 0.00895062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_385_n 0.0216783f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=2.035
cc_30 VNB N_VGND_c_386_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.035
cc_31 VNB N_VGND_c_387_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=2.4 $Y2=2.375
cc_32 VNB N_VGND_c_388_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=2.375
cc_33 VNB N_VGND_c_389_n 0.0474473f $X=-0.19 $Y=-0.245 $X2=2.982 $Y2=0.865
cc_34 VNB N_VGND_c_390_n 0.23222f $X=-0.19 $Y=-0.245 $X2=2.975 $Y2=0.865
cc_35 VNB N_A_251_74#_c_427_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_36 VNB N_A_251_74#_c_428_n 0.0247434f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.65
cc_37 VNB N_A_251_74#_c_429_n 0.00810708f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.95
cc_38 VNB N_A_251_74#_c_430_n 0.00257219f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=2.035
cc_39 VNB N_A_251_74#_c_431_n 0.00456757f $X=-0.19 $Y=-0.245 $X2=2.4 $Y2=2.12
cc_40 VNB N_A_251_74#_c_432_n 0.0049404f $X=-0.19 $Y=-0.245 $X2=3.15 $Y2=1.95
cc_41 VPB N_A_83_264#_c_68_n 0.0297798f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_42 VPB N_A_83_264#_c_70_n 0.00284593f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.95
cc_43 VPB N_A_83_264#_c_76_n 0.00457874f $X=-0.19 $Y=1.66 $X2=2.395 $Y2=2.375
cc_44 VPB N_A_83_264#_c_72_n 0.00142167f $X=-0.19 $Y=1.66 $X2=3.15 $Y2=1.95
cc_45 VPB N_A1_c_150_n 0.0271668f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=0.37
cc_46 VPB N_A1_c_152_n 0.00335979f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.74
cc_47 VPB N_A2_c_185_n 0.0267782f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=0.37
cc_48 VPB N_A2_c_187_n 0.00241789f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.74
cc_49 VPB N_A3_c_215_n 0.0280001f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=0.37
cc_50 VPB N_A3_c_217_n 0.00238456f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.74
cc_51 VPB N_B2_c_246_n 0.027721f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=0.37
cc_52 VPB N_B2_c_248_n 0.00336148f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.74
cc_53 VPB N_B1_c_280_n 7.49372e-19 $X=-0.19 $Y=1.66 $X2=2.2 $Y2=1.84
cc_54 VPB N_B1_c_285_n 0.0250515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB B1 0.011961f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.32
cc_56 VPB N_X_c_315_n 0.041687f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.74
cc_57 VPB N_X_c_316_n 0.0138434f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.65
cc_58 VPB N_X_c_312_n 0.0075617f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.95
cc_59 VPB N_VPWR_c_340_n 0.0143226f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_60 VPB N_VPWR_c_341_n 0.00626527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_342_n 0.0145833f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.65
cc_62 VPB N_VPWR_c_343_n 0.0347679f $X=-0.19 $Y=1.66 $X2=2.205 $Y2=2.035
cc_63 VPB N_VPWR_c_344_n 0.0117986f $X=-0.19 $Y=1.66 $X2=2.4 $Y2=2.375
cc_64 VPB N_VPWR_c_345_n 0.0189171f $X=-0.19 $Y=1.66 $X2=3.15 $Y2=1.18
cc_65 VPB N_VPWR_c_346_n 0.0729976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_347_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_339_n 0.119735f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 N_A_83_264#_c_68_n N_A1_c_150_n 0.0404013f $X=0.505 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_69 N_A_83_264#_c_70_n N_A1_c_150_n 0.00376784f $X=0.7 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_70 N_A_83_264#_c_80_p N_A1_c_150_n 0.0163635f $X=2.205 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_71 N_A_83_264#_c_73_n N_A1_c_150_n 0.00170039f $X=0.7 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_72 N_A_83_264#_c_68_n N_A1_M1009_g 8.96112e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A_83_264#_M1004_g N_A1_M1009_g 0.023959f $X=0.61 $Y=0.74 $X2=0 $Y2=0
cc_74 N_A_83_264#_c_73_n N_A1_M1009_g 5.98792e-19 $X=0.7 $Y=1.485 $X2=0 $Y2=0
cc_75 N_A_83_264#_c_68_n N_A1_c_152_n 3.43727e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A_83_264#_c_70_n N_A1_c_152_n 0.0102525f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_77 N_A_83_264#_c_80_p N_A1_c_152_n 0.023487f $X=2.205 $Y=2.035 $X2=0 $Y2=0
cc_78 N_A_83_264#_c_73_n N_A1_c_152_n 0.0240952f $X=0.7 $Y=1.485 $X2=0 $Y2=0
cc_79 N_A_83_264#_c_80_p N_A2_c_185_n 0.0162159f $X=2.205 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_80 N_A_83_264#_c_80_p N_A2_c_187_n 0.0226548f $X=2.205 $Y=2.035 $X2=0 $Y2=0
cc_81 N_A_83_264#_c_80_p N_A3_c_215_n 0.0135074f $X=2.205 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_82 N_A_83_264#_c_76_n N_A3_c_215_n 0.0012286f $X=2.395 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_83 N_A_83_264#_c_93_p N_A3_c_215_n 8.08813e-19 $X=2.395 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_84 N_A_83_264#_c_80_p N_A3_c_217_n 0.011794f $X=2.205 $Y=2.035 $X2=0 $Y2=0
cc_85 N_A_83_264#_c_93_p N_A3_c_217_n 0.0117765f $X=2.395 $Y=2.035 $X2=0 $Y2=0
cc_86 N_A_83_264#_c_76_n N_B2_c_246_n 0.0154583f $X=2.395 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_87 N_A_83_264#_c_97_p N_B2_c_246_n 0.0144191f $X=3.065 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_88 N_A_83_264#_c_71_n N_B2_c_246_n 0.00152828f $X=3.15 $Y=1.18 $X2=-0.19
+ $Y2=-0.245
cc_89 N_A_83_264#_c_72_n N_B2_c_246_n 0.00539177f $X=3.15 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_90 N_A_83_264#_c_71_n N_B2_M1002_g 0.0135416f $X=3.15 $Y=1.18 $X2=0 $Y2=0
cc_91 N_A_83_264#_c_72_n N_B2_M1002_g 0.00313735f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_92 N_A_83_264#_c_97_p N_B2_c_248_n 0.0208442f $X=3.065 $Y=2.035 $X2=0 $Y2=0
cc_93 N_A_83_264#_c_71_n N_B2_c_248_n 0.0136544f $X=3.15 $Y=1.18 $X2=0 $Y2=0
cc_94 N_A_83_264#_c_72_n N_B2_c_248_n 0.0329498f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_95 N_A_83_264#_c_93_p N_B2_c_248_n 0.00272805f $X=2.395 $Y=2.035 $X2=0 $Y2=0
cc_96 N_A_83_264#_c_72_n N_B1_c_280_n 0.00329951f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_97 N_A_83_264#_c_76_n N_B1_c_285_n 0.00330497f $X=2.395 $Y=2.375 $X2=0 $Y2=0
cc_98 N_A_83_264#_c_97_p N_B1_c_285_n 0.00820643f $X=3.065 $Y=2.035 $X2=0 $Y2=0
cc_99 N_A_83_264#_c_72_n N_B1_c_285_n 0.0115533f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_100 N_A_83_264#_c_71_n N_B1_M1000_g 0.0197418f $X=3.15 $Y=1.18 $X2=0 $Y2=0
cc_101 N_A_83_264#_c_72_n B1 0.042784f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_102 N_A_83_264#_c_71_n N_B1_c_283_n 6.70187e-19 $X=3.15 $Y=1.18 $X2=0 $Y2=0
cc_103 N_A_83_264#_c_72_n N_B1_c_283_n 0.00900681f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_104 N_A_83_264#_c_68_n N_X_c_315_n 0.0130375f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A_83_264#_c_68_n N_X_c_316_n 0.00300223f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_106 N_A_83_264#_c_70_n N_X_c_316_n 0.00565815f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_107 N_A_83_264#_c_73_n N_X_c_316_n 0.00153915f $X=0.7 $Y=1.485 $X2=0 $Y2=0
cc_108 N_A_83_264#_c_68_n N_X_c_312_n 0.0101525f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_109 N_A_83_264#_M1004_g N_X_c_312_n 0.00424574f $X=0.61 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A_83_264#_c_70_n N_X_c_312_n 0.00535848f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_111 N_A_83_264#_c_73_n N_X_c_312_n 0.0249376f $X=0.7 $Y=1.485 $X2=0 $Y2=0
cc_112 N_A_83_264#_M1004_g N_X_c_313_n 0.0075748f $X=0.61 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A_83_264#_c_68_n X 0.00339811f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_114 N_A_83_264#_M1004_g X 0.00423703f $X=0.61 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A_83_264#_c_73_n X 0.0102842f $X=0.7 $Y=1.485 $X2=0 $Y2=0
cc_116 N_A_83_264#_c_70_n N_VPWR_M1007_d 0.00228597f $X=0.7 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_117 N_A_83_264#_c_80_p N_VPWR_M1007_d 0.0133826f $X=2.205 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_118 N_A_83_264#_c_128_p N_VPWR_M1007_d 0.00300113f $X=0.785 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_119 N_A_83_264#_c_68_n N_VPWR_c_340_n 0.0102525f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_120 N_A_83_264#_c_80_p N_VPWR_c_340_n 0.0128995f $X=2.205 $Y=2.035 $X2=0
+ $Y2=0
cc_121 N_A_83_264#_c_128_p N_VPWR_c_340_n 0.0129456f $X=0.785 $Y=2.035 $X2=0
+ $Y2=0
cc_122 N_A_83_264#_c_97_p N_VPWR_c_344_n 0.0118099f $X=3.065 $Y=2.035 $X2=0
+ $Y2=0
cc_123 N_A_83_264#_c_68_n N_VPWR_c_345_n 0.00445602f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_124 N_A_83_264#_c_76_n N_VPWR_c_346_n 0.0123062f $X=2.395 $Y=2.375 $X2=0
+ $Y2=0
cc_125 N_A_83_264#_c_68_n N_VPWR_c_339_n 0.00865213f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_126 N_A_83_264#_c_76_n N_VPWR_c_339_n 0.0134332f $X=2.395 $Y=2.375 $X2=0
+ $Y2=0
cc_127 N_A_83_264#_c_80_p A_248_368# 0.0114366f $X=2.205 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_83_264#_c_80_p A_332_368# 0.018186f $X=2.205 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_129 N_A_83_264#_c_97_p A_548_368# 0.0208204f $X=3.065 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_130 N_A_83_264#_c_72_n A_548_368# 0.00143335f $X=3.15 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_131 N_A_83_264#_c_68_n N_VGND_c_383_n 2.61167e-19 $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A_83_264#_M1004_g N_VGND_c_383_n 0.00737997f $X=0.61 $Y=0.74 $X2=0
+ $Y2=0
cc_133 N_A_83_264#_c_73_n N_VGND_c_383_n 0.00279673f $X=0.7 $Y=1.485 $X2=0 $Y2=0
cc_134 N_A_83_264#_M1004_g N_VGND_c_385_n 0.00434272f $X=0.61 $Y=0.74 $X2=0
+ $Y2=0
cc_135 N_A_83_264#_M1004_g N_VGND_c_390_n 0.00825303f $X=0.61 $Y=0.74 $X2=0
+ $Y2=0
cc_136 N_A_83_264#_c_71_n N_A_251_74#_c_428_n 0.0147887f $X=3.15 $Y=1.18 $X2=0
+ $Y2=0
cc_137 N_A_83_264#_M1004_g N_A_251_74#_c_429_n 5.42515e-19 $X=0.61 $Y=0.74 $X2=0
+ $Y2=0
cc_138 N_A_83_264#_M1002_d N_A_251_74#_c_431_n 0.00431143f $X=2.755 $Y=0.37
+ $X2=0 $Y2=0
cc_139 N_A_83_264#_c_71_n N_A_251_74#_c_431_n 0.0277999f $X=3.15 $Y=1.18 $X2=0
+ $Y2=0
cc_140 N_A1_c_150_n N_A2_c_185_n 0.0847137f $X=1.165 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_141 N_A1_c_152_n N_A2_c_185_n 0.00241815f $X=1.12 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_142 N_A1_M1009_g N_A2_M1001_g 0.0217728f $X=1.18 $Y=0.69 $X2=0 $Y2=0
cc_143 N_A1_c_150_n N_A2_c_187_n 5.31004e-19 $X=1.165 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A1_c_152_n N_A2_c_187_n 0.0328897f $X=1.12 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A1_c_150_n N_X_c_315_n 8.36183e-19 $X=1.165 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A1_M1009_g N_X_c_313_n 4.46111e-19 $X=1.18 $Y=0.69 $X2=0 $Y2=0
cc_147 N_A1_c_150_n N_VPWR_c_340_n 0.0180916f $X=1.165 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A1_c_150_n N_VPWR_c_346_n 0.0049405f $X=1.165 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A1_c_150_n N_VPWR_c_339_n 0.00508379f $X=1.165 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A1_c_150_n N_VGND_c_383_n 7.53427e-19 $X=1.165 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A1_M1009_g N_VGND_c_383_n 0.00606053f $X=1.18 $Y=0.69 $X2=0 $Y2=0
cc_152 N_A1_c_152_n N_VGND_c_383_n 0.00553853f $X=1.12 $Y=1.515 $X2=0 $Y2=0
cc_153 N_A1_M1009_g N_VGND_c_387_n 0.00434272f $X=1.18 $Y=0.69 $X2=0 $Y2=0
cc_154 N_A1_M1009_g N_VGND_c_390_n 0.0082141f $X=1.18 $Y=0.69 $X2=0 $Y2=0
cc_155 N_A1_M1009_g N_A_251_74#_c_427_n 0.00725678f $X=1.18 $Y=0.69 $X2=0 $Y2=0
cc_156 N_A1_c_150_n N_A_251_74#_c_429_n 2.37442e-19 $X=1.165 $Y=1.765 $X2=0
+ $Y2=0
cc_157 N_A1_M1009_g N_A_251_74#_c_429_n 0.0056999f $X=1.18 $Y=0.69 $X2=0 $Y2=0
cc_158 N_A1_c_152_n N_A_251_74#_c_429_n 0.00726085f $X=1.12 $Y=1.515 $X2=0 $Y2=0
cc_159 N_A2_c_185_n N_A3_c_215_n 0.0625522f $X=1.585 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_160 N_A2_c_187_n N_A3_c_215_n 0.00179181f $X=1.66 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_161 N_A2_M1001_g N_A3_M1005_g 0.0261471f $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_162 N_A2_c_185_n N_A3_c_217_n 0.00127792f $X=1.585 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A2_c_187_n N_A3_c_217_n 0.0277337f $X=1.66 $Y=1.515 $X2=0 $Y2=0
cc_164 N_A2_c_185_n N_VPWR_c_346_n 0.0049405f $X=1.585 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A2_c_185_n N_VPWR_c_339_n 0.00508379f $X=1.585 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A2_M1001_g N_VGND_c_384_n 0.00472263f $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_167 N_A2_M1001_g N_VGND_c_387_n 0.00434272f $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_168 N_A2_M1001_g N_VGND_c_390_n 0.0082141f $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_169 N_A2_M1001_g N_A_251_74#_c_427_n 0.00915605f $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_170 N_A2_c_185_n N_A_251_74#_c_428_n 9.79877e-19 $X=1.585 $Y=1.765 $X2=0
+ $Y2=0
cc_171 N_A2_M1001_g N_A_251_74#_c_428_n 0.0117933f $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_172 N_A2_c_187_n N_A_251_74#_c_428_n 0.019847f $X=1.66 $Y=1.515 $X2=0 $Y2=0
cc_173 N_A2_c_185_n N_A_251_74#_c_429_n 3.05922e-19 $X=1.585 $Y=1.765 $X2=0
+ $Y2=0
cc_174 N_A2_M1001_g N_A_251_74#_c_429_n 0.0027332f $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_175 N_A2_c_187_n N_A_251_74#_c_429_n 0.00541082f $X=1.66 $Y=1.515 $X2=0 $Y2=0
cc_176 N_A2_M1001_g N_A_251_74#_c_448_n 6.53479e-19 $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_177 N_A3_c_215_n N_B2_c_246_n 0.0304218f $X=2.125 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_178 N_A3_c_217_n N_B2_c_246_n 7.18891e-19 $X=2.2 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_179 N_A3_M1005_g N_B2_M1002_g 0.0253778f $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_180 N_A3_c_215_n N_B2_c_248_n 0.00214276f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_181 N_A3_c_217_n N_B2_c_248_n 0.0346782f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_182 N_A3_c_215_n N_VPWR_c_346_n 0.0049405f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_183 N_A3_c_215_n N_VPWR_c_339_n 0.00508379f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A3_M1005_g N_VGND_c_384_n 0.00590558f $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_185 N_A3_M1005_g N_VGND_c_389_n 0.00432912f $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_186 N_A3_M1005_g N_VGND_c_390_n 0.00818188f $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_187 N_A3_M1005_g N_A_251_74#_c_427_n 6.8749e-19 $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_188 N_A3_c_215_n N_A_251_74#_c_428_n 0.00134355f $X=2.125 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_A3_M1005_g N_A_251_74#_c_428_n 0.0145861f $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_190 N_A3_c_217_n N_A_251_74#_c_428_n 0.0259036f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_191 N_A3_M1005_g N_A_251_74#_c_430_n 0.00250516f $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_192 N_A3_M1005_g N_A_251_74#_c_448_n 0.00693236f $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_193 N_B2_c_246_n N_B1_c_285_n 0.030825f $X=2.665 $Y=1.765 $X2=0 $Y2=0
cc_194 N_B2_c_248_n N_B1_c_285_n 3.04709e-19 $X=2.74 $Y=1.515 $X2=0 $Y2=0
cc_195 N_B2_M1002_g N_B1_M1000_g 0.0231667f $X=2.68 $Y=0.69 $X2=0 $Y2=0
cc_196 N_B2_c_246_n N_B1_c_283_n 0.0152021f $X=2.665 $Y=1.765 $X2=0 $Y2=0
cc_197 N_B2_M1002_g N_B1_c_283_n 0.00411837f $X=2.68 $Y=0.69 $X2=0 $Y2=0
cc_198 N_B2_c_248_n N_B1_c_283_n 3.40711e-19 $X=2.74 $Y=1.515 $X2=0 $Y2=0
cc_199 N_B2_c_246_n N_VPWR_c_341_n 0.00301068f $X=2.665 $Y=1.765 $X2=0 $Y2=0
cc_200 N_B2_c_246_n N_VPWR_c_346_n 0.00490557f $X=2.665 $Y=1.765 $X2=0 $Y2=0
cc_201 N_B2_c_246_n N_VPWR_c_339_n 0.00508379f $X=2.665 $Y=1.765 $X2=0 $Y2=0
cc_202 N_B2_M1002_g N_VGND_c_389_n 0.00290288f $X=2.68 $Y=0.69 $X2=0 $Y2=0
cc_203 N_B2_M1002_g N_VGND_c_390_n 0.00360251f $X=2.68 $Y=0.69 $X2=0 $Y2=0
cc_204 N_B2_M1002_g N_A_251_74#_c_428_n 0.00155078f $X=2.68 $Y=0.69 $X2=0 $Y2=0
cc_205 N_B2_c_248_n N_A_251_74#_c_428_n 0.00217387f $X=2.74 $Y=1.515 $X2=0 $Y2=0
cc_206 N_B2_M1002_g N_A_251_74#_c_431_n 0.0152406f $X=2.68 $Y=0.69 $X2=0 $Y2=0
cc_207 N_B1_c_285_n N_VPWR_c_341_n 0.0065298f $X=3.26 $Y=1.765 $X2=0 $Y2=0
cc_208 N_B1_c_285_n N_VPWR_c_343_n 0.0141252f $X=3.26 $Y=1.765 $X2=0 $Y2=0
cc_209 B1 N_VPWR_c_344_n 0.020013f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_210 N_B1_c_283_n N_VPWR_c_344_n 0.00105029f $X=3.57 $Y=1.345 $X2=0 $Y2=0
cc_211 N_B1_c_285_n N_VPWR_c_346_n 0.00443511f $X=3.26 $Y=1.765 $X2=0 $Y2=0
cc_212 N_B1_c_285_n N_VPWR_c_339_n 0.00460931f $X=3.26 $Y=1.765 $X2=0 $Y2=0
cc_213 N_B1_M1000_g N_VGND_c_389_n 0.00290288f $X=3.275 $Y=0.69 $X2=0 $Y2=0
cc_214 N_B1_M1000_g N_VGND_c_390_n 0.00363413f $X=3.275 $Y=0.69 $X2=0 $Y2=0
cc_215 N_B1_M1000_g N_A_251_74#_c_431_n 0.0130694f $X=3.275 $Y=0.69 $X2=0 $Y2=0
cc_216 B1 N_A_251_74#_c_432_n 0.0210212f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_217 N_B1_c_283_n N_A_251_74#_c_432_n 0.00210773f $X=3.57 $Y=1.345 $X2=0 $Y2=0
cc_218 N_X_c_315_n N_VPWR_c_340_n 0.027028f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_219 N_X_c_315_n N_VPWR_c_345_n 0.0159324f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_220 N_X_c_315_n N_VPWR_c_339_n 0.0131546f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_221 N_X_c_313_n N_VGND_c_383_n 0.0277278f $X=0.395 $Y=0.515 $X2=0 $Y2=0
cc_222 N_X_c_313_n N_VGND_c_385_n 0.021034f $X=0.395 $Y=0.515 $X2=0 $Y2=0
cc_223 N_X_c_313_n N_VGND_c_390_n 0.0173537f $X=0.395 $Y=0.515 $X2=0 $Y2=0
cc_224 X N_A_251_74#_c_429_n 0.00259535f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_225 N_VGND_c_383_n N_A_251_74#_c_427_n 0.0255177f $X=0.895 $Y=0.515 $X2=0
+ $Y2=0
cc_226 N_VGND_c_384_n N_A_251_74#_c_427_n 0.018426f $X=1.895 $Y=0.655 $X2=0
+ $Y2=0
cc_227 N_VGND_c_387_n N_A_251_74#_c_427_n 0.0144922f $X=1.73 $Y=0 $X2=0 $Y2=0
cc_228 N_VGND_c_390_n N_A_251_74#_c_427_n 0.0118826f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_229 N_VGND_c_384_n N_A_251_74#_c_428_n 0.0241019f $X=1.895 $Y=0.655 $X2=0
+ $Y2=0
cc_230 N_VGND_c_383_n N_A_251_74#_c_429_n 0.00163629f $X=0.895 $Y=0.515 $X2=0
+ $Y2=0
cc_231 N_VGND_c_384_n N_A_251_74#_c_430_n 0.00879395f $X=1.895 $Y=0.655 $X2=0
+ $Y2=0
cc_232 N_VGND_c_389_n N_A_251_74#_c_430_n 0.0152637f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_233 N_VGND_c_390_n N_A_251_74#_c_430_n 0.0121407f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_234 N_VGND_c_389_n N_A_251_74#_c_431_n 0.0348412f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_235 N_VGND_c_390_n N_A_251_74#_c_431_n 0.0286968f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_236 N_VGND_c_389_n N_A_251_74#_c_432_n 0.0116085f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_237 N_VGND_c_390_n N_A_251_74#_c_432_n 0.00928389f $X=3.6 $Y=0 $X2=0 $Y2=0
