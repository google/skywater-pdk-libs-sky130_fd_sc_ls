* File: sky130_fd_sc_ls__einvp_8.pxi.spice
* Created: Wed Sep  2 11:07:25 2020
* 
x_PM_SKY130_FD_SC_LS__EINVP_8%A N_A_c_177_n N_A_M1005_g N_A_c_187_n N_A_M1000_g
+ N_A_c_178_n N_A_M1009_g N_A_c_188_n N_A_M1003_g N_A_c_189_n N_A_M1010_g
+ N_A_c_179_n N_A_M1014_g N_A_c_190_n N_A_M1018_g N_A_c_180_n N_A_M1016_g
+ N_A_c_191_n N_A_M1021_g N_A_c_181_n N_A_M1020_g N_A_c_192_n N_A_M1022_g
+ N_A_c_182_n N_A_M1023_g N_A_c_193_n N_A_M1025_g N_A_c_183_n N_A_M1026_g
+ N_A_c_194_n N_A_M1031_g N_A_c_184_n N_A_M1027_g A A A A A N_A_c_185_n
+ N_A_c_186_n PM_SKY130_FD_SC_LS__EINVP_8%A
x_PM_SKY130_FD_SC_LS__EINVP_8%A_802_323# N_A_802_323#_M1033_s
+ N_A_802_323#_M1013_s N_A_802_323#_c_353_n N_A_802_323#_M1001_g
+ N_A_802_323#_c_334_n N_A_802_323#_c_335_n N_A_802_323#_c_356_n
+ N_A_802_323#_M1002_g N_A_802_323#_c_336_n N_A_802_323#_c_358_n
+ N_A_802_323#_M1006_g N_A_802_323#_c_337_n N_A_802_323#_c_360_n
+ N_A_802_323#_M1007_g N_A_802_323#_c_338_n N_A_802_323#_c_362_n
+ N_A_802_323#_M1008_g N_A_802_323#_c_339_n N_A_802_323#_c_364_n
+ N_A_802_323#_M1011_g N_A_802_323#_c_340_n N_A_802_323#_c_366_n
+ N_A_802_323#_M1019_g N_A_802_323#_c_341_n N_A_802_323#_c_368_n
+ N_A_802_323#_M1028_g N_A_802_323#_c_342_n N_A_802_323#_c_343_n
+ N_A_802_323#_c_344_n N_A_802_323#_c_345_n N_A_802_323#_c_346_n
+ N_A_802_323#_c_347_n N_A_802_323#_c_348_n N_A_802_323#_c_349_n
+ N_A_802_323#_c_350_n N_A_802_323#_c_377_n N_A_802_323#_c_351_n
+ N_A_802_323#_c_352_n PM_SKY130_FD_SC_LS__EINVP_8%A_802_323#
x_PM_SKY130_FD_SC_LS__EINVP_8%TE N_TE_c_514_n N_TE_M1004_g N_TE_c_515_n
+ N_TE_c_516_n N_TE_c_517_n N_TE_M1012_g N_TE_c_518_n N_TE_c_519_n N_TE_M1015_g
+ N_TE_c_520_n N_TE_c_521_n N_TE_M1017_g N_TE_c_522_n N_TE_c_523_n N_TE_M1024_g
+ N_TE_c_524_n N_TE_c_525_n N_TE_M1029_g N_TE_c_526_n N_TE_c_527_n N_TE_M1030_g
+ N_TE_c_528_n N_TE_c_529_n N_TE_M1032_g N_TE_c_530_n N_TE_c_531_n N_TE_M1033_g
+ N_TE_c_532_n N_TE_M1013_g N_TE_c_533_n N_TE_c_534_n N_TE_c_535_n N_TE_c_536_n
+ N_TE_c_537_n N_TE_c_538_n N_TE_c_539_n TE PM_SKY130_FD_SC_LS__EINVP_8%TE
x_PM_SKY130_FD_SC_LS__EINVP_8%A_27_368# N_A_27_368#_M1000_d N_A_27_368#_M1003_d
+ N_A_27_368#_M1018_d N_A_27_368#_M1022_d N_A_27_368#_M1031_d
+ N_A_27_368#_M1002_d N_A_27_368#_M1007_d N_A_27_368#_M1011_d
+ N_A_27_368#_M1028_d N_A_27_368#_c_670_n N_A_27_368#_c_671_n
+ N_A_27_368#_c_672_n N_A_27_368#_c_759_p N_A_27_368#_c_673_n
+ N_A_27_368#_c_763_p N_A_27_368#_c_674_n N_A_27_368#_c_766_p
+ N_A_27_368#_c_675_n N_A_27_368#_c_693_n N_A_27_368#_c_694_n
+ N_A_27_368#_c_697_n N_A_27_368#_c_676_n N_A_27_368#_c_677_n
+ N_A_27_368#_c_664_n N_A_27_368#_c_665_n N_A_27_368#_c_678_n
+ N_A_27_368#_c_666_n N_A_27_368#_c_679_n N_A_27_368#_c_667_n
+ N_A_27_368#_c_680_n N_A_27_368#_c_681_n N_A_27_368#_c_682_n
+ N_A_27_368#_c_683_n N_A_27_368#_c_739_n N_A_27_368#_c_668_n
+ N_A_27_368#_c_669_n PM_SKY130_FD_SC_LS__EINVP_8%A_27_368#
x_PM_SKY130_FD_SC_LS__EINVP_8%Z N_Z_M1005_s N_Z_M1014_s N_Z_M1020_s N_Z_M1026_s
+ N_Z_M1000_s N_Z_M1010_s N_Z_M1021_s N_Z_M1025_s N_Z_c_836_n N_Z_c_829_n
+ N_Z_c_830_n N_Z_c_847_n N_Z_c_831_n N_Z_c_855_n N_Z_c_832_n N_Z_c_863_n
+ N_Z_c_866_n N_Z_c_827_n N_Z_c_873_n N_Z_c_833_n N_Z_c_881_n N_Z_c_885_n
+ N_Z_c_834_n N_Z_c_892_n N_Z_c_895_n N_Z_c_898_n Z
+ PM_SKY130_FD_SC_LS__EINVP_8%Z
x_PM_SKY130_FD_SC_LS__EINVP_8%VPWR N_VPWR_M1001_s N_VPWR_M1006_s N_VPWR_M1008_s
+ N_VPWR_M1019_s N_VPWR_M1013_d N_VPWR_c_958_n N_VPWR_c_959_n N_VPWR_c_960_n
+ N_VPWR_c_961_n N_VPWR_c_962_n N_VPWR_c_963_n N_VPWR_c_964_n N_VPWR_c_965_n
+ N_VPWR_c_966_n N_VPWR_c_967_n N_VPWR_c_968_n VPWR N_VPWR_c_969_n
+ N_VPWR_c_970_n N_VPWR_c_971_n N_VPWR_c_972_n N_VPWR_c_957_n
+ PM_SKY130_FD_SC_LS__EINVP_8%VPWR
x_PM_SKY130_FD_SC_LS__EINVP_8%A_27_74# N_A_27_74#_M1005_d N_A_27_74#_M1009_d
+ N_A_27_74#_M1016_d N_A_27_74#_M1023_d N_A_27_74#_M1027_d N_A_27_74#_M1012_d
+ N_A_27_74#_M1017_d N_A_27_74#_M1029_d N_A_27_74#_M1032_d N_A_27_74#_c_1068_n
+ N_A_27_74#_c_1069_n N_A_27_74#_c_1070_n N_A_27_74#_c_1071_n
+ N_A_27_74#_c_1072_n N_A_27_74#_c_1073_n N_A_27_74#_c_1074_n
+ N_A_27_74#_c_1075_n N_A_27_74#_c_1076_n N_A_27_74#_c_1077_n
+ N_A_27_74#_c_1078_n N_A_27_74#_c_1079_n N_A_27_74#_c_1080_n
+ N_A_27_74#_c_1081_n N_A_27_74#_c_1082_n N_A_27_74#_c_1083_n
+ N_A_27_74#_c_1084_n N_A_27_74#_c_1085_n N_A_27_74#_c_1086_n
+ N_A_27_74#_c_1087_n N_A_27_74#_c_1088_n N_A_27_74#_c_1089_n
+ PM_SKY130_FD_SC_LS__EINVP_8%A_27_74#
x_PM_SKY130_FD_SC_LS__EINVP_8%VGND N_VGND_M1004_s N_VGND_M1015_s N_VGND_M1024_s
+ N_VGND_M1030_s N_VGND_M1033_d N_VGND_c_1240_n N_VGND_c_1241_n N_VGND_c_1242_n
+ N_VGND_c_1243_n N_VGND_c_1244_n N_VGND_c_1245_n N_VGND_c_1246_n
+ N_VGND_c_1247_n VGND N_VGND_c_1248_n N_VGND_c_1249_n N_VGND_c_1250_n
+ N_VGND_c_1251_n N_VGND_c_1252_n N_VGND_c_1253_n N_VGND_c_1254_n
+ N_VGND_c_1255_n PM_SKY130_FD_SC_LS__EINVP_8%VGND
cc_1 VNB N_A_c_177_n 0.0207336f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_A_c_178_n 0.0165475f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.22
cc_3 VNB N_A_c_179_n 0.0171712f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.22
cc_4 VNB N_A_c_180_n 0.0171914f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.22
cc_5 VNB N_A_c_181_n 0.0171712f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=1.22
cc_6 VNB N_A_c_182_n 0.0171914f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=1.22
cc_7 VNB N_A_c_183_n 0.0172959f $X=-0.19 $Y=-0.245 $X2=3.425 $Y2=1.22
cc_8 VNB N_A_c_184_n 0.0165598f $X=-0.19 $Y=-0.245 $X2=3.925 $Y2=1.22
cc_9 VNB N_A_c_185_n 0.0355723f $X=-0.19 $Y=-0.245 $X2=3.295 $Y2=1.385
cc_10 VNB N_A_c_186_n 0.244074f $X=-0.19 $Y=-0.245 $X2=3.65 $Y2=1.492
cc_11 VNB N_A_802_323#_c_334_n 0.00771672f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.765
cc_12 VNB N_A_802_323#_c_335_n 0.00607832f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.4
cc_13 VNB N_A_802_323#_c_336_n 0.00537118f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=2.4
cc_14 VNB N_A_802_323#_c_337_n 0.00494563f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=2.4
cc_15 VNB N_A_802_323#_c_338_n 0.00493383f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.765
cc_16 VNB N_A_802_323#_c_339_n 0.00494563f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=0.74
cc_17 VNB N_A_802_323#_c_340_n 0.00493383f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=0.74
cc_18 VNB N_A_802_323#_c_341_n 0.00494563f $X=-0.19 $Y=-0.245 $X2=3.425 $Y2=1.22
cc_19 VNB N_A_802_323#_c_342_n 0.0150523f $X=-0.19 $Y=-0.245 $X2=3.65 $Y2=2.4
cc_20 VNB N_A_802_323#_c_343_n 0.00348356f $X=-0.19 $Y=-0.245 $X2=3.925 $Y2=0.74
cc_21 VNB N_A_802_323#_c_344_n 0.00247438f $X=-0.19 $Y=-0.245 $X2=3.925 $Y2=0.74
cc_22 VNB N_A_802_323#_c_345_n 0.00247438f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_23 VNB N_A_802_323#_c_346_n 0.00248618f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_24 VNB N_A_802_323#_c_347_n 0.00247438f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_25 VNB N_A_802_323#_c_348_n 0.00248618f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.21
cc_26 VNB N_A_802_323#_c_349_n 0.00247438f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=1.21
cc_27 VNB N_A_802_323#_c_350_n 0.0113187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_802_323#_c_351_n 0.00336983f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=1.385
cc_29 VNB N_A_802_323#_c_352_n 0.0117383f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=1.385
cc_30 VNB N_TE_c_514_n 0.0173552f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_31 VNB N_TE_c_515_n 0.0145237f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.765
cc_32 VNB N_TE_c_516_n 0.00615296f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.4
cc_33 VNB N_TE_c_517_n 0.0171627f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.4
cc_34 VNB N_TE_c_518_n 0.0105631f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_35 VNB N_TE_c_519_n 0.0163632f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.4
cc_36 VNB N_TE_c_520_n 0.0105749f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=2.4
cc_37 VNB N_TE_c_521_n 0.0163604f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.22
cc_38 VNB N_TE_c_522_n 0.0105513f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.765
cc_39 VNB N_TE_c_523_n 0.0163604f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=2.4
cc_40 VNB N_TE_c_524_n 0.0105749f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_41 VNB N_TE_c_525_n 0.0163632f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=2.4
cc_42 VNB N_TE_c_526_n 0.0105631f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=0.74
cc_43 VNB N_TE_c_527_n 0.0171627f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=1.765
cc_44 VNB N_TE_c_528_n 0.0145237f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=1.22
cc_45 VNB N_TE_c_529_n 0.0208358f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=0.74
cc_46 VNB N_TE_c_530_n 0.0528403f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=2.4
cc_47 VNB N_TE_c_531_n 0.0245639f $X=-0.19 $Y=-0.245 $X2=3.425 $Y2=0.74
cc_48 VNB N_TE_c_532_n 0.0443573f $X=-0.19 $Y=-0.245 $X2=3.65 $Y2=2.4
cc_49 VNB N_TE_c_533_n 0.00414591f $X=-0.19 $Y=-0.245 $X2=3.925 $Y2=0.74
cc_50 VNB N_TE_c_534_n 0.00415771f $X=-0.19 $Y=-0.245 $X2=3.925 $Y2=0.74
cc_51 VNB N_TE_c_535_n 0.00415771f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_52 VNB N_TE_c_536_n 0.00415771f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_53 VNB N_TE_c_537_n 0.00415771f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_54 VNB N_TE_c_538_n 0.00414591f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.21
cc_55 VNB N_TE_c_539_n 0.00415771f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=1.21
cc_56 VNB TE 0.0297385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_27_368#_c_664_n 0.00342583f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=1.492
cc_58 VNB N_A_27_368#_c_665_n 0.00250548f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=1.385
cc_59 VNB N_A_27_368#_c_666_n 0.00390912f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.492
cc_60 VNB N_A_27_368#_c_667_n 0.00641513f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=1.385
cc_61 VNB N_A_27_368#_c_668_n 0.00154195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_27_368#_c_669_n 0.00154195f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=1.365
cc_63 VNB N_Z_c_827_n 0.00686569f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.385
cc_64 VNB Z 0.0056279f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=1.385
cc_65 VNB N_VPWR_c_957_n 0.382608f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=1.492
cc_66 VNB N_A_27_74#_c_1068_n 0.0229491f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=0.74
cc_67 VNB N_A_27_74#_c_1069_n 0.00254822f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=2.4
cc_68 VNB N_A_27_74#_c_1070_n 0.00971634f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=2.4
cc_69 VNB N_A_27_74#_c_1071_n 0.00304663f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=1.22
cc_70 VNB N_A_27_74#_c_1072_n 0.00304663f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=0.74
cc_71 VNB N_A_27_74#_c_1073_n 0.00499169f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=2.4
cc_72 VNB N_A_27_74#_c_1074_n 0.00162809f $X=-0.19 $Y=-0.245 $X2=3.65 $Y2=1.765
cc_73 VNB N_A_27_74#_c_1075_n 0.0122249f $X=-0.19 $Y=-0.245 $X2=3.65 $Y2=2.4
cc_74 VNB N_A_27_74#_c_1076_n 0.00255778f $X=-0.19 $Y=-0.245 $X2=3.65 $Y2=2.4
cc_75 VNB N_A_27_74#_c_1077_n 0.00299989f $X=-0.19 $Y=-0.245 $X2=3.925 $Y2=0.74
cc_76 VNB N_A_27_74#_c_1078_n 0.010543f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_77 VNB N_A_27_74#_c_1079_n 0.00356911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_27_74#_c_1080_n 0.010543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_27_74#_c_1081_n 0.00299989f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.492
cc_80 VNB N_A_27_74#_c_1082_n 0.0133095f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.385
cc_81 VNB N_A_27_74#_c_1083_n 0.0102993f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=1.492
cc_82 VNB N_A_27_74#_c_1084_n 0.00240543f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=1.385
cc_83 VNB N_A_27_74#_c_1085_n 0.00240543f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.385
cc_84 VNB N_A_27_74#_c_1086_n 0.00240543f $X=-0.19 $Y=-0.245 $X2=2.275 $Y2=1.385
cc_85 VNB N_A_27_74#_c_1087_n 0.00158451f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=1.385
cc_86 VNB N_A_27_74#_c_1088_n 0.00107773f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=1.492
cc_87 VNB N_A_27_74#_c_1089_n 0.0015849f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=1.492
cc_88 VNB N_VGND_c_1240_n 0.00558127f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_89 VNB N_VGND_c_1241_n 0.002601f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.22
cc_90 VNB N_VGND_c_1242_n 0.002601f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=2.4
cc_91 VNB N_VGND_c_1243_n 0.00558127f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=0.74
cc_92 VNB N_VGND_c_1244_n 0.0131032f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=2.4
cc_93 VNB N_VGND_c_1245_n 0.0361666f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=1.22
cc_94 VNB N_VGND_c_1246_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=1.765
cc_95 VNB N_VGND_c_1247_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=2.4
cc_96 VNB N_VGND_c_1248_n 0.102301f $X=-0.19 $Y=-0.245 $X2=3.425 $Y2=0.74
cc_97 VNB N_VGND_c_1249_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_98 VNB N_VGND_c_1250_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1251_n 0.0331641f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.385
cc_100 VNB N_VGND_c_1252_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=1.385
cc_101 VNB N_VGND_c_1253_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.492
cc_102 VNB N_VGND_c_1254_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.492
cc_103 VNB N_VGND_c_1255_n 0.488212f $X=-0.19 $Y=-0.245 $X2=2.275 $Y2=1.385
cc_104 VPB N_A_c_187_n 0.0181192f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.765
cc_105 VPB N_A_c_188_n 0.0141098f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.765
cc_106 VPB N_A_c_189_n 0.0141098f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.765
cc_107 VPB N_A_c_190_n 0.0141098f $X=-0.19 $Y=1.66 $X2=1.85 $Y2=1.765
cc_108 VPB N_A_c_191_n 0.0141098f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.765
cc_109 VPB N_A_c_192_n 0.0141098f $X=-0.19 $Y=1.66 $X2=2.75 $Y2=1.765
cc_110 VPB N_A_c_193_n 0.0141098f $X=-0.19 $Y=1.66 $X2=3.2 $Y2=1.765
cc_111 VPB N_A_c_194_n 0.0141395f $X=-0.19 $Y=1.66 $X2=3.65 $Y2=1.765
cc_112 VPB N_A_c_186_n 0.0521263f $X=-0.19 $Y=1.66 $X2=3.65 $Y2=1.492
cc_113 VPB N_A_802_323#_c_353_n 0.0146233f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.22
cc_114 VPB N_A_802_323#_c_334_n 0.0062311f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.765
cc_115 VPB N_A_802_323#_c_335_n 0.00362133f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.4
cc_116 VPB N_A_802_323#_c_356_n 0.015069f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.4
cc_117 VPB N_A_802_323#_c_336_n 0.00675749f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=2.4
cc_118 VPB N_A_802_323#_c_358_n 0.0152877f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_119 VPB N_A_802_323#_c_337_n 0.00593398f $X=-0.19 $Y=1.66 $X2=1.85 $Y2=2.4
cc_120 VPB N_A_802_323#_c_360_n 0.0152877f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=1.22
cc_121 VPB N_A_802_323#_c_338_n 0.00675749f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.765
cc_122 VPB N_A_802_323#_c_362_n 0.0150768f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=2.4
cc_123 VPB N_A_802_323#_c_339_n 0.00593398f $X=-0.19 $Y=1.66 $X2=2.425 $Y2=0.74
cc_124 VPB N_A_802_323#_c_364_n 0.01529f $X=-0.19 $Y=1.66 $X2=2.75 $Y2=2.4
cc_125 VPB N_A_802_323#_c_340_n 0.00675749f $X=-0.19 $Y=1.66 $X2=2.925 $Y2=0.74
cc_126 VPB N_A_802_323#_c_366_n 0.0150768f $X=-0.19 $Y=1.66 $X2=3.2 $Y2=1.765
cc_127 VPB N_A_802_323#_c_341_n 0.00593398f $X=-0.19 $Y=1.66 $X2=3.425 $Y2=1.22
cc_128 VPB N_A_802_323#_c_368_n 0.0189382f $X=-0.19 $Y=1.66 $X2=3.425 $Y2=0.74
cc_129 VPB N_A_802_323#_c_342_n 0.0206571f $X=-0.19 $Y=1.66 $X2=3.65 $Y2=2.4
cc_130 VPB N_A_802_323#_c_343_n 0.00167153f $X=-0.19 $Y=1.66 $X2=3.925 $Y2=0.74
cc_131 VPB N_A_802_323#_c_344_n 0.00167153f $X=-0.19 $Y=1.66 $X2=3.925 $Y2=0.74
cc_132 VPB N_A_802_323#_c_345_n 0.00167153f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.21
cc_133 VPB N_A_802_323#_c_346_n 0.00167153f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.21
cc_134 VPB N_A_802_323#_c_347_n 0.00167153f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.21
cc_135 VPB N_A_802_323#_c_348_n 0.00167153f $X=-0.19 $Y=1.66 $X2=2.555 $Y2=1.21
cc_136 VPB N_A_802_323#_c_349_n 0.00167153f $X=-0.19 $Y=1.66 $X2=3.035 $Y2=1.21
cc_137 VPB N_A_802_323#_c_377_n 0.0967593f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.492
cc_138 VPB N_A_802_323#_c_351_n 0.0222215f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=1.385
cc_139 VPB N_TE_c_532_n 0.0321294f $X=-0.19 $Y=1.66 $X2=3.65 $Y2=2.4
cc_140 VPB N_A_27_368#_c_670_n 0.051291f $X=-0.19 $Y=1.66 $X2=2.425 $Y2=0.74
cc_141 VPB N_A_27_368#_c_671_n 0.0027982f $X=-0.19 $Y=1.66 $X2=2.925 $Y2=1.22
cc_142 VPB N_A_27_368#_c_672_n 0.00947786f $X=-0.19 $Y=1.66 $X2=2.925 $Y2=0.74
cc_143 VPB N_A_27_368#_c_673_n 0.0027982f $X=-0.19 $Y=1.66 $X2=3.425 $Y2=1.22
cc_144 VPB N_A_27_368#_c_674_n 0.002727f $X=-0.19 $Y=1.66 $X2=3.925 $Y2=1.22
cc_145 VPB N_A_27_368#_c_675_n 0.00512904f $X=-0.19 $Y=1.66 $X2=2.555 $Y2=1.21
cc_146 VPB N_A_27_368#_c_676_n 6.40903e-19 $X=-0.19 $Y=1.66 $X2=0.915 $Y2=1.492
cc_147 VPB N_A_27_368#_c_677_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.492
cc_148 VPB N_A_27_368#_c_678_n 0.00280674f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.492
cc_149 VPB N_A_27_368#_c_679_n 0.00280674f $X=-0.19 $Y=1.66 $X2=2.275 $Y2=1.385
cc_150 VPB N_A_27_368#_c_680_n 0.00283383f $X=-0.19 $Y=1.66 $X2=3.2 $Y2=1.492
cc_151 VPB N_A_27_368#_c_681_n 0.00149233f $X=-0.19 $Y=1.66 $X2=3.425 $Y2=1.492
cc_152 VPB N_A_27_368#_c_682_n 0.00160153f $X=-0.19 $Y=1.66 $X2=3.65 $Y2=1.492
cc_153 VPB N_A_27_368#_c_683_n 0.00145593f $X=-0.19 $Y=1.66 $X2=3.925 $Y2=1.22
cc_154 VPB N_Z_c_829_n 0.00219429f $X=-0.19 $Y=1.66 $X2=2.75 $Y2=2.4
cc_155 VPB N_Z_c_830_n 0.00224287f $X=-0.19 $Y=1.66 $X2=2.925 $Y2=1.22
cc_156 VPB N_Z_c_831_n 0.00219429f $X=-0.19 $Y=1.66 $X2=3.425 $Y2=0.74
cc_157 VPB N_Z_c_832_n 0.00219429f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.21
cc_158 VPB N_Z_c_833_n 0.00224287f $X=-0.19 $Y=1.66 $X2=1.255 $Y2=1.385
cc_159 VPB N_Z_c_834_n 0.00224287f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.385
cc_160 VPB Z 0.00582828f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=1.385
cc_161 VPB N_VPWR_c_958_n 0.00339119f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_162 VPB N_VPWR_c_959_n 0.00670059f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=1.22
cc_163 VPB N_VPWR_c_960_n 0.0185253f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=2.4
cc_164 VPB N_VPWR_c_961_n 0.00444486f $X=-0.19 $Y=1.66 $X2=2.425 $Y2=0.74
cc_165 VPB N_VPWR_c_962_n 0.00514362f $X=-0.19 $Y=1.66 $X2=2.925 $Y2=0.74
cc_166 VPB N_VPWR_c_963_n 0.0103331f $X=-0.19 $Y=1.66 $X2=3.425 $Y2=1.22
cc_167 VPB N_VPWR_c_964_n 0.0587564f $X=-0.19 $Y=1.66 $X2=3.425 $Y2=0.74
cc_168 VPB N_VPWR_c_965_n 0.0971135f $X=-0.19 $Y=1.66 $X2=3.925 $Y2=0.74
cc_169 VPB N_VPWR_c_966_n 0.00601644f $X=-0.19 $Y=1.66 $X2=3.925 $Y2=0.74
cc_170 VPB N_VPWR_c_967_n 0.0185253f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.21
cc_171 VPB N_VPWR_c_968_n 0.00324402f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.21
cc_172 VPB N_VPWR_c_969_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=1.385
cc_173 VPB N_VPWR_c_970_n 0.0445971f $X=-0.19 $Y=1.66 $X2=1.255 $Y2=1.385
cc_174 VPB N_VPWR_c_971_n 0.00460249f $X=-0.19 $Y=1.66 $X2=2.275 $Y2=1.385
cc_175 VPB N_VPWR_c_972_n 0.00460249f $X=-0.19 $Y=1.66 $X2=2.425 $Y2=1.492
cc_176 VPB N_VPWR_c_957_n 0.110506f $X=-0.19 $Y=1.66 $X2=2.75 $Y2=1.492
cc_177 N_A_c_194_n N_A_802_323#_c_353_n 0.0222615f $X=3.65 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A_c_186_n N_A_802_323#_c_335_n 0.00713346f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_179 N_A_c_184_n N_TE_c_514_n 0.00900363f $X=3.925 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_180 N_A_c_186_n N_TE_c_516_n 0.00900363f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_181 N_A_c_187_n N_A_27_368#_c_670_n 0.00141178f $X=0.5 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A_c_187_n N_A_27_368#_c_671_n 0.0136604f $X=0.5 $Y=1.765 $X2=0 $Y2=0
cc_183 N_A_c_188_n N_A_27_368#_c_671_n 0.0128349f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A_c_189_n N_A_27_368#_c_673_n 0.0128349f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_185 N_A_c_190_n N_A_27_368#_c_673_n 0.0128349f $X=1.85 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A_c_191_n N_A_27_368#_c_674_n 0.0128349f $X=2.3 $Y=1.765 $X2=0 $Y2=0
cc_187 N_A_c_192_n N_A_27_368#_c_674_n 0.0128349f $X=2.75 $Y=1.765 $X2=0 $Y2=0
cc_188 N_A_c_193_n N_A_27_368#_c_675_n 0.0127839f $X=3.2 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A_c_194_n N_A_27_368#_c_675_n 0.012504f $X=3.65 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A_c_186_n N_A_27_368#_c_693_n 3.56962e-19 $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_191 N_A_c_194_n N_A_27_368#_c_694_n 0.0057515f $X=3.65 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A_c_187_n N_Z_c_836_n 0.00892248f $X=0.5 $Y=1.765 $X2=0 $Y2=0
cc_193 N_A_c_188_n N_Z_c_836_n 0.00968252f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_194 N_A_c_189_n N_Z_c_836_n 6.21854e-19 $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_195 N_A_c_188_n N_Z_c_829_n 0.00903574f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A_c_189_n N_Z_c_829_n 0.00903574f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_197 N_A_c_185_n N_Z_c_829_n 0.042029f $X=3.295 $Y=1.385 $X2=0 $Y2=0
cc_198 N_A_c_186_n N_Z_c_829_n 0.00885373f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_199 N_A_c_187_n N_Z_c_830_n 0.00415728f $X=0.5 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A_c_188_n N_Z_c_830_n 0.00109449f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A_c_185_n N_Z_c_830_n 0.0277828f $X=3.295 $Y=1.385 $X2=0 $Y2=0
cc_202 N_A_c_186_n N_Z_c_830_n 0.00708762f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_203 N_A_c_188_n N_Z_c_847_n 6.26672e-19 $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_204 N_A_c_189_n N_Z_c_847_n 0.00976089f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_205 N_A_c_190_n N_Z_c_847_n 0.00968252f $X=1.85 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A_c_191_n N_Z_c_847_n 6.21854e-19 $X=2.3 $Y=1.765 $X2=0 $Y2=0
cc_207 N_A_c_190_n N_Z_c_831_n 0.00903574f $X=1.85 $Y=1.765 $X2=0 $Y2=0
cc_208 N_A_c_191_n N_Z_c_831_n 0.00903574f $X=2.3 $Y=1.765 $X2=0 $Y2=0
cc_209 N_A_c_185_n N_Z_c_831_n 0.042029f $X=3.295 $Y=1.385 $X2=0 $Y2=0
cc_210 N_A_c_186_n N_Z_c_831_n 0.00909013f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_211 N_A_c_190_n N_Z_c_855_n 6.12174e-19 $X=1.85 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A_c_191_n N_Z_c_855_n 0.00952605f $X=2.3 $Y=1.765 $X2=0 $Y2=0
cc_213 N_A_c_192_n N_Z_c_855_n 0.00976089f $X=2.75 $Y=1.765 $X2=0 $Y2=0
cc_214 N_A_c_193_n N_Z_c_855_n 6.26672e-19 $X=3.2 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A_c_192_n N_Z_c_832_n 0.00903574f $X=2.75 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A_c_193_n N_Z_c_832_n 0.00903574f $X=3.2 $Y=1.765 $X2=0 $Y2=0
cc_217 N_A_c_185_n N_Z_c_832_n 0.042029f $X=3.295 $Y=1.385 $X2=0 $Y2=0
cc_218 N_A_c_186_n N_Z_c_832_n 0.00920833f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_219 N_A_c_182_n N_Z_c_863_n 0.00874124f $X=2.925 $Y=1.22 $X2=0 $Y2=0
cc_220 N_A_c_183_n N_Z_c_863_n 0.0121141f $X=3.425 $Y=1.22 $X2=0 $Y2=0
cc_221 N_A_c_186_n N_Z_c_863_n 0.0010599f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_222 N_A_c_192_n N_Z_c_866_n 6.26672e-19 $X=2.75 $Y=1.765 $X2=0 $Y2=0
cc_223 N_A_c_193_n N_Z_c_866_n 0.00976089f $X=3.2 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A_c_194_n N_Z_c_866_n 0.0100248f $X=3.65 $Y=1.765 $X2=0 $Y2=0
cc_225 N_A_c_183_n N_Z_c_827_n 0.00374449f $X=3.425 $Y=1.22 $X2=0 $Y2=0
cc_226 N_A_c_184_n N_Z_c_827_n 0.00399031f $X=3.925 $Y=1.22 $X2=0 $Y2=0
cc_227 N_A_c_185_n N_Z_c_827_n 0.021022f $X=3.295 $Y=1.385 $X2=0 $Y2=0
cc_228 N_A_c_186_n N_Z_c_827_n 0.0169783f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_229 N_A_c_178_n N_Z_c_873_n 0.00582792f $X=0.925 $Y=1.22 $X2=0 $Y2=0
cc_230 N_A_c_179_n N_Z_c_873_n 4.41837e-19 $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_231 N_A_c_185_n N_Z_c_873_n 0.0182538f $X=3.295 $Y=1.385 $X2=0 $Y2=0
cc_232 N_A_c_186_n N_Z_c_873_n 6.73904e-19 $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_233 N_A_c_189_n N_Z_c_833_n 0.00109449f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A_c_190_n N_Z_c_833_n 0.00109449f $X=1.85 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A_c_185_n N_Z_c_833_n 0.0277828f $X=3.295 $Y=1.385 $X2=0 $Y2=0
cc_236 N_A_c_186_n N_Z_c_833_n 0.00505568f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_237 N_A_c_178_n N_Z_c_881_n 0.00935149f $X=0.925 $Y=1.22 $X2=0 $Y2=0
cc_238 N_A_c_179_n N_Z_c_881_n 0.0123177f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_239 N_A_c_185_n N_Z_c_881_n 0.180071f $X=3.295 $Y=1.385 $X2=0 $Y2=0
cc_240 N_A_c_186_n N_Z_c_881_n 0.00106692f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_241 N_A_c_180_n N_Z_c_885_n 0.00553813f $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_242 N_A_c_181_n N_Z_c_885_n 3.58423e-19 $X=2.425 $Y=1.22 $X2=0 $Y2=0
cc_243 N_A_c_186_n N_Z_c_885_n 0.00113983f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_244 N_A_c_191_n N_Z_c_834_n 0.00109449f $X=2.3 $Y=1.765 $X2=0 $Y2=0
cc_245 N_A_c_192_n N_Z_c_834_n 0.00109449f $X=2.75 $Y=1.765 $X2=0 $Y2=0
cc_246 N_A_c_185_n N_Z_c_834_n 0.0277828f $X=3.295 $Y=1.385 $X2=0 $Y2=0
cc_247 N_A_c_186_n N_Z_c_834_n 0.00536838f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_248 N_A_c_180_n N_Z_c_892_n 0.00775967f $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_249 N_A_c_181_n N_Z_c_892_n 0.0122113f $X=2.425 $Y=1.22 $X2=0 $Y2=0
cc_250 N_A_c_186_n N_Z_c_892_n 0.00106239f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_251 N_A_c_182_n N_Z_c_895_n 0.00554054f $X=2.925 $Y=1.22 $X2=0 $Y2=0
cc_252 N_A_c_183_n N_Z_c_895_n 3.58587e-19 $X=3.425 $Y=1.22 $X2=0 $Y2=0
cc_253 N_A_c_186_n N_Z_c_895_n 0.00113363f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_254 N_A_c_184_n N_Z_c_898_n 0.00527055f $X=3.925 $Y=1.22 $X2=0 $Y2=0
cc_255 N_A_c_186_n N_Z_c_898_n 0.00501495f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_256 N_A_c_193_n Z 0.00109449f $X=3.2 $Y=1.765 $X2=0 $Y2=0
cc_257 N_A_c_194_n Z 0.0103343f $X=3.65 $Y=1.765 $X2=0 $Y2=0
cc_258 N_A_c_185_n Z 0.0168664f $X=3.295 $Y=1.385 $X2=0 $Y2=0
cc_259 N_A_c_186_n Z 0.0253351f $X=3.65 $Y=1.492 $X2=0 $Y2=0
cc_260 N_A_c_187_n N_VPWR_c_965_n 0.00278271f $X=0.5 $Y=1.765 $X2=0 $Y2=0
cc_261 N_A_c_188_n N_VPWR_c_965_n 0.00278271f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_262 N_A_c_189_n N_VPWR_c_965_n 0.00278271f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_263 N_A_c_190_n N_VPWR_c_965_n 0.00278271f $X=1.85 $Y=1.765 $X2=0 $Y2=0
cc_264 N_A_c_191_n N_VPWR_c_965_n 0.00278271f $X=2.3 $Y=1.765 $X2=0 $Y2=0
cc_265 N_A_c_192_n N_VPWR_c_965_n 0.00278271f $X=2.75 $Y=1.765 $X2=0 $Y2=0
cc_266 N_A_c_193_n N_VPWR_c_965_n 0.00278271f $X=3.2 $Y=1.765 $X2=0 $Y2=0
cc_267 N_A_c_194_n N_VPWR_c_965_n 0.00278271f $X=3.65 $Y=1.765 $X2=0 $Y2=0
cc_268 N_A_c_187_n N_VPWR_c_957_n 0.003573f $X=0.5 $Y=1.765 $X2=0 $Y2=0
cc_269 N_A_c_188_n N_VPWR_c_957_n 0.00353823f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_270 N_A_c_189_n N_VPWR_c_957_n 0.00353823f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_271 N_A_c_190_n N_VPWR_c_957_n 0.00353823f $X=1.85 $Y=1.765 $X2=0 $Y2=0
cc_272 N_A_c_191_n N_VPWR_c_957_n 0.00353823f $X=2.3 $Y=1.765 $X2=0 $Y2=0
cc_273 N_A_c_192_n N_VPWR_c_957_n 0.00353823f $X=2.75 $Y=1.765 $X2=0 $Y2=0
cc_274 N_A_c_193_n N_VPWR_c_957_n 0.00353823f $X=3.2 $Y=1.765 $X2=0 $Y2=0
cc_275 N_A_c_194_n N_VPWR_c_957_n 0.00353907f $X=3.65 $Y=1.765 $X2=0 $Y2=0
cc_276 N_A_c_177_n N_A_27_74#_c_1068_n 0.00791306f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_277 N_A_c_178_n N_A_27_74#_c_1068_n 6.43486e-19 $X=0.925 $Y=1.22 $X2=0 $Y2=0
cc_278 N_A_c_185_n N_A_27_74#_c_1068_n 0.00231504f $X=3.295 $Y=1.385 $X2=0 $Y2=0
cc_279 N_A_c_177_n N_A_27_74#_c_1069_n 0.0100245f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_280 N_A_c_178_n N_A_27_74#_c_1069_n 0.00926373f $X=0.925 $Y=1.22 $X2=0 $Y2=0
cc_281 N_A_c_177_n N_A_27_74#_c_1070_n 0.00282152f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_282 N_A_c_179_n N_A_27_74#_c_1071_n 0.00823735f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_283 N_A_c_180_n N_A_27_74#_c_1071_n 0.0107668f $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_284 N_A_c_181_n N_A_27_74#_c_1072_n 0.00834679f $X=2.425 $Y=1.22 $X2=0 $Y2=0
cc_285 N_A_c_182_n N_A_27_74#_c_1072_n 0.00967244f $X=2.925 $Y=1.22 $X2=0 $Y2=0
cc_286 N_A_c_183_n N_A_27_74#_c_1073_n 0.00829802f $X=3.425 $Y=1.22 $X2=0 $Y2=0
cc_287 N_A_c_184_n N_A_27_74#_c_1073_n 0.0123973f $X=3.925 $Y=1.22 $X2=0 $Y2=0
cc_288 N_A_c_184_n N_A_27_74#_c_1074_n 9.60276e-19 $X=3.925 $Y=1.22 $X2=0 $Y2=0
cc_289 N_A_c_184_n N_A_27_74#_c_1076_n 0.00159361f $X=3.925 $Y=1.22 $X2=0 $Y2=0
cc_290 N_A_c_178_n N_A_27_74#_c_1084_n 4.46617e-19 $X=0.925 $Y=1.22 $X2=0 $Y2=0
cc_291 N_A_c_179_n N_A_27_74#_c_1084_n 0.00707613f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_292 N_A_c_180_n N_A_27_74#_c_1084_n 6.08486e-19 $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_293 N_A_c_180_n N_A_27_74#_c_1085_n 4.46617e-19 $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_294 N_A_c_181_n N_A_27_74#_c_1085_n 0.00707613f $X=2.425 $Y=1.22 $X2=0 $Y2=0
cc_295 N_A_c_182_n N_A_27_74#_c_1085_n 6.08486e-19 $X=2.925 $Y=1.22 $X2=0 $Y2=0
cc_296 N_A_c_182_n N_A_27_74#_c_1086_n 4.46617e-19 $X=2.925 $Y=1.22 $X2=0 $Y2=0
cc_297 N_A_c_183_n N_A_27_74#_c_1086_n 0.00675729f $X=3.425 $Y=1.22 $X2=0 $Y2=0
cc_298 N_A_c_184_n N_A_27_74#_c_1086_n 8.16033e-19 $X=3.925 $Y=1.22 $X2=0 $Y2=0
cc_299 N_A_c_177_n N_VGND_c_1248_n 0.00278247f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_300 N_A_c_178_n N_VGND_c_1248_n 0.00278271f $X=0.925 $Y=1.22 $X2=0 $Y2=0
cc_301 N_A_c_179_n N_VGND_c_1248_n 0.00279469f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_302 N_A_c_180_n N_VGND_c_1248_n 0.00278271f $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_303 N_A_c_181_n N_VGND_c_1248_n 0.00279469f $X=2.425 $Y=1.22 $X2=0 $Y2=0
cc_304 N_A_c_182_n N_VGND_c_1248_n 0.00278271f $X=2.925 $Y=1.22 $X2=0 $Y2=0
cc_305 N_A_c_183_n N_VGND_c_1248_n 0.00279469f $X=3.425 $Y=1.22 $X2=0 $Y2=0
cc_306 N_A_c_184_n N_VGND_c_1248_n 0.00278271f $X=3.925 $Y=1.22 $X2=0 $Y2=0
cc_307 N_A_c_177_n N_VGND_c_1255_n 0.00357084f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_308 N_A_c_178_n N_VGND_c_1255_n 0.00353178f $X=0.925 $Y=1.22 $X2=0 $Y2=0
cc_309 N_A_c_179_n N_VGND_c_1255_n 0.00353834f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_310 N_A_c_180_n N_VGND_c_1255_n 0.00354745f $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_311 N_A_c_181_n N_VGND_c_1255_n 0.00353834f $X=2.425 $Y=1.22 $X2=0 $Y2=0
cc_312 N_A_c_182_n N_VGND_c_1255_n 0.00354745f $X=2.925 $Y=1.22 $X2=0 $Y2=0
cc_313 N_A_c_183_n N_VGND_c_1255_n 0.00353834f $X=3.425 $Y=1.22 $X2=0 $Y2=0
cc_314 N_A_c_184_n N_VGND_c_1255_n 0.00354184f $X=3.925 $Y=1.22 $X2=0 $Y2=0
cc_315 N_A_802_323#_c_343_n N_TE_c_515_n 0.0135815f $X=4.55 $Y=1.69 $X2=0 $Y2=0
cc_316 N_A_802_323#_c_334_n N_TE_c_516_n 0.0135815f $X=4.475 $Y=1.69 $X2=0 $Y2=0
cc_317 N_A_802_323#_c_344_n N_TE_c_518_n 0.0135815f $X=5 $Y=1.69 $X2=0 $Y2=0
cc_318 N_A_802_323#_c_345_n N_TE_c_520_n 0.0135815f $X=5.45 $Y=1.69 $X2=0 $Y2=0
cc_319 N_A_802_323#_c_346_n N_TE_c_522_n 0.0135815f $X=5.9 $Y=1.69 $X2=0 $Y2=0
cc_320 N_A_802_323#_c_347_n N_TE_c_524_n 0.0135815f $X=6.35 $Y=1.69 $X2=0 $Y2=0
cc_321 N_A_802_323#_c_348_n N_TE_c_526_n 0.0135815f $X=6.8 $Y=1.69 $X2=0 $Y2=0
cc_322 N_A_802_323#_c_349_n N_TE_c_528_n 0.0135815f $X=7.25 $Y=1.69 $X2=0 $Y2=0
cc_323 N_A_802_323#_c_352_n N_TE_c_529_n 0.00128937f $X=8.34 $Y=0.515 $X2=0
+ $Y2=0
cc_324 N_A_802_323#_c_350_n N_TE_c_530_n 0.0141302f $X=8.14 $Y=1.615 $X2=0 $Y2=0
cc_325 N_A_802_323#_c_351_n N_TE_c_530_n 0.00787748f $X=7.94 $Y=2.8 $X2=0 $Y2=0
cc_326 N_A_802_323#_c_352_n N_TE_c_530_n 0.00642168f $X=8.34 $Y=0.515 $X2=0
+ $Y2=0
cc_327 N_A_802_323#_c_350_n N_TE_c_531_n 0.00414962f $X=8.14 $Y=1.615 $X2=0
+ $Y2=0
cc_328 N_A_802_323#_c_352_n N_TE_c_531_n 0.00801467f $X=8.34 $Y=0.515 $X2=0
+ $Y2=0
cc_329 N_A_802_323#_c_342_n N_TE_c_532_n 0.00348971f $X=7.775 $Y=1.69 $X2=0
+ $Y2=0
cc_330 N_A_802_323#_c_350_n N_TE_c_532_n 0.00315476f $X=8.14 $Y=1.615 $X2=0
+ $Y2=0
cc_331 N_A_802_323#_c_377_n N_TE_c_532_n 0.0155693f $X=7.94 $Y=1.78 $X2=0 $Y2=0
cc_332 N_A_802_323#_c_351_n N_TE_c_532_n 0.0202334f $X=7.94 $Y=2.8 $X2=0 $Y2=0
cc_333 N_A_802_323#_c_336_n N_TE_c_533_n 0.0135815f $X=4.925 $Y=1.69 $X2=0 $Y2=0
cc_334 N_A_802_323#_c_337_n N_TE_c_534_n 0.0135815f $X=5.375 $Y=1.69 $X2=0 $Y2=0
cc_335 N_A_802_323#_c_338_n N_TE_c_535_n 0.0135815f $X=5.825 $Y=1.69 $X2=0 $Y2=0
cc_336 N_A_802_323#_c_339_n N_TE_c_536_n 0.0135815f $X=6.275 $Y=1.69 $X2=0 $Y2=0
cc_337 N_A_802_323#_c_340_n N_TE_c_537_n 0.0135815f $X=6.725 $Y=1.69 $X2=0 $Y2=0
cc_338 N_A_802_323#_c_341_n N_TE_c_538_n 0.0135815f $X=7.175 $Y=1.69 $X2=0 $Y2=0
cc_339 N_A_802_323#_c_342_n N_TE_c_539_n 0.0135815f $X=7.775 $Y=1.69 $X2=0 $Y2=0
cc_340 N_A_802_323#_c_350_n TE 0.0240474f $X=8.14 $Y=1.615 $X2=0 $Y2=0
cc_341 N_A_802_323#_c_351_n TE 0.00778046f $X=7.94 $Y=2.8 $X2=0 $Y2=0
cc_342 N_A_802_323#_c_352_n TE 0.00381888f $X=8.34 $Y=0.515 $X2=0 $Y2=0
cc_343 N_A_802_323#_c_353_n N_A_27_368#_c_675_n 0.00125031f $X=4.1 $Y=1.765
+ $X2=0 $Y2=0
cc_344 N_A_802_323#_c_353_n N_A_27_368#_c_694_n 0.0057515f $X=4.1 $Y=1.765 $X2=0
+ $Y2=0
cc_345 N_A_802_323#_c_353_n N_A_27_368#_c_697_n 0.0126791f $X=4.1 $Y=1.765 $X2=0
+ $Y2=0
cc_346 N_A_802_323#_c_334_n N_A_27_368#_c_697_n 0.00359456f $X=4.475 $Y=1.69
+ $X2=0 $Y2=0
cc_347 N_A_802_323#_c_356_n N_A_27_368#_c_697_n 0.0139616f $X=4.55 $Y=1.765
+ $X2=0 $Y2=0
cc_348 N_A_802_323#_c_356_n N_A_27_368#_c_676_n 0.0048514f $X=4.55 $Y=1.765
+ $X2=0 $Y2=0
cc_349 N_A_802_323#_c_336_n N_A_27_368#_c_676_n 0.00495792f $X=4.925 $Y=1.69
+ $X2=0 $Y2=0
cc_350 N_A_802_323#_c_358_n N_A_27_368#_c_676_n 0.00460318f $X=5 $Y=1.765 $X2=0
+ $Y2=0
cc_351 N_A_802_323#_c_360_n N_A_27_368#_c_676_n 3.53158e-19 $X=5.45 $Y=1.765
+ $X2=0 $Y2=0
cc_352 N_A_802_323#_c_344_n N_A_27_368#_c_676_n 0.00119837f $X=5 $Y=1.69 $X2=0
+ $Y2=0
cc_353 N_A_802_323#_c_356_n N_A_27_368#_c_677_n 0.00578756f $X=4.55 $Y=1.765
+ $X2=0 $Y2=0
cc_354 N_A_802_323#_c_358_n N_A_27_368#_c_677_n 0.00817025f $X=5 $Y=1.765 $X2=0
+ $Y2=0
cc_355 N_A_802_323#_c_337_n N_A_27_368#_c_664_n 0.0113135f $X=5.375 $Y=1.69
+ $X2=0 $Y2=0
cc_356 N_A_802_323#_c_344_n N_A_27_368#_c_664_n 0.00779896f $X=5 $Y=1.69 $X2=0
+ $Y2=0
cc_357 N_A_802_323#_c_345_n N_A_27_368#_c_664_n 0.00779896f $X=5.45 $Y=1.69
+ $X2=0 $Y2=0
cc_358 N_A_802_323#_c_336_n N_A_27_368#_c_665_n 0.0060478f $X=4.925 $Y=1.69
+ $X2=0 $Y2=0
cc_359 N_A_802_323#_c_344_n N_A_27_368#_c_665_n 2.1146e-19 $X=5 $Y=1.69 $X2=0
+ $Y2=0
cc_360 N_A_802_323#_c_358_n N_A_27_368#_c_678_n 6.35084e-19 $X=5 $Y=1.765 $X2=0
+ $Y2=0
cc_361 N_A_802_323#_c_360_n N_A_27_368#_c_678_n 0.014764f $X=5.45 $Y=1.765 $X2=0
+ $Y2=0
cc_362 N_A_802_323#_c_338_n N_A_27_368#_c_678_n 0.00508612f $X=5.825 $Y=1.69
+ $X2=0 $Y2=0
cc_363 N_A_802_323#_c_362_n N_A_27_368#_c_678_n 0.00554458f $X=5.9 $Y=1.765
+ $X2=0 $Y2=0
cc_364 N_A_802_323#_c_345_n N_A_27_368#_c_678_n 0.00119837f $X=5.45 $Y=1.69
+ $X2=0 $Y2=0
cc_365 N_A_802_323#_c_338_n N_A_27_368#_c_666_n 0.00366668f $X=5.825 $Y=1.69
+ $X2=0 $Y2=0
cc_366 N_A_802_323#_c_339_n N_A_27_368#_c_666_n 0.00932562f $X=6.275 $Y=1.69
+ $X2=0 $Y2=0
cc_367 N_A_802_323#_c_346_n N_A_27_368#_c_666_n 0.00830203f $X=5.9 $Y=1.69 $X2=0
+ $Y2=0
cc_368 N_A_802_323#_c_347_n N_A_27_368#_c_666_n 0.00779896f $X=6.35 $Y=1.69
+ $X2=0 $Y2=0
cc_369 N_A_802_323#_c_362_n N_A_27_368#_c_679_n 6.54939e-19 $X=5.9 $Y=1.765
+ $X2=0 $Y2=0
cc_370 N_A_802_323#_c_364_n N_A_27_368#_c_679_n 0.0149123f $X=6.35 $Y=1.765
+ $X2=0 $Y2=0
cc_371 N_A_802_323#_c_340_n N_A_27_368#_c_679_n 0.00508612f $X=6.725 $Y=1.69
+ $X2=0 $Y2=0
cc_372 N_A_802_323#_c_366_n N_A_27_368#_c_679_n 0.00554458f $X=6.8 $Y=1.765
+ $X2=0 $Y2=0
cc_373 N_A_802_323#_c_347_n N_A_27_368#_c_679_n 0.00128795f $X=6.35 $Y=1.69
+ $X2=0 $Y2=0
cc_374 N_A_802_323#_c_340_n N_A_27_368#_c_667_n 0.00366668f $X=6.725 $Y=1.69
+ $X2=0 $Y2=0
cc_375 N_A_802_323#_c_341_n N_A_27_368#_c_667_n 0.00932562f $X=7.175 $Y=1.69
+ $X2=0 $Y2=0
cc_376 N_A_802_323#_c_342_n N_A_27_368#_c_667_n 0.00501819f $X=7.775 $Y=1.69
+ $X2=0 $Y2=0
cc_377 N_A_802_323#_c_348_n N_A_27_368#_c_667_n 0.00830203f $X=6.8 $Y=1.69 $X2=0
+ $Y2=0
cc_378 N_A_802_323#_c_349_n N_A_27_368#_c_667_n 0.00801042f $X=7.25 $Y=1.69
+ $X2=0 $Y2=0
cc_379 N_A_802_323#_c_350_n N_A_27_368#_c_667_n 0.00259598f $X=8.14 $Y=1.615
+ $X2=0 $Y2=0
cc_380 N_A_802_323#_c_351_n N_A_27_368#_c_667_n 0.00712759f $X=7.94 $Y=2.8 $X2=0
+ $Y2=0
cc_381 N_A_802_323#_c_366_n N_A_27_368#_c_680_n 6.54939e-19 $X=6.8 $Y=1.765
+ $X2=0 $Y2=0
cc_382 N_A_802_323#_c_368_n N_A_27_368#_c_680_n 0.0153683f $X=7.25 $Y=1.765
+ $X2=0 $Y2=0
cc_383 N_A_802_323#_c_342_n N_A_27_368#_c_680_n 0.0051257f $X=7.775 $Y=1.69
+ $X2=0 $Y2=0
cc_384 N_A_802_323#_c_349_n N_A_27_368#_c_680_n 0.00128795f $X=7.25 $Y=1.69
+ $X2=0 $Y2=0
cc_385 N_A_802_323#_c_377_n N_A_27_368#_c_680_n 0.00471029f $X=7.94 $Y=1.78
+ $X2=0 $Y2=0
cc_386 N_A_802_323#_c_351_n N_A_27_368#_c_680_n 0.0840207f $X=7.94 $Y=2.8 $X2=0
+ $Y2=0
cc_387 N_A_802_323#_c_358_n N_A_27_368#_c_739_n 0.00205171f $X=5 $Y=1.765 $X2=0
+ $Y2=0
cc_388 N_A_802_323#_c_338_n N_A_27_368#_c_668_n 0.00329878f $X=5.825 $Y=1.69
+ $X2=0 $Y2=0
cc_389 N_A_802_323#_c_345_n N_A_27_368#_c_668_n 2.1146e-19 $X=5.45 $Y=1.69 $X2=0
+ $Y2=0
cc_390 N_A_802_323#_c_340_n N_A_27_368#_c_669_n 0.00329878f $X=6.725 $Y=1.69
+ $X2=0 $Y2=0
cc_391 N_A_802_323#_c_347_n N_A_27_368#_c_669_n 2.1146e-19 $X=6.35 $Y=1.69 $X2=0
+ $Y2=0
cc_392 N_A_802_323#_c_353_n N_Z_c_866_n 7.39283e-19 $X=4.1 $Y=1.765 $X2=0 $Y2=0
cc_393 N_A_802_323#_c_353_n Z 0.00588952f $X=4.1 $Y=1.765 $X2=0 $Y2=0
cc_394 N_A_802_323#_c_334_n Z 0.00444898f $X=4.475 $Y=1.69 $X2=0 $Y2=0
cc_395 N_A_802_323#_c_335_n Z 0.00686281f $X=4.175 $Y=1.69 $X2=0 $Y2=0
cc_396 N_A_802_323#_c_356_n Z 8.3084e-19 $X=4.55 $Y=1.765 $X2=0 $Y2=0
cc_397 N_A_802_323#_c_353_n N_VPWR_c_958_n 0.00923031f $X=4.1 $Y=1.765 $X2=0
+ $Y2=0
cc_398 N_A_802_323#_c_356_n N_VPWR_c_958_n 0.0100415f $X=4.55 $Y=1.765 $X2=0
+ $Y2=0
cc_399 N_A_802_323#_c_358_n N_VPWR_c_958_n 5.32848e-19 $X=5 $Y=1.765 $X2=0 $Y2=0
cc_400 N_A_802_323#_c_358_n N_VPWR_c_959_n 0.00492639f $X=5 $Y=1.765 $X2=0 $Y2=0
cc_401 N_A_802_323#_c_337_n N_VPWR_c_959_n 0.00253179f $X=5.375 $Y=1.69 $X2=0
+ $Y2=0
cc_402 N_A_802_323#_c_360_n N_VPWR_c_959_n 0.00492882f $X=5.45 $Y=1.765 $X2=0
+ $Y2=0
cc_403 N_A_802_323#_c_360_n N_VPWR_c_960_n 0.00445602f $X=5.45 $Y=1.765 $X2=0
+ $Y2=0
cc_404 N_A_802_323#_c_362_n N_VPWR_c_960_n 0.00413917f $X=5.9 $Y=1.765 $X2=0
+ $Y2=0
cc_405 N_A_802_323#_c_360_n N_VPWR_c_961_n 7.01758e-19 $X=5.45 $Y=1.765 $X2=0
+ $Y2=0
cc_406 N_A_802_323#_c_362_n N_VPWR_c_961_n 0.0148284f $X=5.9 $Y=1.765 $X2=0
+ $Y2=0
cc_407 N_A_802_323#_c_339_n N_VPWR_c_961_n 0.00253179f $X=6.275 $Y=1.69 $X2=0
+ $Y2=0
cc_408 N_A_802_323#_c_364_n N_VPWR_c_961_n 0.00533258f $X=6.35 $Y=1.765 $X2=0
+ $Y2=0
cc_409 N_A_802_323#_c_364_n N_VPWR_c_962_n 7.01758e-19 $X=6.35 $Y=1.765 $X2=0
+ $Y2=0
cc_410 N_A_802_323#_c_366_n N_VPWR_c_962_n 0.0148284f $X=6.8 $Y=1.765 $X2=0
+ $Y2=0
cc_411 N_A_802_323#_c_341_n N_VPWR_c_962_n 0.00253179f $X=7.175 $Y=1.69 $X2=0
+ $Y2=0
cc_412 N_A_802_323#_c_368_n N_VPWR_c_962_n 0.00664113f $X=7.25 $Y=1.765 $X2=0
+ $Y2=0
cc_413 N_A_802_323#_c_351_n N_VPWR_c_964_n 0.0825826f $X=7.94 $Y=2.8 $X2=0 $Y2=0
cc_414 N_A_802_323#_c_353_n N_VPWR_c_965_n 0.00413917f $X=4.1 $Y=1.765 $X2=0
+ $Y2=0
cc_415 N_A_802_323#_c_356_n N_VPWR_c_967_n 0.00413917f $X=4.55 $Y=1.765 $X2=0
+ $Y2=0
cc_416 N_A_802_323#_c_358_n N_VPWR_c_967_n 0.00445602f $X=5 $Y=1.765 $X2=0 $Y2=0
cc_417 N_A_802_323#_c_364_n N_VPWR_c_969_n 0.00445602f $X=6.35 $Y=1.765 $X2=0
+ $Y2=0
cc_418 N_A_802_323#_c_366_n N_VPWR_c_969_n 0.00413917f $X=6.8 $Y=1.765 $X2=0
+ $Y2=0
cc_419 N_A_802_323#_c_368_n N_VPWR_c_970_n 0.00445602f $X=7.25 $Y=1.765 $X2=0
+ $Y2=0
cc_420 N_A_802_323#_c_377_n N_VPWR_c_970_n 0.00182254f $X=7.94 $Y=1.78 $X2=0
+ $Y2=0
cc_421 N_A_802_323#_c_351_n N_VPWR_c_970_n 0.0330759f $X=7.94 $Y=2.8 $X2=0 $Y2=0
cc_422 N_A_802_323#_c_353_n N_VPWR_c_957_n 0.0081781f $X=4.1 $Y=1.765 $X2=0
+ $Y2=0
cc_423 N_A_802_323#_c_356_n N_VPWR_c_957_n 0.00817726f $X=4.55 $Y=1.765 $X2=0
+ $Y2=0
cc_424 N_A_802_323#_c_358_n N_VPWR_c_957_n 0.00857589f $X=5 $Y=1.765 $X2=0 $Y2=0
cc_425 N_A_802_323#_c_360_n N_VPWR_c_957_n 0.00857589f $X=5.45 $Y=1.765 $X2=0
+ $Y2=0
cc_426 N_A_802_323#_c_362_n N_VPWR_c_957_n 0.00817726f $X=5.9 $Y=1.765 $X2=0
+ $Y2=0
cc_427 N_A_802_323#_c_364_n N_VPWR_c_957_n 0.00857589f $X=6.35 $Y=1.765 $X2=0
+ $Y2=0
cc_428 N_A_802_323#_c_366_n N_VPWR_c_957_n 0.00817726f $X=6.8 $Y=1.765 $X2=0
+ $Y2=0
cc_429 N_A_802_323#_c_368_n N_VPWR_c_957_n 0.00862391f $X=7.25 $Y=1.765 $X2=0
+ $Y2=0
cc_430 N_A_802_323#_c_351_n N_VPWR_c_957_n 0.0286723f $X=7.94 $Y=2.8 $X2=0 $Y2=0
cc_431 N_A_802_323#_c_334_n N_A_27_74#_c_1075_n 0.0100464f $X=4.475 $Y=1.69
+ $X2=0 $Y2=0
cc_432 N_A_802_323#_c_336_n N_A_27_74#_c_1075_n 5.53729e-19 $X=4.925 $Y=1.69
+ $X2=0 $Y2=0
cc_433 N_A_802_323#_c_334_n N_A_27_74#_c_1076_n 0.00135362f $X=4.475 $Y=1.69
+ $X2=0 $Y2=0
cc_434 N_A_802_323#_c_335_n N_A_27_74#_c_1076_n 9.19439e-19 $X=4.175 $Y=1.69
+ $X2=0 $Y2=0
cc_435 N_A_802_323#_c_337_n N_A_27_74#_c_1078_n 0.00178447f $X=5.375 $Y=1.69
+ $X2=0 $Y2=0
cc_436 N_A_802_323#_c_339_n N_A_27_74#_c_1080_n 0.00178512f $X=6.275 $Y=1.69
+ $X2=0 $Y2=0
cc_437 N_A_802_323#_c_341_n N_A_27_74#_c_1082_n 0.00156528f $X=7.175 $Y=1.69
+ $X2=0 $Y2=0
cc_438 N_A_802_323#_c_342_n N_A_27_74#_c_1082_n 0.00548254f $X=7.775 $Y=1.69
+ $X2=0 $Y2=0
cc_439 N_A_802_323#_c_350_n N_A_27_74#_c_1082_n 0.0131155f $X=8.14 $Y=1.615
+ $X2=0 $Y2=0
cc_440 N_A_802_323#_c_351_n N_A_27_74#_c_1082_n 0.00768298f $X=7.94 $Y=2.8 $X2=0
+ $Y2=0
cc_441 N_A_802_323#_c_352_n N_A_27_74#_c_1083_n 0.0705816f $X=8.34 $Y=0.515
+ $X2=0 $Y2=0
cc_442 N_A_802_323#_c_336_n N_A_27_74#_c_1087_n 8.34684e-19 $X=4.925 $Y=1.69
+ $X2=0 $Y2=0
cc_443 N_A_802_323#_c_346_n N_A_27_74#_c_1088_n 5.66069e-19 $X=5.9 $Y=1.69 $X2=0
+ $Y2=0
cc_444 N_A_802_323#_c_340_n N_A_27_74#_c_1089_n 8.32109e-19 $X=6.725 $Y=1.69
+ $X2=0 $Y2=0
cc_445 N_A_802_323#_c_352_n N_VGND_c_1245_n 0.0267305f $X=8.34 $Y=0.515 $X2=0
+ $Y2=0
cc_446 N_A_802_323#_c_352_n N_VGND_c_1251_n 0.0198916f $X=8.34 $Y=0.515 $X2=0
+ $Y2=0
cc_447 N_A_802_323#_c_352_n N_VGND_c_1255_n 0.0164199f $X=8.34 $Y=0.515 $X2=0
+ $Y2=0
cc_448 N_TE_c_515_n N_A_27_368#_c_697_n 3.68831e-19 $X=4.78 $Y=1.295 $X2=0 $Y2=0
cc_449 N_TE_c_516_n N_A_27_368#_c_697_n 3.73472e-19 $X=4.43 $Y=1.295 $X2=0 $Y2=0
cc_450 N_TE_c_518_n N_A_27_368#_c_664_n 0.00168303f $X=5.21 $Y=1.295 $X2=0 $Y2=0
cc_451 N_TE_c_515_n N_A_27_368#_c_665_n 9.49246e-19 $X=4.78 $Y=1.295 $X2=0 $Y2=0
cc_452 N_TE_c_535_n N_A_27_368#_c_666_n 0.00192358f $X=5.715 $Y=1.295 $X2=0
+ $Y2=0
cc_453 N_TE_c_526_n N_A_27_368#_c_667_n 0.00192473f $X=6.93 $Y=1.295 $X2=0 $Y2=0
cc_454 N_TE_c_528_n N_A_27_368#_c_667_n 9.48235e-19 $X=7.43 $Y=1.295 $X2=0 $Y2=0
cc_455 N_TE_c_520_n N_A_27_368#_c_668_n 9.48557e-19 $X=5.64 $Y=1.295 $X2=0 $Y2=0
cc_456 N_TE_c_524_n N_A_27_368#_c_669_n 9.46462e-19 $X=6.5 $Y=1.295 $X2=0 $Y2=0
cc_457 N_TE_c_532_n N_VPWR_c_964_n 0.0100734f $X=8.625 $Y=1.765 $X2=0 $Y2=0
cc_458 TE N_VPWR_c_964_n 0.0107485f $X=8.795 $Y=1.21 $X2=0 $Y2=0
cc_459 N_TE_c_532_n N_VPWR_c_970_n 0.00444469f $X=8.625 $Y=1.765 $X2=0 $Y2=0
cc_460 N_TE_c_532_n N_VPWR_c_957_n 0.00862183f $X=8.625 $Y=1.765 $X2=0 $Y2=0
cc_461 N_TE_c_514_n N_A_27_74#_c_1073_n 9.48753e-19 $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_462 N_TE_c_514_n N_A_27_74#_c_1074_n 0.00259974f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_463 N_TE_c_514_n N_A_27_74#_c_1075_n 0.00620031f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_464 N_TE_c_515_n N_A_27_74#_c_1075_n 0.00808852f $X=4.78 $Y=1.295 $X2=0 $Y2=0
cc_465 N_TE_c_516_n N_A_27_74#_c_1075_n 0.00382439f $X=4.43 $Y=1.295 $X2=0 $Y2=0
cc_466 N_TE_c_517_n N_A_27_74#_c_1075_n 0.00569215f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_467 N_TE_c_533_n N_A_27_74#_c_1075_n 0.00203633f $X=4.855 $Y=1.295 $X2=0
+ $Y2=0
cc_468 N_TE_c_514_n N_A_27_74#_c_1077_n 8.24514e-19 $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_469 N_TE_c_517_n N_A_27_74#_c_1077_n 0.0120759f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_470 N_TE_c_519_n N_A_27_74#_c_1077_n 0.00292368f $X=5.285 $Y=1.22 $X2=0 $Y2=0
cc_471 N_TE_c_518_n N_A_27_74#_c_1078_n 8.70366e-19 $X=5.21 $Y=1.295 $X2=0 $Y2=0
cc_472 N_TE_c_519_n N_A_27_74#_c_1078_n 0.00620454f $X=5.285 $Y=1.22 $X2=0 $Y2=0
cc_473 N_TE_c_520_n N_A_27_74#_c_1078_n 0.00596159f $X=5.64 $Y=1.295 $X2=0 $Y2=0
cc_474 N_TE_c_521_n N_A_27_74#_c_1078_n 0.00620454f $X=5.715 $Y=1.22 $X2=0 $Y2=0
cc_475 N_TE_c_522_n N_A_27_74#_c_1078_n 8.70366e-19 $X=6.07 $Y=1.295 $X2=0 $Y2=0
cc_476 N_TE_c_534_n N_A_27_74#_c_1078_n 0.0024633f $X=5.285 $Y=1.295 $X2=0 $Y2=0
cc_477 N_TE_c_535_n N_A_27_74#_c_1078_n 0.0024633f $X=5.715 $Y=1.295 $X2=0 $Y2=0
cc_478 N_TE_c_521_n N_A_27_74#_c_1079_n 0.00273953f $X=5.715 $Y=1.22 $X2=0 $Y2=0
cc_479 N_TE_c_523_n N_A_27_74#_c_1079_n 0.00273953f $X=6.145 $Y=1.22 $X2=0 $Y2=0
cc_480 N_TE_c_522_n N_A_27_74#_c_1080_n 8.70366e-19 $X=6.07 $Y=1.295 $X2=0 $Y2=0
cc_481 N_TE_c_523_n N_A_27_74#_c_1080_n 0.00620454f $X=6.145 $Y=1.22 $X2=0 $Y2=0
cc_482 N_TE_c_524_n N_A_27_74#_c_1080_n 0.00596159f $X=6.5 $Y=1.295 $X2=0 $Y2=0
cc_483 N_TE_c_525_n N_A_27_74#_c_1080_n 0.00620454f $X=6.575 $Y=1.22 $X2=0 $Y2=0
cc_484 N_TE_c_526_n N_A_27_74#_c_1080_n 8.70366e-19 $X=6.93 $Y=1.295 $X2=0 $Y2=0
cc_485 N_TE_c_536_n N_A_27_74#_c_1080_n 0.0024633f $X=6.145 $Y=1.295 $X2=0 $Y2=0
cc_486 N_TE_c_537_n N_A_27_74#_c_1080_n 0.0024633f $X=6.575 $Y=1.295 $X2=0 $Y2=0
cc_487 N_TE_c_525_n N_A_27_74#_c_1081_n 0.00292368f $X=6.575 $Y=1.22 $X2=0 $Y2=0
cc_488 N_TE_c_527_n N_A_27_74#_c_1081_n 0.0120759f $X=7.005 $Y=1.22 $X2=0 $Y2=0
cc_489 N_TE_c_529_n N_A_27_74#_c_1081_n 8.24514e-19 $X=7.505 $Y=1.22 $X2=0 $Y2=0
cc_490 N_TE_c_527_n N_A_27_74#_c_1082_n 0.00569215f $X=7.005 $Y=1.22 $X2=0 $Y2=0
cc_491 N_TE_c_528_n N_A_27_74#_c_1082_n 0.00808852f $X=7.43 $Y=1.295 $X2=0 $Y2=0
cc_492 N_TE_c_529_n N_A_27_74#_c_1082_n 0.00628935f $X=7.505 $Y=1.22 $X2=0 $Y2=0
cc_493 N_TE_c_530_n N_A_27_74#_c_1082_n 0.0123389f $X=8.435 $Y=1.295 $X2=0 $Y2=0
cc_494 N_TE_c_538_n N_A_27_74#_c_1082_n 0.00203633f $X=7.005 $Y=1.295 $X2=0
+ $Y2=0
cc_495 N_TE_c_539_n N_A_27_74#_c_1082_n 0.0024633f $X=7.505 $Y=1.295 $X2=0 $Y2=0
cc_496 N_TE_c_529_n N_A_27_74#_c_1083_n 0.00561403f $X=7.505 $Y=1.22 $X2=0 $Y2=0
cc_497 N_TE_c_531_n N_A_27_74#_c_1083_n 7.7288e-19 $X=8.555 $Y=1.22 $X2=0 $Y2=0
cc_498 N_TE_c_518_n N_A_27_74#_c_1087_n 0.00609583f $X=5.21 $Y=1.295 $X2=0 $Y2=0
cc_499 N_TE_c_533_n N_A_27_74#_c_1087_n 4.11475e-19 $X=4.855 $Y=1.295 $X2=0
+ $Y2=0
cc_500 N_TE_c_522_n N_A_27_74#_c_1088_n 0.00520704f $X=6.07 $Y=1.295 $X2=0 $Y2=0
cc_501 N_TE_c_526_n N_A_27_74#_c_1089_n 0.00609583f $X=6.93 $Y=1.295 $X2=0 $Y2=0
cc_502 N_TE_c_538_n N_A_27_74#_c_1089_n 4.11475e-19 $X=7.005 $Y=1.295 $X2=0
+ $Y2=0
cc_503 N_TE_c_514_n N_VGND_c_1240_n 0.0110591f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_504 N_TE_c_515_n N_VGND_c_1240_n 0.00132661f $X=4.78 $Y=1.295 $X2=0 $Y2=0
cc_505 N_TE_c_517_n N_VGND_c_1240_n 0.00528159f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_506 N_TE_c_517_n N_VGND_c_1241_n 5.77505e-19 $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_507 N_TE_c_519_n N_VGND_c_1241_n 0.0118161f $X=5.285 $Y=1.22 $X2=0 $Y2=0
cc_508 N_TE_c_520_n N_VGND_c_1241_n 7.80356e-19 $X=5.64 $Y=1.295 $X2=0 $Y2=0
cc_509 N_TE_c_521_n N_VGND_c_1241_n 0.0116953f $X=5.715 $Y=1.22 $X2=0 $Y2=0
cc_510 N_TE_c_523_n N_VGND_c_1241_n 5.3132e-19 $X=6.145 $Y=1.22 $X2=0 $Y2=0
cc_511 N_TE_c_521_n N_VGND_c_1242_n 5.3132e-19 $X=5.715 $Y=1.22 $X2=0 $Y2=0
cc_512 N_TE_c_523_n N_VGND_c_1242_n 0.0116953f $X=6.145 $Y=1.22 $X2=0 $Y2=0
cc_513 N_TE_c_524_n N_VGND_c_1242_n 7.80356e-19 $X=6.5 $Y=1.295 $X2=0 $Y2=0
cc_514 N_TE_c_525_n N_VGND_c_1242_n 0.0118161f $X=6.575 $Y=1.22 $X2=0 $Y2=0
cc_515 N_TE_c_527_n N_VGND_c_1242_n 5.77505e-19 $X=7.005 $Y=1.22 $X2=0 $Y2=0
cc_516 N_TE_c_527_n N_VGND_c_1243_n 0.00528159f $X=7.005 $Y=1.22 $X2=0 $Y2=0
cc_517 N_TE_c_528_n N_VGND_c_1243_n 0.00132661f $X=7.43 $Y=1.295 $X2=0 $Y2=0
cc_518 N_TE_c_529_n N_VGND_c_1243_n 0.0148634f $X=7.505 $Y=1.22 $X2=0 $Y2=0
cc_519 N_TE_c_531_n N_VGND_c_1245_n 0.00495522f $X=8.555 $Y=1.22 $X2=0 $Y2=0
cc_520 N_TE_c_532_n N_VGND_c_1245_n 5.98351e-19 $X=8.625 $Y=1.765 $X2=0 $Y2=0
cc_521 TE N_VGND_c_1245_n 0.0217001f $X=8.795 $Y=1.21 $X2=0 $Y2=0
cc_522 N_TE_c_521_n N_VGND_c_1246_n 0.00383152f $X=5.715 $Y=1.22 $X2=0 $Y2=0
cc_523 N_TE_c_523_n N_VGND_c_1246_n 0.00383152f $X=6.145 $Y=1.22 $X2=0 $Y2=0
cc_524 N_TE_c_514_n N_VGND_c_1248_n 0.00383152f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_525 N_TE_c_517_n N_VGND_c_1249_n 0.00434272f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_526 N_TE_c_519_n N_VGND_c_1249_n 0.00383152f $X=5.285 $Y=1.22 $X2=0 $Y2=0
cc_527 N_TE_c_525_n N_VGND_c_1250_n 0.00383152f $X=6.575 $Y=1.22 $X2=0 $Y2=0
cc_528 N_TE_c_527_n N_VGND_c_1250_n 0.00434272f $X=7.005 $Y=1.22 $X2=0 $Y2=0
cc_529 N_TE_c_529_n N_VGND_c_1251_n 0.00383152f $X=7.505 $Y=1.22 $X2=0 $Y2=0
cc_530 N_TE_c_531_n N_VGND_c_1251_n 0.00434272f $X=8.555 $Y=1.22 $X2=0 $Y2=0
cc_531 N_TE_c_514_n N_VGND_c_1255_n 0.00757637f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_532 N_TE_c_517_n N_VGND_c_1255_n 0.00820718f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_533 N_TE_c_519_n N_VGND_c_1255_n 0.0075754f $X=5.285 $Y=1.22 $X2=0 $Y2=0
cc_534 N_TE_c_521_n N_VGND_c_1255_n 0.0075754f $X=5.715 $Y=1.22 $X2=0 $Y2=0
cc_535 N_TE_c_523_n N_VGND_c_1255_n 0.0075754f $X=6.145 $Y=1.22 $X2=0 $Y2=0
cc_536 N_TE_c_525_n N_VGND_c_1255_n 0.0075754f $X=6.575 $Y=1.22 $X2=0 $Y2=0
cc_537 N_TE_c_527_n N_VGND_c_1255_n 0.00820718f $X=7.005 $Y=1.22 $X2=0 $Y2=0
cc_538 N_TE_c_529_n N_VGND_c_1255_n 0.00762539f $X=7.505 $Y=1.22 $X2=0 $Y2=0
cc_539 N_TE_c_531_n N_VGND_c_1255_n 0.00828933f $X=8.555 $Y=1.22 $X2=0 $Y2=0
cc_540 N_A_27_368#_c_671_n N_Z_M1000_s 0.00197722f $X=1.07 $Y=2.99 $X2=0 $Y2=0
cc_541 N_A_27_368#_c_673_n N_Z_M1010_s 0.00197722f $X=1.97 $Y=2.99 $X2=0 $Y2=0
cc_542 N_A_27_368#_c_674_n N_Z_M1021_s 0.00197722f $X=2.875 $Y=2.99 $X2=0 $Y2=0
cc_543 N_A_27_368#_c_675_n N_Z_M1025_s 0.00197722f $X=3.79 $Y=2.99 $X2=0 $Y2=0
cc_544 N_A_27_368#_c_671_n N_Z_c_836_n 0.0160777f $X=1.07 $Y=2.99 $X2=0 $Y2=0
cc_545 N_A_27_368#_M1003_d N_Z_c_829_n 0.00197722f $X=1.025 $Y=1.84 $X2=0 $Y2=0
cc_546 N_A_27_368#_c_759_p N_Z_c_829_n 0.0151327f $X=1.175 $Y=2.225 $X2=0 $Y2=0
cc_547 N_A_27_368#_c_670_n N_Z_c_830_n 0.00347751f $X=0.275 $Y=1.985 $X2=0 $Y2=0
cc_548 N_A_27_368#_c_673_n N_Z_c_847_n 0.0160777f $X=1.97 $Y=2.99 $X2=0 $Y2=0
cc_549 N_A_27_368#_M1018_d N_Z_c_831_n 0.00197722f $X=1.925 $Y=1.84 $X2=0 $Y2=0
cc_550 N_A_27_368#_c_763_p N_Z_c_831_n 0.0151327f $X=2.075 $Y=2.225 $X2=0 $Y2=0
cc_551 N_A_27_368#_c_674_n N_Z_c_855_n 0.0160777f $X=2.875 $Y=2.99 $X2=0 $Y2=0
cc_552 N_A_27_368#_M1022_d N_Z_c_832_n 0.00197722f $X=2.825 $Y=1.84 $X2=0 $Y2=0
cc_553 N_A_27_368#_c_766_p N_Z_c_832_n 0.0151327f $X=2.975 $Y=2.225 $X2=0 $Y2=0
cc_554 N_A_27_368#_c_675_n N_Z_c_866_n 0.0160777f $X=3.79 $Y=2.99 $X2=0 $Y2=0
cc_555 N_A_27_368#_c_693_n N_Z_c_866_n 0.0123817f $X=3.875 $Y=2.23 $X2=0 $Y2=0
cc_556 N_A_27_368#_c_694_n N_Z_c_866_n 0.0328619f $X=3.875 $Y=2.905 $X2=0 $Y2=0
cc_557 N_A_27_368#_M1031_d Z 0.00230936f $X=3.725 $Y=1.84 $X2=0 $Y2=0
cc_558 N_A_27_368#_c_693_n Z 0.0149531f $X=3.875 $Y=2.23 $X2=0 $Y2=0
cc_559 N_A_27_368#_c_697_n Z 0.011339f $X=4.69 $Y=2.145 $X2=0 $Y2=0
cc_560 N_A_27_368#_c_676_n Z 0.00537822f $X=4.775 $Y=1.985 $X2=0 $Y2=0
cc_561 N_A_27_368#_c_665_n Z 0.00643084f $X=4.94 $Y=1.635 $X2=0 $Y2=0
cc_562 N_A_27_368#_c_697_n N_VPWR_M1001_s 0.00536623f $X=4.69 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_563 N_A_27_368#_c_675_n N_VPWR_c_958_n 0.0125885f $X=3.79 $Y=2.99 $X2=0 $Y2=0
cc_564 N_A_27_368#_c_694_n N_VPWR_c_958_n 0.0328619f $X=3.875 $Y=2.905 $X2=0
+ $Y2=0
cc_565 N_A_27_368#_c_697_n N_VPWR_c_958_n 0.0171814f $X=4.69 $Y=2.145 $X2=0
+ $Y2=0
cc_566 N_A_27_368#_c_677_n N_VPWR_c_958_n 0.0389192f $X=4.775 $Y=2.4 $X2=0 $Y2=0
cc_567 N_A_27_368#_c_676_n N_VPWR_c_959_n 0.0108084f $X=4.775 $Y=1.985 $X2=0
+ $Y2=0
cc_568 N_A_27_368#_c_677_n N_VPWR_c_959_n 0.0478192f $X=4.775 $Y=2.4 $X2=0 $Y2=0
cc_569 N_A_27_368#_c_664_n N_VPWR_c_959_n 0.0132604f $X=5.51 $Y=1.635 $X2=0
+ $Y2=0
cc_570 N_A_27_368#_c_678_n N_VPWR_c_959_n 0.0695307f $X=5.675 $Y=1.985 $X2=0
+ $Y2=0
cc_571 N_A_27_368#_c_739_n N_VPWR_c_959_n 0.0117758f $X=4.815 $Y=2.145 $X2=0
+ $Y2=0
cc_572 N_A_27_368#_c_678_n N_VPWR_c_960_n 0.0110241f $X=5.675 $Y=1.985 $X2=0
+ $Y2=0
cc_573 N_A_27_368#_c_678_n N_VPWR_c_961_n 0.0716194f $X=5.675 $Y=1.985 $X2=0
+ $Y2=0
cc_574 N_A_27_368#_c_666_n N_VPWR_c_961_n 0.016902f $X=6.41 $Y=1.635 $X2=0 $Y2=0
cc_575 N_A_27_368#_c_679_n N_VPWR_c_961_n 0.0716194f $X=6.575 $Y=1.985 $X2=0
+ $Y2=0
cc_576 N_A_27_368#_c_679_n N_VPWR_c_962_n 0.0716194f $X=6.575 $Y=1.985 $X2=0
+ $Y2=0
cc_577 N_A_27_368#_c_667_n N_VPWR_c_962_n 0.016902f $X=7.31 $Y=1.635 $X2=0 $Y2=0
cc_578 N_A_27_368#_c_680_n N_VPWR_c_962_n 0.0716194f $X=7.475 $Y=1.985 $X2=0
+ $Y2=0
cc_579 N_A_27_368#_c_671_n N_VPWR_c_965_n 0.0438391f $X=1.07 $Y=2.99 $X2=0 $Y2=0
cc_580 N_A_27_368#_c_672_n N_VPWR_c_965_n 0.018997f $X=0.375 $Y=2.99 $X2=0 $Y2=0
cc_581 N_A_27_368#_c_673_n N_VPWR_c_965_n 0.0438391f $X=1.97 $Y=2.99 $X2=0 $Y2=0
cc_582 N_A_27_368#_c_674_n N_VPWR_c_965_n 0.043195f $X=2.875 $Y=2.99 $X2=0 $Y2=0
cc_583 N_A_27_368#_c_675_n N_VPWR_c_965_n 0.0573142f $X=3.79 $Y=2.99 $X2=0 $Y2=0
cc_584 N_A_27_368#_c_681_n N_VPWR_c_965_n 0.0146958f $X=1.172 $Y=2.99 $X2=0
+ $Y2=0
cc_585 N_A_27_368#_c_682_n N_VPWR_c_965_n 0.0157711f $X=2.08 $Y=2.99 $X2=0 $Y2=0
cc_586 N_A_27_368#_c_683_n N_VPWR_c_965_n 0.0143373f $X=2.975 $Y=2.99 $X2=0
+ $Y2=0
cc_587 N_A_27_368#_c_677_n N_VPWR_c_967_n 0.0110241f $X=4.775 $Y=2.4 $X2=0 $Y2=0
cc_588 N_A_27_368#_c_679_n N_VPWR_c_969_n 0.0110241f $X=6.575 $Y=1.985 $X2=0
+ $Y2=0
cc_589 N_A_27_368#_c_680_n N_VPWR_c_970_n 0.0110241f $X=7.475 $Y=1.985 $X2=0
+ $Y2=0
cc_590 N_A_27_368#_c_671_n N_VPWR_c_957_n 0.0247572f $X=1.07 $Y=2.99 $X2=0 $Y2=0
cc_591 N_A_27_368#_c_672_n N_VPWR_c_957_n 0.0103026f $X=0.375 $Y=2.99 $X2=0
+ $Y2=0
cc_592 N_A_27_368#_c_673_n N_VPWR_c_957_n 0.0247572f $X=1.97 $Y=2.99 $X2=0 $Y2=0
cc_593 N_A_27_368#_c_674_n N_VPWR_c_957_n 0.0243813f $X=2.875 $Y=2.99 $X2=0
+ $Y2=0
cc_594 N_A_27_368#_c_675_n N_VPWR_c_957_n 0.0321184f $X=3.79 $Y=2.99 $X2=0 $Y2=0
cc_595 N_A_27_368#_c_677_n N_VPWR_c_957_n 0.00909194f $X=4.775 $Y=2.4 $X2=0
+ $Y2=0
cc_596 N_A_27_368#_c_678_n N_VPWR_c_957_n 0.00909194f $X=5.675 $Y=1.985 $X2=0
+ $Y2=0
cc_597 N_A_27_368#_c_679_n N_VPWR_c_957_n 0.00909194f $X=6.575 $Y=1.985 $X2=0
+ $Y2=0
cc_598 N_A_27_368#_c_680_n N_VPWR_c_957_n 0.00909194f $X=7.475 $Y=1.985 $X2=0
+ $Y2=0
cc_599 N_A_27_368#_c_681_n N_VPWR_c_957_n 0.00796993f $X=1.172 $Y=2.99 $X2=0
+ $Y2=0
cc_600 N_A_27_368#_c_682_n N_VPWR_c_957_n 0.00855309f $X=2.08 $Y=2.99 $X2=0
+ $Y2=0
cc_601 N_A_27_368#_c_683_n N_VPWR_c_957_n 0.00777554f $X=2.975 $Y=2.99 $X2=0
+ $Y2=0
cc_602 N_A_27_368#_c_665_n N_A_27_74#_c_1075_n 0.018115f $X=4.94 $Y=1.635 $X2=0
+ $Y2=0
cc_603 N_A_27_368#_c_664_n N_A_27_74#_c_1078_n 0.0266476f $X=5.51 $Y=1.635 $X2=0
+ $Y2=0
cc_604 N_A_27_368#_c_666_n N_A_27_74#_c_1078_n 0.00632315f $X=6.41 $Y=1.635
+ $X2=0 $Y2=0
cc_605 N_A_27_368#_c_668_n N_A_27_74#_c_1078_n 0.0211079f $X=5.635 $Y=1.635
+ $X2=0 $Y2=0
cc_606 N_A_27_368#_c_666_n N_A_27_74#_c_1080_n 0.0296586f $X=6.41 $Y=1.635 $X2=0
+ $Y2=0
cc_607 N_A_27_368#_c_667_n N_A_27_74#_c_1080_n 0.00331213f $X=7.31 $Y=1.635
+ $X2=0 $Y2=0
cc_608 N_A_27_368#_c_669_n N_A_27_74#_c_1080_n 0.0211079f $X=6.535 $Y=1.635
+ $X2=0 $Y2=0
cc_609 N_A_27_368#_c_667_n N_A_27_74#_c_1082_n 0.0477555f $X=7.31 $Y=1.635 $X2=0
+ $Y2=0
cc_610 N_A_27_368#_c_664_n N_A_27_74#_c_1087_n 0.0181153f $X=5.51 $Y=1.635 $X2=0
+ $Y2=0
cc_611 N_A_27_368#_c_665_n N_A_27_74#_c_1087_n 0.00327833f $X=4.94 $Y=1.635
+ $X2=0 $Y2=0
cc_612 N_A_27_368#_c_666_n N_A_27_74#_c_1088_n 0.0143536f $X=6.41 $Y=1.635 $X2=0
+ $Y2=0
cc_613 N_A_27_368#_c_667_n N_A_27_74#_c_1089_n 0.0211082f $X=7.31 $Y=1.635 $X2=0
+ $Y2=0
cc_614 N_Z_c_881_n N_A_27_74#_M1009_d 0.00462121f $X=1.545 $Y=0.812 $X2=0 $Y2=0
cc_615 N_Z_c_892_n N_A_27_74#_M1016_d 0.00462121f $X=2.545 $Y=0.812 $X2=0 $Y2=0
cc_616 N_Z_c_863_n N_A_27_74#_M1023_d 0.00462121f $X=3.545 $Y=0.925 $X2=0 $Y2=0
cc_617 N_Z_M1005_s N_A_27_74#_c_1069_n 0.00184993f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_618 N_Z_c_873_n N_A_27_74#_c_1069_n 0.0124744f $X=0.71 $Y=0.78 $X2=0 $Y2=0
cc_619 N_Z_c_881_n N_A_27_74#_c_1069_n 0.00352531f $X=1.545 $Y=0.812 $X2=0 $Y2=0
cc_620 N_Z_M1014_s N_A_27_74#_c_1071_n 0.00263602f $X=1.5 $Y=0.37 $X2=0 $Y2=0
cc_621 N_Z_c_881_n N_A_27_74#_c_1071_n 0.00352531f $X=1.545 $Y=0.812 $X2=0 $Y2=0
cc_622 N_Z_c_885_n N_A_27_74#_c_1071_n 0.0171011f $X=1.875 $Y=0.812 $X2=0 $Y2=0
cc_623 N_Z_c_892_n N_A_27_74#_c_1071_n 0.00211519f $X=2.545 $Y=0.812 $X2=0 $Y2=0
cc_624 N_Z_M1020_s N_A_27_74#_c_1072_n 0.00263602f $X=2.5 $Y=0.37 $X2=0 $Y2=0
cc_625 N_Z_c_863_n N_A_27_74#_c_1072_n 0.0035136f $X=3.545 $Y=0.925 $X2=0 $Y2=0
cc_626 N_Z_c_892_n N_A_27_74#_c_1072_n 0.0033843f $X=2.545 $Y=0.812 $X2=0 $Y2=0
cc_627 N_Z_c_895_n N_A_27_74#_c_1072_n 0.0171011f $X=2.875 $Y=0.812 $X2=0 $Y2=0
cc_628 N_Z_M1026_s N_A_27_74#_c_1073_n 0.00250873f $X=3.5 $Y=0.37 $X2=0 $Y2=0
cc_629 N_Z_c_863_n N_A_27_74#_c_1073_n 0.00352531f $X=3.545 $Y=0.925 $X2=0 $Y2=0
cc_630 N_Z_c_898_n N_A_27_74#_c_1073_n 0.0192212f $X=3.71 $Y=0.76 $X2=0 $Y2=0
cc_631 N_Z_c_898_n N_A_27_74#_c_1074_n 0.0248574f $X=3.71 $Y=0.76 $X2=0 $Y2=0
cc_632 N_Z_c_827_n N_A_27_74#_c_1076_n 0.0131434f $X=3.79 $Y=1.55 $X2=0 $Y2=0
cc_633 Z N_A_27_74#_c_1076_n 0.0124668f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_634 N_Z_c_881_n N_A_27_74#_c_1084_n 0.0197079f $X=1.545 $Y=0.812 $X2=0 $Y2=0
cc_635 N_Z_c_892_n N_A_27_74#_c_1085_n 0.0197079f $X=2.545 $Y=0.812 $X2=0 $Y2=0
cc_636 N_Z_c_863_n N_A_27_74#_c_1086_n 0.0197079f $X=3.545 $Y=0.925 $X2=0 $Y2=0
cc_637 N_Z_c_863_n N_VGND_c_1255_n 0.00142691f $X=3.545 $Y=0.925 $X2=0 $Y2=0
cc_638 N_Z_c_881_n N_VGND_c_1255_n 0.00142621f $X=1.545 $Y=0.812 $X2=0 $Y2=0
cc_639 N_Z_c_892_n N_VGND_c_1255_n 0.00114754f $X=2.545 $Y=0.812 $X2=0 $Y2=0
cc_640 N_A_27_74#_c_1073_n N_VGND_c_1240_n 0.0112234f $X=4.055 $Y=0.34 $X2=0
+ $Y2=0
cc_641 N_A_27_74#_c_1075_n N_VGND_c_1240_n 0.0238715f $X=4.905 $Y=1.295 $X2=0
+ $Y2=0
cc_642 N_A_27_74#_c_1077_n N_VGND_c_1240_n 0.0256025f $X=5.07 $Y=0.515 $X2=0
+ $Y2=0
cc_643 N_A_27_74#_c_1077_n N_VGND_c_1241_n 0.0254585f $X=5.07 $Y=0.515 $X2=0
+ $Y2=0
cc_644 N_A_27_74#_c_1078_n N_VGND_c_1241_n 0.0216086f $X=5.845 $Y=1.295 $X2=0
+ $Y2=0
cc_645 N_A_27_74#_c_1079_n N_VGND_c_1241_n 0.0254171f $X=5.93 $Y=0.515 $X2=0
+ $Y2=0
cc_646 N_A_27_74#_c_1079_n N_VGND_c_1242_n 0.0254171f $X=5.93 $Y=0.515 $X2=0
+ $Y2=0
cc_647 N_A_27_74#_c_1080_n N_VGND_c_1242_n 0.0216086f $X=6.705 $Y=1.295 $X2=0
+ $Y2=0
cc_648 N_A_27_74#_c_1081_n N_VGND_c_1242_n 0.0254585f $X=6.79 $Y=0.515 $X2=0
+ $Y2=0
cc_649 N_A_27_74#_c_1081_n N_VGND_c_1243_n 0.0256025f $X=6.79 $Y=0.515 $X2=0
+ $Y2=0
cc_650 N_A_27_74#_c_1082_n N_VGND_c_1243_n 0.0238715f $X=7.635 $Y=1.295 $X2=0
+ $Y2=0
cc_651 N_A_27_74#_c_1083_n N_VGND_c_1243_n 0.0254585f $X=7.72 $Y=0.515 $X2=0
+ $Y2=0
cc_652 N_A_27_74#_c_1079_n N_VGND_c_1246_n 0.00749631f $X=5.93 $Y=0.515 $X2=0
+ $Y2=0
cc_653 N_A_27_74#_c_1069_n N_VGND_c_1248_n 0.0378242f $X=1.045 $Y=0.34 $X2=0
+ $Y2=0
cc_654 N_A_27_74#_c_1070_n N_VGND_c_1248_n 0.0235688f $X=0.445 $Y=0.34 $X2=0
+ $Y2=0
cc_655 N_A_27_74#_c_1071_n N_VGND_c_1248_n 0.0423597f $X=2.045 $Y=0.34 $X2=0
+ $Y2=0
cc_656 N_A_27_74#_c_1072_n N_VGND_c_1248_n 0.0423597f $X=3.045 $Y=0.34 $X2=0
+ $Y2=0
cc_657 N_A_27_74#_c_1073_n N_VGND_c_1248_n 0.0551615f $X=4.055 $Y=0.34 $X2=0
+ $Y2=0
cc_658 N_A_27_74#_c_1084_n N_VGND_c_1248_n 0.0225845f $X=1.21 $Y=0.34 $X2=0
+ $Y2=0
cc_659 N_A_27_74#_c_1085_n N_VGND_c_1248_n 0.0225845f $X=2.21 $Y=0.34 $X2=0
+ $Y2=0
cc_660 N_A_27_74#_c_1086_n N_VGND_c_1248_n 0.0225845f $X=3.21 $Y=0.34 $X2=0
+ $Y2=0
cc_661 N_A_27_74#_c_1077_n N_VGND_c_1249_n 0.0109942f $X=5.07 $Y=0.515 $X2=0
+ $Y2=0
cc_662 N_A_27_74#_c_1081_n N_VGND_c_1250_n 0.0109942f $X=6.79 $Y=0.515 $X2=0
+ $Y2=0
cc_663 N_A_27_74#_c_1083_n N_VGND_c_1251_n 0.011066f $X=7.72 $Y=0.515 $X2=0
+ $Y2=0
cc_664 N_A_27_74#_c_1069_n N_VGND_c_1255_n 0.0213038f $X=1.045 $Y=0.34 $X2=0
+ $Y2=0
cc_665 N_A_27_74#_c_1070_n N_VGND_c_1255_n 0.0127152f $X=0.445 $Y=0.34 $X2=0
+ $Y2=0
cc_666 N_A_27_74#_c_1071_n N_VGND_c_1255_n 0.0239391f $X=2.045 $Y=0.34 $X2=0
+ $Y2=0
cc_667 N_A_27_74#_c_1072_n N_VGND_c_1255_n 0.0239391f $X=3.045 $Y=0.34 $X2=0
+ $Y2=0
cc_668 N_A_27_74#_c_1073_n N_VGND_c_1255_n 0.0309203f $X=4.055 $Y=0.34 $X2=0
+ $Y2=0
cc_669 N_A_27_74#_c_1077_n N_VGND_c_1255_n 0.00904371f $X=5.07 $Y=0.515 $X2=0
+ $Y2=0
cc_670 N_A_27_74#_c_1079_n N_VGND_c_1255_n 0.0062048f $X=5.93 $Y=0.515 $X2=0
+ $Y2=0
cc_671 N_A_27_74#_c_1081_n N_VGND_c_1255_n 0.00904371f $X=6.79 $Y=0.515 $X2=0
+ $Y2=0
cc_672 N_A_27_74#_c_1083_n N_VGND_c_1255_n 0.00915947f $X=7.72 $Y=0.515 $X2=0
+ $Y2=0
cc_673 N_A_27_74#_c_1084_n N_VGND_c_1255_n 0.0124836f $X=1.21 $Y=0.34 $X2=0
+ $Y2=0
cc_674 N_A_27_74#_c_1085_n N_VGND_c_1255_n 0.0124836f $X=2.21 $Y=0.34 $X2=0
+ $Y2=0
cc_675 N_A_27_74#_c_1086_n N_VGND_c_1255_n 0.0124836f $X=3.21 $Y=0.34 $X2=0
+ $Y2=0
