* File: sky130_fd_sc_ls__dlrtp_1.pex.spice
* Created: Wed Sep  2 11:03:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__DLRTP_1%D 2 3 5 8 10 14 15
r30 13 15 33.413 $w=3.39e-07 $l=2.35e-07 $layer=POLY_cond $X=0.27 $Y=1.54
+ $X2=0.505 $Y2=1.54
r31 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r32 10 14 8.53661 $w=2.68e-07 $l=2e-07 $layer=LI1_cond $X=0.24 $Y=1.665 $X2=0.24
+ $Y2=1.465
r33 6 15 13.5074 $w=3.39e-07 $l=2.83549e-07 $layer=POLY_cond $X=0.6 $Y=1.3
+ $X2=0.505 $Y2=1.54
r34 6 8 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.6 $Y=1.3 $X2=0.6
+ $Y2=0.835
r35 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=2.045
+ $X2=0.505 $Y2=2.54
r36 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.955 $X2=0.505
+ $Y2=2.045
r37 1 15 17.5597 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=0.505 $Y=1.78
+ $X2=0.505 $Y2=1.54
r38 1 2 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=0.505 $Y=1.78
+ $X2=0.505 $Y2=1.955
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_1%GATE 2 3 5 8 10 17
c40 8 0 7.12951e-20 $X=1.185 $Y=0.74
r41 15 17 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.095 $Y=1.615
+ $X2=1.185 $Y2=1.615
r42 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.095
+ $Y=1.615 $X2=1.095 $Y2=1.615
r43 12 15 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.005 $Y=1.615
+ $X2=1.095 $Y2=1.615
r44 10 16 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.095 $Y2=1.615
r45 6 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.45
+ $X2=1.185 $Y2=1.615
r46 6 8 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.185 $Y=1.45
+ $X2=1.185 $Y2=0.74
r47 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.005 $Y=2.045
+ $X2=1.005 $Y2=2.54
r48 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.005 $Y=1.955 $X2=1.005
+ $Y2=2.045
r49 1 12 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.78
+ $X2=1.005 $Y2=1.615
r50 1 2 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=1.005 $Y=1.78
+ $X2=1.005 $Y2=1.955
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_1%A_216_424# 1 2 7 10 11 13 16 18 20 21 22 25
+ 27 28 34 39 40 44 45 48 51 53 56 57 58 60
c149 57 0 1.3812e-19 $X=3.93 $Y=1.39
c150 56 0 6.93786e-20 $X=3.93 $Y=1.39
c151 43 0 5.47968e-20 $X=2.935 $Y=0.77
c152 22 0 1.98637e-19 $X=3.275 $Y=1.765
c153 18 0 1.76514e-19 $X=3.185 $Y=1.885
r154 56 58 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.965 $Y=1.39
+ $X2=3.965 $Y2=1.225
r155 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.93
+ $Y=1.39 $X2=3.93 $Y2=1.39
r156 52 60 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.665 $Y=1.615
+ $X2=1.665 $Y2=1.525
r157 51 54 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.642 $Y=1.615
+ $X2=1.642 $Y2=1.78
r158 51 53 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.642 $Y=1.615
+ $X2=1.642 $Y2=1.45
r159 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.665
+ $Y=1.615 $X2=1.665 $Y2=1.615
r160 49 53 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.54 $Y=1.13
+ $X2=1.54 $Y2=1.45
r161 48 49 11.8581 $w=3.88e-07 $l=2.75e-07 $layer=LI1_cond $X=1.43 $Y=0.855
+ $X2=1.43 $Y2=1.13
r162 46 58 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.92 $Y=0.425
+ $X2=3.92 $Y2=1.225
r163 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.835 $Y=0.34
+ $X2=3.92 $Y2=0.425
r164 44 45 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=3.835 $Y=0.34
+ $X2=3.02 $Y2=0.34
r165 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.935 $Y=0.425
+ $X2=3.02 $Y2=0.34
r166 42 43 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.935 $Y=0.425
+ $X2=2.935 $Y2=0.77
r167 41 48 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.625 $Y=0.855
+ $X2=1.43 $Y2=0.855
r168 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.85 $Y=0.855
+ $X2=2.935 $Y2=0.77
r169 40 41 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=2.85 $Y=0.855
+ $X2=1.625 $Y2=0.855
r170 39 54 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.54 $Y=1.97
+ $X2=1.54 $Y2=1.78
r171 32 48 2.51173 $w=3.88e-07 $l=8.5e-08 $layer=LI1_cond $X=1.43 $Y=0.77
+ $X2=1.43 $Y2=0.855
r172 32 34 7.5352 $w=3.88e-07 $l=2.55e-07 $layer=LI1_cond $X=1.43 $Y=0.77
+ $X2=1.43 $Y2=0.515
r173 28 39 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.455 $Y=2.095
+ $X2=1.54 $Y2=1.97
r174 28 30 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=1.455 $Y=2.095
+ $X2=1.355 $Y2=2.095
r175 23 57 38.6777 $w=2.84e-07 $l=2.18746e-07 $layer=POLY_cond $X=3.77 $Y=1.225
+ $X2=3.895 $Y2=1.39
r176 23 25 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.77 $Y=1.225
+ $X2=3.77 $Y2=0.58
r177 21 57 63.6444 $w=2.84e-07 $l=4.64354e-07 $layer=POLY_cond $X=3.695 $Y=1.765
+ $X2=3.895 $Y2=1.39
r178 21 22 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.695 $Y=1.765
+ $X2=3.275 $Y2=1.765
r179 18 22 26.9307 $w=1.5e-07 $l=1.58745e-07 $layer=POLY_cond $X=3.185 $Y=1.885
+ $X2=3.275 $Y2=1.765
r180 18 20 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.185 $Y=1.885
+ $X2=3.185 $Y2=2.46
r181 14 27 18.8402 $w=1.65e-07 $l=9.08295e-08 $layer=POLY_cond $X=2.24 $Y=1.45
+ $X2=2.205 $Y2=1.525
r182 14 16 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.24 $Y=1.45
+ $X2=2.24 $Y2=0.74
r183 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.185 $Y=1.885
+ $X2=2.185 $Y2=2.38
r184 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.185 $Y=1.795
+ $X2=2.185 $Y2=1.885
r185 9 27 18.8402 $w=1.65e-07 $l=8.44097e-08 $layer=POLY_cond $X=2.185 $Y=1.6
+ $X2=2.205 $Y2=1.525
r186 9 10 75.7984 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=2.185 $Y=1.6
+ $X2=2.185 $Y2=1.795
r187 8 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.525
+ $X2=1.665 $Y2=1.525
r188 7 27 6.66866 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=2.095 $Y=1.525
+ $X2=2.205 $Y2=1.525
r189 7 8 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=2.095 $Y=1.525
+ $X2=1.83 $Y2=1.525
r190 2 30 600 $w=1.7e-07 $l=2.824e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=2.12 $X2=1.355 $Y2=2.135
r191 1 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.26
+ $Y=0.37 $X2=1.4 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_1%A_27_424# 1 2 9 11 13 17 18 21 23 26 30 33
c91 33 0 1.20405e-19 $X=2.69 $Y=1.635
c92 21 0 1.2531e-19 $X=2.61 $Y=2.39
c93 11 0 1.81262e-19 $X=2.765 $Y=1.885
c94 9 0 1.71716e-19 $X=2.75 $Y=0.69
r95 33 36 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=1.635
+ $X2=2.69 $Y2=1.8
r96 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.635 $X2=2.69 $Y2=1.635
r97 28 30 4.96677 $w=5.88e-07 $l=2.45e-07 $layer=LI1_cond $X=0.385 $Y=0.835
+ $X2=0.63 $Y2=0.835
r98 25 26 7.19996 $w=4.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=2.33
+ $X2=0.715 $Y2=2.33
r99 23 25 9.1006 $w=4.58e-07 $l=3.5e-07 $layer=LI1_cond $X=0.28 $Y=2.33 $X2=0.63
+ $Y2=2.33
r100 21 36 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.61 $Y=2.39
+ $X2=2.61 $Y2=1.8
r101 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.525 $Y=2.475
+ $X2=2.61 $Y2=2.39
r102 18 26 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=2.525 $Y=2.475
+ $X2=0.715 $Y2=2.475
r103 17 25 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.63 $Y=2.1 $X2=0.63
+ $Y2=2.33
r104 16 30 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=0.63 $Y=1.13
+ $X2=0.63 $Y2=0.835
r105 16 17 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=0.63 $Y=1.13
+ $X2=0.63 $Y2=2.1
r106 11 34 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.765 $Y=1.885
+ $X2=2.69 $Y2=1.635
r107 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.765 $Y=1.885
+ $X2=2.765 $Y2=2.46
r108 7 34 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.75 $Y=1.47
+ $X2=2.69 $Y2=1.635
r109 7 9 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.75 $Y=1.47 $X2=2.75
+ $Y2=0.69
r110 2 23 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
r111 1 28 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.24
+ $Y=0.56 $X2=0.385 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_1%A_363_74# 1 2 9 10 12 14 15 16 18 20 21 22
+ 25 35 39 41 45 48
c113 45 0 1.95222e-19 $X=3.23 $Y=1.285
c114 35 0 1.81262e-19 $X=2.085 $Y=2.12
c115 25 0 1.3812e-19 $X=3.88 $Y=2.215
c116 20 0 1.90301e-19 $X=3.11 $Y=1.97
c117 16 0 7.12951e-20 $X=2.17 $Y=1.195
r118 45 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.23 $Y=1.285
+ $X2=3.23 $Y2=1.12
r119 44 46 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=1.285
+ $X2=3.175 $Y2=1.45
r120 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.23
+ $Y=1.285 $X2=3.23 $Y2=1.285
r121 41 44 3.45733 $w=2.98e-07 $l=9e-08 $layer=LI1_cond $X=3.175 $Y=1.195
+ $X2=3.175 $Y2=1.285
r122 37 39 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.99 $Y=2.055
+ $X2=3.11 $Y2=2.055
r123 33 35 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=1.96 $Y=2.12
+ $X2=2.085 $Y2=2.12
r124 29 31 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.96 $Y=1.195
+ $X2=2.085 $Y2=1.195
r125 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.88
+ $Y=2.215 $X2=3.88 $Y2=2.215
r126 23 25 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.88 $Y=2.905
+ $X2=3.88 $Y2=2.215
r127 21 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.715 $Y=2.99
+ $X2=3.88 $Y2=2.905
r128 21 22 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.715 $Y=2.99
+ $X2=3.075 $Y2=2.99
r129 20 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.11 $Y=1.97
+ $X2=3.11 $Y2=2.055
r130 20 46 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.11 $Y=1.97
+ $X2=3.11 $Y2=1.45
r131 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.99 $Y=2.905
+ $X2=3.075 $Y2=2.99
r132 17 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=2.14
+ $X2=2.99 $Y2=2.055
r133 17 18 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.99 $Y=2.14
+ $X2=2.99 $Y2=2.905
r134 16 31 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=1.195
+ $X2=2.085 $Y2=1.195
r135 15 41 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.025 $Y=1.195
+ $X2=3.175 $Y2=1.195
r136 15 16 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=3.025 $Y=1.195
+ $X2=2.17 $Y2=1.195
r137 14 35 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.085 $Y=2.02
+ $X2=2.085 $Y2=2.12
r138 13 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=1.28
+ $X2=2.085 $Y2=1.195
r139 13 14 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.085 $Y=1.28
+ $X2=2.085 $Y2=2.02
r140 10 26 50.1894 $w=3.66e-07 $l=3.02903e-07 $layer=POLY_cond $X=3.72 $Y=2.465
+ $X2=3.837 $Y2=2.215
r141 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.72 $Y=2.465
+ $X2=3.72 $Y2=2.75
r142 9 48 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.14 $Y=0.69
+ $X2=3.14 $Y2=1.12
r143 2 33 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.815
+ $Y=1.96 $X2=1.96 $Y2=2.12
r144 1 29 182 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_NDIFF $count=1 $X=1.815
+ $Y=0.37 $X2=1.96 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_1%A_817_48# 1 2 7 9 10 12 14 15 17 18 20 23 25
+ 32 38 40 44 47 49 50
c106 23 0 6.93786e-20 $X=4.38 $Y=0.94
c107 14 0 1.44303e-19 $X=4.38 $Y=2.05
r108 51 52 5.11481 $w=4.78e-07 $l=1.58e-07 $layer=LI1_cond $X=5.335 $Y=2.222
+ $X2=5.335 $Y2=2.38
r109 49 51 2.66626 $w=4.78e-07 $l=1.07e-07 $layer=LI1_cond $X=5.335 $Y=2.115
+ $X2=5.335 $Y2=2.222
r110 49 50 9.39634 $w=4.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=2.115
+ $X2=5.335 $Y2=1.95
r111 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.14
+ $Y=1.385 $X2=6.14 $Y2=1.385
r112 42 44 7.38284 $w=3.18e-07 $l=2.05e-07 $layer=LI1_cond $X=6.135 $Y=1.18
+ $X2=6.135 $Y2=1.385
r113 41 47 2.76166 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=5.265 $Y=1.095
+ $X2=5.017 $Y2=1.095
r114 40 42 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=5.975 $Y=1.095
+ $X2=6.135 $Y2=1.18
r115 40 41 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.975 $Y=1.095
+ $X2=5.265 $Y2=1.095
r116 38 52 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=2.465
+ $X2=5.41 $Y2=2.38
r117 34 47 3.70735 $w=2.5e-07 $l=2.01057e-07 $layer=LI1_cond $X=5.18 $Y=1.18
+ $X2=5.017 $Y2=1.095
r118 34 50 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.18 $Y=1.18
+ $X2=5.18 $Y2=1.95
r119 30 47 3.70735 $w=2.5e-07 $l=1.19143e-07 $layer=LI1_cond $X=4.935 $Y=1.01
+ $X2=5.017 $Y2=1.095
r120 30 32 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.935 $Y=1.01
+ $X2=4.935 $Y2=0.515
r121 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.47
+ $Y=2.215 $X2=4.47 $Y2=2.215
r122 25 51 3.21507 $w=3.15e-07 $l=2.4e-07 $layer=LI1_cond $X=5.095 $Y=2.222
+ $X2=5.335 $Y2=2.222
r123 25 27 22.8659 $w=3.13e-07 $l=6.25e-07 $layer=LI1_cond $X=5.095 $Y=2.222
+ $X2=4.47 $Y2=2.222
r124 21 23 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=4.16 $Y=0.94
+ $X2=4.38 $Y2=0.94
r125 18 45 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=6.215 $Y=1.765
+ $X2=6.14 $Y2=1.385
r126 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.215 $Y=1.765
+ $X2=6.215 $Y2=2.4
r127 15 45 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=6.05 $Y=1.22
+ $X2=6.14 $Y2=1.385
r128 15 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.05 $Y=1.22
+ $X2=6.05 $Y2=0.74
r129 14 28 38.535 $w=3.06e-07 $l=2.0106e-07 $layer=POLY_cond $X=4.38 $Y=2.05
+ $X2=4.46 $Y2=2.215
r130 13 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.38 $Y=1.015
+ $X2=4.38 $Y2=0.94
r131 13 14 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=4.38 $Y=1.015
+ $X2=4.38 $Y2=2.05
r132 10 28 51.9239 $w=3.06e-07 $l=2.89396e-07 $layer=POLY_cond $X=4.375 $Y=2.465
+ $X2=4.46 $Y2=2.215
r133 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.375 $Y=2.465
+ $X2=4.375 $Y2=2.75
r134 7 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.16 $Y=0.865
+ $X2=4.16 $Y2=0.94
r135 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.16 $Y=0.865 $X2=4.16
+ $Y2=0.58
r136 2 49 600 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=1 $X=5.21
+ $Y=1.96 $X2=5.41 $Y2=2.115
r137 2 38 300 $w=1.7e-07 $l=5.96678e-07 $layer=licon1_PDIFF $count=2 $X=5.21
+ $Y=1.96 $X2=5.41 $Y2=2.465
r138 1 32 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.79
+ $Y=0.37 $X2=4.935 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_1%A_643_74# 1 2 7 9 12 14 15 19 20 21 25 28 29
+ 35
c83 29 0 4.70777e-20 $X=3.39 $Y=2.405
c84 25 0 1.71716e-19 $X=3.58 $Y=0.76
c85 21 0 3.71736e-19 $X=3.665 $Y=1.81
c86 19 0 1.44303e-19 $X=3.58 $Y=1.725
r87 35 38 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=4.795 $Y=1.635
+ $X2=4.795 $Y2=1.81
r88 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.83
+ $Y=1.635 $X2=4.83 $Y2=1.635
r89 31 33 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.45 $Y=1.81
+ $X2=3.58 $Y2=1.81
r90 28 29 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.39 $Y=2.57
+ $X2=3.39 $Y2=2.405
r91 23 25 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=0.76
+ $X2=3.58 $Y2=0.76
r92 21 33 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.665 $Y=1.81
+ $X2=3.58 $Y2=1.81
r93 20 38 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.665 $Y=1.81
+ $X2=4.795 $Y2=1.81
r94 20 21 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=4.665 $Y=1.81
+ $X2=3.665 $Y2=1.81
r95 19 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=1.725
+ $X2=3.58 $Y2=1.81
r96 18 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.58 $Y=0.925
+ $X2=3.58 $Y2=0.76
r97 18 19 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.58 $Y=0.925 $X2=3.58
+ $Y2=1.725
r98 16 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.45 $Y=1.895
+ $X2=3.45 $Y2=1.81
r99 16 29 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.45 $Y=1.895
+ $X2=3.45 $Y2=2.405
r100 14 36 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.045 $Y=1.635
+ $X2=4.83 $Y2=1.635
r101 14 15 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=5.045 $Y=1.635
+ $X2=5.135 $Y2=1.677
r102 10 15 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=5.15 $Y=1.47
+ $X2=5.135 $Y2=1.677
r103 10 12 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=5.15 $Y=1.47
+ $X2=5.15 $Y2=0.74
r104 7 15 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.135 $Y=1.885
+ $X2=5.135 $Y2=1.677
r105 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.135 $Y=1.885
+ $X2=5.135 $Y2=2.46
r106 2 28 600 $w=1.7e-07 $l=6.80882e-07 $layer=licon1_PDIFF $count=1 $X=3.26
+ $Y=1.96 $X2=3.41 $Y2=2.57
r107 1 23 182 $w=1.7e-07 $l=4.79687e-07 $layer=licon1_NDIFF $count=1 $X=3.215
+ $Y=0.37 $X2=3.415 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_1%RESET_B 3 5 7 8 12
c36 3 0 1.77844e-19 $X=5.54 $Y=0.74
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.6
+ $Y=1.515 $X2=5.6 $Y2=1.515
r38 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=5.6 $Y=1.665 $X2=5.6
+ $Y2=1.515
r39 5 11 75.1901 $w=2.72e-07 $l=3.87105e-07 $layer=POLY_cond $X=5.635 $Y=1.885
+ $X2=5.6 $Y2=1.515
r40 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.635 $Y=1.885
+ $X2=5.635 $Y2=2.46
r41 1 11 38.8629 $w=2.72e-07 $l=1.92678e-07 $layer=POLY_cond $X=5.54 $Y=1.35
+ $X2=5.6 $Y2=1.515
r42 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.54 $Y=1.35 $X2=5.54
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_1%VPWR 1 2 3 4 15 19 23 28 29 30 32 37 45 55
+ 56 59 62 65
r75 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r76 65 68 9.62469 $w=6.38e-07 $l=5.15e-07 $layer=LI1_cond $X=4.755 $Y=2.815
+ $X2=4.755 $Y2=3.33
r77 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r78 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r80 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r81 53 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r82 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r83 50 68 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=5.075 $Y=3.33
+ $X2=4.755 $Y2=3.33
r84 50 52 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=5.075 $Y=3.33
+ $X2=5.52 $Y2=3.33
r85 49 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r86 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r87 46 62 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=2.517 $Y2=3.33
r88 46 48 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r89 45 68 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=4.435 $Y=3.33
+ $X2=4.755 $Y2=3.33
r90 45 48 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.435 $Y=3.33
+ $X2=4.08 $Y2=3.33
r91 44 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r92 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r93 41 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r94 41 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r95 40 43 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r96 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r97 38 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r98 38 40 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r99 37 62 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.517 $Y2=3.33
r100 37 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.16 $Y2=3.33
r101 35 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r103 32 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r104 32 34 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r105 30 49 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r106 30 63 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=2.64 $Y2=3.33
r107 28 52 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.745 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.745 $Y=3.33
+ $X2=5.91 $Y2=3.33
r109 27 55 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.075 $Y=3.33
+ $X2=6.48 $Y2=3.33
r110 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.075 $Y=3.33
+ $X2=5.91 $Y2=3.33
r111 23 26 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=5.91 $Y=2.115
+ $X2=5.91 $Y2=2.815
r112 21 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.91 $Y=3.245
+ $X2=5.91 $Y2=3.33
r113 21 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.91 $Y=3.245
+ $X2=5.91 $Y2=2.815
r114 17 62 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.517 $Y=3.245
+ $X2=2.517 $Y2=3.33
r115 17 19 13.2147 $w=3.73e-07 $l=4.3e-07 $layer=LI1_cond $X=2.517 $Y=3.245
+ $X2=2.517 $Y2=2.815
r116 13 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r117 13 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.815
r118 4 26 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=5.71
+ $Y=1.96 $X2=5.91 $Y2=2.815
r119 4 23 400 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=1 $X=5.71
+ $Y=1.96 $X2=5.91 $Y2=2.115
r120 3 65 600 $w=1.7e-07 $l=4.20595e-07 $layer=licon1_PDIFF $count=1 $X=4.45
+ $Y=2.54 $X2=4.755 $Y2=2.815
r121 2 19 600 $w=1.7e-07 $l=9.74192e-07 $layer=licon1_PDIFF $count=1 $X=2.26
+ $Y=1.96 $X2=2.515 $Y2=2.815
r122 1 15 600 $w=1.7e-07 $l=7.88686e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.12 $X2=0.78 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_1%Q 1 2 9 14 15 16
c23 16 0 1.77844e-19 $X=6.48 $Y=0.555
r24 22 23 9.7361 $w=5.33e-07 $l=1.65e-07 $layer=LI1_cond $X=6.367 $Y=0.675
+ $X2=6.367 $Y2=0.84
r25 16 22 2.68279 $w=5.33e-07 $l=1.2e-07 $layer=LI1_cond $X=6.367 $Y=0.555
+ $X2=6.367 $Y2=0.675
r26 15 23 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=6.55 $Y=1.82
+ $X2=6.55 $Y2=0.84
r27 14 15 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.455 $Y=1.985
+ $X2=6.455 $Y2=1.82
r28 7 14 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=6.455 $Y=2 $X2=6.455
+ $Y2=1.985
r29 7 9 26.09 $w=3.58e-07 $l=8.15e-07 $layer=LI1_cond $X=6.455 $Y=2 $X2=6.455
+ $Y2=2.815
r30 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.84 $X2=6.44 $Y2=1.985
r31 2 9 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.84 $X2=6.44 $Y2=2.815
r32 1 22 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=6.125
+ $Y=0.37 $X2=6.265 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LS__DLRTP_1%VGND 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 38 44 62 63 66
r74 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r75 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r76 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r77 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r78 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r79 56 59 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r80 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r81 54 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r82 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r83 51 66 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.68 $Y=0 $X2=2.487
+ $Y2=0
r84 51 53 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.68 $Y=0 $X2=4.08
+ $Y2=0
r85 50 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r86 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r87 47 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r88 46 49 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r89 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r90 44 66 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.487
+ $Y2=0
r91 44 49 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.16
+ $Y2=0
r92 42 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r93 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r94 38 54 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r95 38 67 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=2.64
+ $Y2=0
r96 36 59 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.52
+ $Y2=0
r97 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.755
+ $Y2=0
r98 35 62 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.92 $Y=0 $X2=6.48
+ $Y2=0
r99 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.92 $Y=0 $X2=5.755
+ $Y2=0
r100 33 53 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.08
+ $Y2=0
r101 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.375
+ $Y2=0
r102 32 56 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=4.54 $Y=0 $X2=4.56
+ $Y2=0
r103 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.54 $Y=0 $X2=4.375
+ $Y2=0
r104 30 41 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=0
+ $X2=0.72 $Y2=0
r105 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.885 $Y=0 $X2=0.97
+ $Y2=0
r106 29 46 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.2
+ $Y2=0
r107 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=0 $X2=0.97
+ $Y2=0
r108 25 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.755 $Y=0.085
+ $X2=5.755 $Y2=0
r109 25 27 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=5.755 $Y=0.085
+ $X2=5.755 $Y2=0.675
r110 21 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.375 $Y=0.085
+ $X2=4.375 $Y2=0
r111 21 23 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.375 $Y=0.085
+ $X2=4.375 $Y2=0.58
r112 17 66 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.487 $Y=0.085
+ $X2=2.487 $Y2=0
r113 17 19 12.8714 $w=3.83e-07 $l=4.3e-07 $layer=LI1_cond $X=2.487 $Y=0.085
+ $X2=2.487 $Y2=0.515
r114 13 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.97 $Y=0.085
+ $X2=0.97 $Y2=0
r115 13 15 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=0.97 $Y=0.085
+ $X2=0.97 $Y2=0.515
r116 4 27 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=5.615
+ $Y=0.37 $X2=5.755 $Y2=0.675
r117 3 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.235
+ $Y=0.37 $X2=4.375 $Y2=0.58
r118 2 19 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=2.315
+ $Y=0.37 $X2=2.485 $Y2=0.515
r119 1 15 91 $w=1.7e-07 $l=3.16702e-07 $layer=licon1_NDIFF $count=2 $X=0.675
+ $Y=0.56 $X2=0.97 $Y2=0.515
.ends

