* File: sky130_fd_sc_ls__clkinv_1.pex.spice
* Created: Fri Aug 28 13:10:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__CLKINV_1%A 1 3 6 8 10 11 12 18 21 25
r34 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.765 $X2=0.59 $Y2=1.765
r35 21 23 50.3829 $w=6.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.72 $Y=1.085
+ $X2=0.72 $Y2=0.92
r36 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.085 $X2=0.59 $Y2=1.085
r37 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.425 $X2=0.59 $Y2=1.425
r38 16 25 12.2422 $w=6.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.72 $Y=1.615
+ $X2=0.72 $Y2=1.765
r39 16 18 16.1358 $w=6.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.72 $Y=1.615
+ $X2=0.72 $Y2=1.425
r40 15 21 12.7388 $w=6.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.72 $Y=1.235
+ $X2=0.72 $Y2=1.085
r41 15 18 16.1358 $w=6.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.72 $Y=1.235
+ $X2=0.72 $Y2=1.425
r42 12 26 2.40157 $w=5.08e-07 $l=1e-07 $layer=LI1_cond $X=0.44 $Y=1.665 $X2=0.44
+ $Y2=1.765
r43 12 19 5.76378 $w=5.08e-07 $l=2.4e-07 $layer=LI1_cond $X=0.44 $Y=1.665
+ $X2=0.44 $Y2=1.425
r44 11 19 3.12205 $w=5.08e-07 $l=1.3e-07 $layer=LI1_cond $X=0.44 $Y=1.295
+ $X2=0.44 $Y2=1.425
r45 11 22 5.04331 $w=5.08e-07 $l=2.1e-07 $layer=LI1_cond $X=0.44 $Y=1.295
+ $X2=0.44 $Y2=1.085
r46 8 25 50.8109 $w=2.78e-07 $l=3.76032e-07 $layer=POLY_cond $X=0.945 $Y=2.045
+ $X2=0.72 $Y2=1.765
r47 8 10 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.945 $Y=2.045
+ $X2=0.945 $Y2=2.54
r48 6 23 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.565 $Y=0.58
+ $X2=0.565 $Y2=0.92
r49 1 25 50.8109 $w=2.78e-07 $l=3.76032e-07 $layer=POLY_cond $X=0.495 $Y=2.045
+ $X2=0.72 $Y2=1.765
r50 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=2.045
+ $X2=0.495 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_1%VPWR 1 2 7 9 11 13 15 17 27
r21 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r22 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r23 18 23 4.02368 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.177 $Y2=3.33
r24 18 20 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.72 $Y2=3.33
r25 17 26 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.222 $Y2=3.33
r26 17 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r28 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r29 15 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 11 26 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.222 $Y2=3.33
r31 11 13 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.79
r32 7 23 3.11948 $w=2.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.177 $Y2=3.33
r33 7 9 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=0.23 $Y=3.245 $X2=0.23
+ $Y2=2.265
r34 2 13 600 $w=1.7e-07 $l=7.41215e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=2.12 $X2=1.17 $Y2=2.79
r35 1 9 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.27 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_1%Y 1 2 9 11 15 16 17 18 19 26 36 45
r28 40 43 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.695 $Y=2.265
+ $X2=0.72 $Y2=2.265
r29 27 45 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=1.205 $Y=2.1
+ $X2=1.205 $Y2=2.265
r30 27 36 3.1212 $w=2.38e-07 $l=6.5e-08 $layer=LI1_cond $X=1.205 $Y=2.1
+ $X2=1.205 $Y2=2.035
r31 19 45 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.2 $Y=2.265
+ $X2=1.205 $Y2=2.265
r32 19 43 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=2.265
+ $X2=0.72 $Y2=2.265
r33 19 36 0.480185 $w=2.38e-07 $l=1e-08 $layer=LI1_cond $X=1.205 $Y=2.025
+ $X2=1.205 $Y2=2.035
r34 18 19 17.2866 $w=2.38e-07 $l=3.6e-07 $layer=LI1_cond $X=1.205 $Y=1.665
+ $X2=1.205 $Y2=2.025
r35 17 18 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.205 $Y=1.295
+ $X2=1.205 $Y2=1.665
r36 16 17 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.205 $Y=0.925
+ $X2=1.205 $Y2=1.295
r37 16 26 11.7645 $w=2.38e-07 $l=2.45e-07 $layer=LI1_cond $X=1.205 $Y=0.925
+ $X2=1.205 $Y2=0.68
r38 15 26 4.07572 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=1.205 $Y=0.515
+ $X2=1.205 $Y2=0.68
r39 11 15 2.96416 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=1.085 $Y=0.515
+ $X2=1.205 $Y2=0.515
r40 11 13 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.085 $Y=0.515
+ $X2=0.78 $Y2=0.515
r41 7 40 1.70047 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.695 $Y=2.43
+ $X2=0.695 $Y2=2.265
r42 7 9 14.8171 $w=2.78e-07 $l=3.6e-07 $layer=LI1_cond $X=0.695 $Y=2.43
+ $X2=0.695 $Y2=2.79
r43 2 43 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=2.12 $X2=0.72 $Y2=2.265
r44 2 9 600 $w=1.7e-07 $l=7.41215e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=2.12 $X2=0.72 $Y2=2.79
r45 1 15 182 $w=1.7e-07 $l=5.88048e-07 $layer=licon1_NDIFF $count=1 $X=0.64
+ $Y=0.37 $X2=1.16 $Y2=0.515
r46 1 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__CLKINV_1%VGND 1 4 6 8 12 13
r14 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r15 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r16 10 16 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r17 10 12 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=1.2
+ $Y2=0
r18 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r19 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r20 4 16 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r21 4 6 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.55
r22 1 6 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.55
.ends

