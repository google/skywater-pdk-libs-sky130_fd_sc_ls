* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ls__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
M1000 VGND a_1598_93# a_1550_119# VNB nshort w=420000u l=150000u
+  ad=1.4689e+12p pd=1.212e+07u as=1.008e+11p ps=1.32e+06u
M1001 a_1598_93# a_1266_119# a_1736_119# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1002 a_1266_119# a_507_347# a_841_288# VPB phighvt w=1e+06u l=150000u
+  ad=4.477e+11p pd=3.4e+06u as=7.8e+11p ps=3.56e+06u
M1003 VPWR a_1598_93# a_1547_508# VPB phighvt w=420000u l=150000u
+  ad=1.83395e+12p pd=1.721e+07u as=1.134e+11p ps=1.38e+06u
M1004 Q a_1934_94# VPWR VPB phighvt w=1.12e+06u l=150000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1005 a_507_347# a_300_74# VGND VNB nshort w=740000u l=150000u
+  ad=2.479e+11p pd=2.15e+06u as=0p ps=0u
M1006 a_1266_119# a_300_74# a_841_288# VNB nshort w=740000u l=150000u
+  ad=6.134e+11p pd=4.02e+06u as=2.146e+11p ps=2.06e+06u
M1007 a_300_74# CLK_N VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.9e+11p pd=2.58e+06u as=0p ps=0u
M1008 a_841_288# a_714_127# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_714_127# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.478e+11p pd=2.86e+06u as=0p ps=0u
M1010 a_1736_119# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_714_127# a_300_74# a_33_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.499e+11p ps=2.87e+06u
M1012 a_1547_508# a_300_74# a_1266_119# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_714_127# a_507_347# a_33_74# VNB nshort w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=2.31e+11p ps=2.78e+06u
M1014 VPWR a_1266_119# a_1598_93# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1015 VPWR a_1266_119# a_1934_94# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.31e+11p ps=2.23e+06u
M1016 VGND RESET_B a_922_127# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1017 a_507_347# a_300_74# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=4.0345e+11p pd=2.86e+06u as=0p ps=0u
M1018 a_817_463# a_507_347# a_714_127# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1019 a_1598_93# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_841_288# a_714_127# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_1266_119# a_1934_94# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1022 a_1550_119# a_507_347# a_1266_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_33_74# D VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR RESET_B a_33_74# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND RESET_B a_120_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1026 a_922_127# a_841_288# a_850_127# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1027 a_300_74# CLK_N VGND VNB nshort w=740000u l=150000u
+  ad=2.035e+11p pd=2.03e+06u as=0p ps=0u
M1028 Q a_1934_94# VGND VNB nshort w=740000u l=150000u
+  ad=2.146e+11p pd=2.06e+06u as=0p ps=0u
M1029 a_120_74# D a_33_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_850_127# a_300_74# a_714_127# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_841_288# a_817_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
