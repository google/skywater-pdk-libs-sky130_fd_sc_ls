* File: sky130_fd_sc_ls__o22a_4.pex.spice
* Created: Wed Sep  2 11:20:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__O22A_4%A2 1 3 6 8 10 11 13 14 20 21
r57 21 22 3.70769 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=1.425 $Y=1.64
+ $X2=1.455 $Y2=1.64
r58 19 21 9.26923 $w=3.9e-07 $l=7.5e-08 $layer=POLY_cond $X=1.35 $Y=1.64
+ $X2=1.425 $Y2=1.64
r59 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.35
+ $Y=1.615 $X2=1.35 $Y2=1.615
r60 14 20 0.892596 $w=6.68e-07 $l=5e-08 $layer=LI1_cond $X=1.18 $Y=1.665
+ $X2=1.18 $Y2=1.615
r61 11 22 25.2441 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.455 $Y=1.885
+ $X2=1.455 $Y2=1.64
r62 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.885
+ $X2=1.455 $Y2=2.46
r63 8 21 25.2441 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.425 $Y=1.395
+ $X2=1.425 $Y2=1.64
r64 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.425 $Y=1.395
+ $X2=1.425 $Y2=1
r65 4 19 43.8744 $w=3.9e-07 $l=3.55e-07 $layer=POLY_cond $X=0.995 $Y=1.64
+ $X2=1.35 $Y2=1.64
r66 4 16 4.94359 $w=3.9e-07 $l=4e-08 $layer=POLY_cond $X=0.995 $Y=1.64 $X2=0.955
+ $Y2=1.64
r67 4 6 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.995 $Y=1.45
+ $X2=0.995 $Y2=1
r68 1 16 25.2441 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=0.955 $Y=1.885
+ $X2=0.955 $Y2=1.64
r69 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.955 $Y=1.885
+ $X2=0.955 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_4%A1 2 4 6 7 9 10 11 12 14 18 19
r67 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.01
+ $Y=1.615 $X2=2.01 $Y2=1.615
r68 19 23 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.16 $Y=1.615
+ $X2=2.01 $Y2=1.615
r69 16 22 38.5916 $w=2.93e-07 $l=1.86145e-07 $layer=POLY_cond $X=1.965 $Y=1.45
+ $X2=2.01 $Y2=1.615
r70 16 18 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.965 $Y=1.45
+ $X2=1.965 $Y2=1
r71 15 18 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.965 $Y=0.31
+ $X2=1.965 $Y2=1
r72 12 22 55.8646 $w=2.93e-07 $l=2.96226e-07 $layer=POLY_cond $X=1.955 $Y=1.885
+ $X2=2.01 $Y2=1.615
r73 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.885
+ $X2=1.955 $Y2=2.46
r74 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.89 $Y=0.235
+ $X2=1.965 $Y2=0.31
r75 10 11 676.851 $w=1.5e-07 $l=1.32e-06 $layer=POLY_cond $X=1.89 $Y=0.235
+ $X2=0.57 $Y2=0.235
r76 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.46
r77 4 6 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.395
+ $X2=0.495 $Y2=1
r78 3 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.495 $Y=0.31
+ $X2=0.57 $Y2=0.235
r79 3 6 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=0.31
+ $X2=0.495 $Y2=1
r80 2 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.795 $X2=0.505
+ $Y2=1.885
r81 1 4 70.5366 $w=1.64e-07 $l=2.44949e-07 $layer=POLY_cond $X=0.505 $Y=1.635
+ $X2=0.495 $Y2=1.395
r82 1 2 62.1936 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=0.505 $Y=1.635
+ $X2=0.505 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_4%B2 3 5 7 8 10 11 13 14 15 22 23
c59 22 0 1.52901e-19 $X=3.34 $Y=1.615
c60 3 0 1.28833e-19 $X=2.925 $Y=1
r61 23 24 3.03526 $w=3.97e-07 $l=2.5e-08 $layer=POLY_cond $X=3.43 $Y=1.64
+ $X2=3.455 $Y2=1.64
r62 21 23 10.927 $w=3.97e-07 $l=9e-08 $layer=POLY_cond $X=3.34 $Y=1.64 $X2=3.43
+ $Y2=1.64
r63 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.34
+ $Y=1.615 $X2=3.34 $Y2=1.615
r64 19 21 46.7431 $w=3.97e-07 $l=3.85e-07 $layer=POLY_cond $X=2.955 $Y=1.64
+ $X2=3.34 $Y2=1.64
r65 15 22 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=3.12 $Y=1.615
+ $X2=3.34 $Y2=1.615
r66 14 15 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.615
+ $X2=3.12 $Y2=1.615
r67 11 24 25.678 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=3.455 $Y=1.885
+ $X2=3.455 $Y2=1.64
r68 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.455 $Y=1.885
+ $X2=3.455 $Y2=2.46
r69 8 23 25.678 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=3.43 $Y=1.395
+ $X2=3.43 $Y2=1.64
r70 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.43 $Y=1.395
+ $X2=3.43 $Y2=1
r71 5 19 25.678 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=2.955 $Y=1.885
+ $X2=2.955 $Y2=1.64
r72 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.955 $Y=1.885
+ $X2=2.955 $Y2=2.46
r73 1 19 3.64232 $w=3.97e-07 $l=3e-08 $layer=POLY_cond $X=2.925 $Y=1.64
+ $X2=2.955 $Y2=1.64
r74 1 3 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.925 $Y=1.45
+ $X2=2.925 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_4%B1 4 5 6 7 9 10 15 17 18 20 23 24 26
c81 24 0 1.28833e-19 $X=2.16 $Y=0.555
c82 17 0 1.52901e-19 $X=3.955 $Y=1.795
r83 29 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.445 $Y=0.405
+ $X2=2.445 $Y2=0.57
r84 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.445
+ $Y=0.405 $X2=2.445 $Y2=0.405
r85 26 29 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.445 $Y=0.235
+ $X2=2.445 $Y2=0.405
r86 24 30 9.79437 $w=3.55e-07 $l=2.85e-07 $layer=LI1_cond $X=2.16 $Y=0.462
+ $X2=2.445 $Y2=0.462
r87 22 23 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.915 $Y=1.395
+ $X2=3.915 $Y2=1.545
r88 18 20 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.955 $Y=1.885
+ $X2=3.955 $Y2=2.46
r89 17 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.955 $Y=1.795
+ $X2=3.955 $Y2=1.885
r90 17 23 97.1774 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=3.955 $Y=1.795
+ $X2=3.955 $Y2=1.545
r91 15 22 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.86 $Y=1 $X2=3.86
+ $Y2=1.395
r92 12 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.86 $Y=0.31
+ $X2=3.86 $Y2=1
r93 11 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.61 $Y=0.235
+ $X2=2.445 $Y2=0.235
r94 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.785 $Y=0.235
+ $X2=3.86 $Y2=0.31
r95 10 11 602.5 $w=1.5e-07 $l=1.175e-06 $layer=POLY_cond $X=3.785 $Y=0.235
+ $X2=2.61 $Y2=0.235
r96 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.505 $Y=1.885
+ $X2=2.505 $Y2=2.46
r97 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.505 $Y=1.795 $X2=2.505
+ $Y2=1.885
r98 5 21 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.505 $Y=1.485
+ $X2=2.505 $Y2=1.395
r99 5 6 120.5 $w=1.8e-07 $l=3.1e-07 $layer=POLY_cond $X=2.505 $Y=1.485 $X2=2.505
+ $Y2=1.795
r100 4 21 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.49 $Y=1 $X2=2.49
+ $Y2=1.395
r101 4 31 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.49 $Y=1 $X2=2.49
+ $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_4%A_206_392# 1 2 3 4 13 15 18 20 22 25 27 29 32
+ 34 36 39 43 51 54 55 57 58 60 63 67 69 72 73 75 85
c176 58 0 1.20589e-19 $X=3.845 $Y=1.595
r177 85 86 7.40503 $w=3.58e-07 $l=5.5e-08 $layer=POLY_cond $X=6.165 $Y=1.557
+ $X2=6.22 $Y2=1.557
r178 84 85 50.4888 $w=3.58e-07 $l=3.75e-07 $layer=POLY_cond $X=5.79 $Y=1.557
+ $X2=6.165 $Y2=1.557
r179 83 84 10.0978 $w=3.58e-07 $l=7.5e-08 $layer=POLY_cond $X=5.715 $Y=1.557
+ $X2=5.79 $Y2=1.557
r180 80 81 49.8156 $w=3.58e-07 $l=3.7e-07 $layer=POLY_cond $X=4.99 $Y=1.557
+ $X2=5.36 $Y2=1.557
r181 79 80 8.07821 $w=3.58e-07 $l=6e-08 $layer=POLY_cond $X=4.93 $Y=1.557
+ $X2=4.99 $Y2=1.557
r182 76 79 47.1229 $w=3.58e-07 $l=3.5e-07 $layer=POLY_cond $X=4.58 $Y=1.557
+ $X2=4.93 $Y2=1.557
r183 76 77 10.0978 $w=3.58e-07 $l=7.5e-08 $layer=POLY_cond $X=4.58 $Y=1.557
+ $X2=4.505 $Y2=1.557
r184 75 76 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.58
+ $Y=1.515 $X2=4.58 $Y2=1.515
r185 71 73 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=0.79
+ $X2=3.81 $Y2=0.79
r186 71 72 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=0.79
+ $X2=3.48 $Y2=0.79
r187 64 83 15.4832 $w=3.58e-07 $l=1.15e-07 $layer=POLY_cond $X=5.6 $Y=1.557
+ $X2=5.715 $Y2=1.557
r188 64 81 32.3129 $w=3.58e-07 $l=2.4e-07 $layer=POLY_cond $X=5.6 $Y=1.557
+ $X2=5.36 $Y2=1.557
r189 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.6
+ $Y=1.515 $X2=5.6 $Y2=1.515
r190 61 75 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.585 $Y=1.515
+ $X2=4.5 $Y2=1.515
r191 61 63 35.4464 $w=3.28e-07 $l=1.015e-06 $layer=LI1_cond $X=4.585 $Y=1.515
+ $X2=5.6 $Y2=1.515
r192 60 75 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.5 $Y=1.35 $X2=4.5
+ $Y2=1.515
r193 59 60 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.5 $Y=0.92 $X2=4.5
+ $Y2=1.35
r194 57 75 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.415 $Y=1.595
+ $X2=4.5 $Y2=1.515
r195 57 58 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.415 $Y=1.595
+ $X2=3.845 $Y2=1.595
r196 55 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.415 $Y=0.835
+ $X2=4.5 $Y2=0.92
r197 55 73 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.415 $Y=0.835
+ $X2=3.81 $Y2=0.835
r198 53 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.76 $Y=1.68
+ $X2=3.845 $Y2=1.595
r199 53 54 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.76 $Y=1.68
+ $X2=3.76 $Y2=1.95
r200 52 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.395 $Y=2.035
+ $X2=3.23 $Y2=2.035
r201 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.675 $Y=2.035
+ $X2=3.76 $Y2=1.95
r202 51 52 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.675 $Y=2.035
+ $X2=3.395 $Y2=2.035
r203 47 72 47.4444 $w=1.78e-07 $l=7.7e-07 $layer=LI1_cond $X=2.71 $Y=0.83
+ $X2=3.48 $Y2=0.83
r204 44 67 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=2.035
+ $X2=1.23 $Y2=2.035
r205 43 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.065 $Y=2.035
+ $X2=3.23 $Y2=2.035
r206 43 44 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=3.065 $Y=2.035
+ $X2=1.395 $Y2=2.035
r207 37 86 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.22 $Y=1.35
+ $X2=6.22 $Y2=1.557
r208 37 39 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.22 $Y=1.35
+ $X2=6.22 $Y2=0.74
r209 34 85 23.1716 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.165 $Y=1.765
+ $X2=6.165 $Y2=1.557
r210 34 36 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.165 $Y=1.765
+ $X2=6.165 $Y2=2.4
r211 30 84 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.79 $Y=1.35
+ $X2=5.79 $Y2=1.557
r212 30 32 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.79 $Y=1.35
+ $X2=5.79 $Y2=0.74
r213 27 83 23.1716 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.715 $Y=1.765
+ $X2=5.715 $Y2=1.557
r214 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.715 $Y=1.765
+ $X2=5.715 $Y2=2.4
r215 23 81 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.36 $Y=1.35
+ $X2=5.36 $Y2=1.557
r216 23 25 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.36 $Y=1.35
+ $X2=5.36 $Y2=0.74
r217 20 80 23.1716 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.99 $Y=1.765
+ $X2=4.99 $Y2=1.557
r218 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.99 $Y=1.765
+ $X2=4.99 $Y2=2.4
r219 16 79 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.93 $Y=1.35
+ $X2=4.93 $Y2=1.557
r220 16 18 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.93 $Y=1.35
+ $X2=4.93 $Y2=0.74
r221 13 77 23.1716 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.505 $Y=1.765
+ $X2=4.505 $Y2=1.557
r222 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.505 $Y=1.765
+ $X2=4.505 $Y2=2.4
r223 4 69 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=3.03
+ $Y=1.96 $X2=3.23 $Y2=2.115
r224 3 67 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.96 $X2=1.23 $Y2=2.115
r225 2 71 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.68 $X2=3.645 $Y2=0.83
r226 1 47 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=2.565
+ $Y=0.68 $X2=2.71 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_4%VPWR 1 2 3 4 5 16 18 24 28 34 36 38 43 44 46
+ 47 48 50 68 76 80
r81 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r82 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r83 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r84 71 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r85 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r86 68 79 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6.497 $Y2=3.33
r87 68 70 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.275 $Y=3.33 $X2=6
+ $Y2=3.33
r88 67 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r89 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r90 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r91 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r92 61 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r93 60 63 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r94 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r95 58 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.23 $Y2=3.33
r96 58 60 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.64 $Y2=3.33
r97 57 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r98 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r99 54 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 54 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r101 53 56 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r102 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 51 73 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r104 51 53 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r105 50 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=2.23 $Y2=3.33
r106 50 56 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=1.68 $Y2=3.33
r107 48 64 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r108 48 61 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=2.64 $Y2=3.33
r109 46 66 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.2 $Y=3.33
+ $X2=5.04 $Y2=3.33
r110 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.2 $Y=3.33
+ $X2=5.365 $Y2=3.33
r111 45 70 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=5.53 $Y=3.33 $X2=6
+ $Y2=3.33
r112 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.53 $Y=3.33
+ $X2=5.365 $Y2=3.33
r113 43 63 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=4.1 $Y=3.33 $X2=4.08
+ $Y2=3.33
r114 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.1 $Y=3.33
+ $X2=4.265 $Y2=3.33
r115 42 66 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=5.04 $Y2=3.33
r116 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.265 $Y2=3.33
r117 38 41 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.44 $Y=1.985
+ $X2=6.44 $Y2=2.815
r118 36 79 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.497 $Y2=3.33
r119 36 41 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.44 $Y2=2.815
r120 32 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.365 $Y=3.245
+ $X2=5.365 $Y2=3.33
r121 32 34 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=5.365 $Y=3.245
+ $X2=5.365 $Y2=2.355
r122 28 31 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=4.265 $Y=2.015
+ $X2=4.265 $Y2=2.415
r123 26 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.265 $Y=3.245
+ $X2=4.265 $Y2=3.33
r124 26 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.265 $Y=3.245
+ $X2=4.265 $Y2=2.415
r125 22 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=3.33
r126 22 24 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=2.455
r127 18 21 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.24 $Y=2.105
+ $X2=0.24 $Y2=2.815
r128 16 73 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r129 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r130 5 41 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=1.84 $X2=6.44 $Y2=2.815
r131 5 38 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=1.84 $X2=6.44 $Y2=1.985
r132 4 34 300 $w=1.7e-07 $l=6.47862e-07 $layer=licon1_PDIFF $count=2 $X=5.065
+ $Y=1.84 $X2=5.365 $Y2=2.355
r133 3 31 300 $w=1.7e-07 $l=5.60312e-07 $layer=licon1_PDIFF $count=2 $X=4.03
+ $Y=1.96 $X2=4.265 $Y2=2.415
r134 3 28 600 $w=1.7e-07 $l=2.61056e-07 $layer=licon1_PDIFF $count=1 $X=4.03
+ $Y=1.96 $X2=4.265 $Y2=2.015
r135 2 24 300 $w=1.7e-07 $l=5.86536e-07 $layer=licon1_PDIFF $count=2 $X=2.03
+ $Y=1.96 $X2=2.23 $Y2=2.455
r136 1 21 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r137 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_4%A_116_392# 1 2 9 13 14 17
r27 15 17 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.73 $Y=2.905
+ $X2=1.73 $Y2=2.455
r28 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.565 $Y=2.99
+ $X2=1.73 $Y2=2.905
r29 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=2.99
+ $X2=0.895 $Y2=2.99
r30 9 12 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.73 $Y=2.115 $X2=0.73
+ $Y2=2.815
r31 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.73 $Y=2.905
+ $X2=0.895 $Y2=2.99
r32 7 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.73 $Y=2.905 $X2=0.73
+ $Y2=2.815
r33 2 17 300 $w=1.7e-07 $l=5.86536e-07 $layer=licon1_PDIFF $count=2 $X=1.53
+ $Y=1.96 $X2=1.73 $Y2=2.455
r34 1 12 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.96 $X2=0.73 $Y2=2.815
r35 1 9 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.96 $X2=0.73 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_4%A_516_392# 1 2 9 11 12 15
r25 13 15 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.73 $Y=2.905
+ $X2=3.73 $Y2=2.455
r26 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.565 $Y=2.99
+ $X2=3.73 $Y2=2.905
r27 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.565 $Y=2.99
+ $X2=2.895 $Y2=2.99
r28 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.73 $Y=2.905
+ $X2=2.895 $Y2=2.99
r29 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.73 $Y=2.905 $X2=2.73
+ $Y2=2.455
r30 2 15 300 $w=1.7e-07 $l=5.86536e-07 $layer=licon1_PDIFF $count=2 $X=3.53
+ $Y=1.96 $X2=3.73 $Y2=2.455
r31 1 9 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=2.58
+ $Y=1.96 $X2=2.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_4%X 1 2 3 4 13 15 17 21 23 24 27 31 33 34 38 42
r70 41 42 18.7898 $w=2.28e-07 $l=3.75e-07 $layer=LI1_cond $X=6.105 $Y=1.295
+ $X2=6.48 $Y2=1.295
r71 39 41 13.8636 $w=1.76e-07 $l=2e-07 $layer=LI1_cond $X=6.012 $Y=1.095
+ $X2=6.012 $Y2=1.295
r72 34 38 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=6.02 $Y=1.85
+ $X2=5.94 $Y2=1.935
r73 33 41 7.97159 $w=1.76e-07 $l=1.18933e-07 $layer=LI1_cond $X=6.02 $Y=1.41
+ $X2=6.012 $Y2=1.295
r74 33 34 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=6.02 $Y=1.41
+ $X2=6.02 $Y2=1.85
r75 29 39 5.6459 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=6.012 $Y=1.01
+ $X2=6.012 $Y2=1.095
r76 29 31 29.6757 $w=1.83e-07 $l=4.95e-07 $layer=LI1_cond $X=6.012 $Y=1.01
+ $X2=6.012 $Y2=0.515
r77 25 38 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=2.02 $X2=5.94
+ $Y2=1.935
r78 25 27 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=5.94 $Y=2.02
+ $X2=5.94 $Y2=2.815
r79 23 39 0.927112 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=5.92 $Y=1.095
+ $X2=6.012 $Y2=1.095
r80 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.92 $Y=1.095
+ $X2=5.23 $Y2=1.095
r81 19 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.105 $Y=1.01
+ $X2=5.23 $Y2=1.095
r82 19 21 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=5.105 $Y=1.01
+ $X2=5.105 $Y2=0.515
r83 18 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.93 $Y=1.935
+ $X2=4.765 $Y2=1.935
r84 17 38 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.775 $Y=1.935
+ $X2=5.94 $Y2=1.935
r85 17 18 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=5.775 $Y=1.935
+ $X2=4.93 $Y2=1.935
r86 13 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.765 $Y=2.02
+ $X2=4.765 $Y2=1.935
r87 13 15 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=4.765 $Y=2.02
+ $X2=4.765 $Y2=2.815
r88 4 38 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.84 $X2=5.94 $Y2=2.015
r89 4 27 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.84 $X2=5.94 $Y2=2.815
r90 3 36 400 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_PDIFF $count=1 $X=4.58
+ $Y=1.84 $X2=4.765 $Y2=2.015
r91 3 15 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=4.58
+ $Y=1.84 $X2=4.765 $Y2=2.815
r92 2 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.865
+ $Y=0.37 $X2=6.005 $Y2=0.515
r93 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.005
+ $Y=0.37 $X2=5.145 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_4%A_27_136# 1 2 3 4 5 18 20 21 24 32 35 36 38
+ 39
r62 38 39 8.29777 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=1.215
+ $X2=3.91 $Y2=1.215
r63 34 36 8.11354 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=1.06
+ $X2=2.375 $Y2=1.06
r64 34 35 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=1.06
+ $X2=2.045 $Y2=1.06
r65 31 39 42.9043 $w=1.88e-07 $l=7.35e-07 $layer=LI1_cond $X=3.175 $Y=1.185
+ $X2=3.91 $Y2=1.185
r66 31 36 46.6986 $w=1.88e-07 $l=8e-07 $layer=LI1_cond $X=3.175 $Y=1.185
+ $X2=2.375 $Y2=1.185
r67 27 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.375 $Y=1.195
+ $X2=1.25 $Y2=1.195
r68 27 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.375 $Y=1.195
+ $X2=2.045 $Y2=1.195
r69 22 32 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=1.11
+ $X2=1.25 $Y2=1.195
r70 22 24 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=1.25 $Y=1.11
+ $X2=1.25 $Y2=0.97
r71 20 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.125 $Y=1.195
+ $X2=1.25 $Y2=1.195
r72 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.125 $Y=1.195
+ $X2=0.445 $Y2=1.195
r73 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.11
+ $X2=0.445 $Y2=1.195
r74 16 18 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.28 $Y=1.11
+ $X2=0.28 $Y2=0.825
r75 5 38 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=3.935
+ $Y=0.68 $X2=4.075 $Y2=1.175
r76 4 31 182 $w=1.7e-07 $l=5.75891e-07 $layer=licon1_NDIFF $count=1 $X=3 $Y=0.68
+ $X2=3.175 $Y2=1.175
r77 3 34 182 $w=1.7e-07 $l=4.57165e-07 $layer=licon1_NDIFF $count=1 $X=2.04
+ $Y=0.68 $X2=2.21 $Y2=1.06
r78 2 24 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.68 $X2=1.21 $Y2=0.97
r79 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.68 $X2=0.28 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LS__O22A_4%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43 48
+ 56 61 67 70 73 76 80
r86 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r87 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r88 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r89 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r90 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r91 65 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r92 65 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r93 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r94 62 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.74 $Y=0 $X2=5.575
+ $Y2=0
r95 62 64 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.74 $Y=0 $X2=6
+ $Y2=0
r96 61 79 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.275 $Y=0 $X2=6.497
+ $Y2=0
r97 61 64 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.275 $Y=0 $X2=6
+ $Y2=0
r98 60 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r99 60 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r100 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r101 57 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.8 $Y=0 $X2=4.635
+ $Y2=0
r102 57 59 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.8 $Y=0 $X2=5.04
+ $Y2=0
r103 56 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.41 $Y=0 $X2=5.575
+ $Y2=0
r104 56 59 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.41 $Y=0 $X2=5.04
+ $Y2=0
r105 55 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r106 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r107 52 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r108 51 54 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r109 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r110 49 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.71
+ $Y2=0
r111 49 51 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=2.16 $Y2=0
r112 48 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.47 $Y=0 $X2=4.635
+ $Y2=0
r113 48 54 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.47 $Y=0 $X2=4.08
+ $Y2=0
r114 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r115 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r116 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r118 44 46 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r119 43 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.71
+ $Y2=0
r120 43 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.2
+ $Y2=0
r121 41 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r122 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r123 38 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r124 38 40 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r125 36 55 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r126 36 52 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=2.16
+ $Y2=0
r127 32 79 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.497 $Y2=0
r128 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.44 $Y2=0.515
r129 28 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.575 $Y=0.085
+ $X2=5.575 $Y2=0
r130 28 30 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=5.575 $Y=0.085
+ $X2=5.575 $Y2=0.625
r131 24 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.635 $Y=0.085
+ $X2=4.635 $Y2=0
r132 24 26 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=4.635 $Y=0.085
+ $X2=4.635 $Y2=0.415
r133 20 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r134 20 22 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.84
r135 16 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r136 16 18 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.84
r137 5 34 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=6.295
+ $Y=0.37 $X2=6.44 $Y2=0.515
r138 4 30 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=5.435
+ $Y=0.37 $X2=5.575 $Y2=0.625
r139 3 26 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.49
+ $Y=0.27 $X2=4.635 $Y2=0.415
r140 2 22 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.68 $X2=1.71 $Y2=0.84
r141 1 18 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.68 $X2=0.78 $Y2=0.84
.ends

