* File: sky130_fd_sc_ls__or2_1.pex.spice
* Created: Wed Sep  2 11:24:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LS__OR2_1%B 1 3 5 8 9 12 14
c27 3 0 8.55747e-20 $X=0.685 $Y=1.765
r28 9 14 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.61 $Y2=1.365
r29 8 12 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.7 $Y=0.835 $X2=0.7
+ $Y2=1.22
r30 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.685 $Y=1.765
+ $X2=0.685 $Y2=2.26
r31 1 3 149.859 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=0.685 $Y=1.385
+ $X2=0.685 $Y2=1.765
r32 1 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.385 $X2=0.61 $Y2=1.385
r33 1 12 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.685 $Y=1.385
+ $X2=0.685 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_1%A 1 3 6 8 12
c36 12 0 8.55747e-20 $X=1.21 $Y=1.515
c37 6 0 7.78164e-20 $X=1.325 $Y=0.835
c38 1 0 6.83128e-20 $X=1.105 $Y=1.765
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.21
+ $Y=1.515 $X2=1.21 $Y2=1.515
r40 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.21 $Y=1.665
+ $X2=1.21 $Y2=1.515
r41 4 11 38.6002 $w=3.3e-07 $l=2.1609e-07 $layer=POLY_cond $X=1.325 $Y=1.35
+ $X2=1.207 $Y2=1.515
r42 4 6 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.325 $Y=1.35
+ $X2=1.325 $Y2=0.835
r43 1 11 51.0153 $w=3.3e-07 $l=2.96648e-07 $layer=POLY_cond $X=1.105 $Y=1.765
+ $X2=1.207 $Y2=1.515
r44 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.105 $Y=1.765
+ $X2=1.105 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_1%A_63_368# 1 2 7 9 12 16 20 22 23 24 25 27
c67 22 0 6.83128e-20 $X=1.615 $Y=1.095
r68 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.805
+ $Y=1.465 $X2=1.805 $Y2=1.465
r69 24 30 9.13575 $w=2.68e-07 $l=2.05925e-07 $layer=LI1_cond $X=1.7 $Y=1.63
+ $X2=1.792 $Y2=1.465
r70 24 25 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.7 $Y=1.63 $X2=1.7
+ $Y2=1.95
r71 22 30 16.8433 $w=2.68e-07 $l=4.49878e-07 $layer=LI1_cond $X=1.615 $Y=1.095
+ $X2=1.792 $Y2=1.465
r72 22 23 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.615 $Y=1.095
+ $X2=1.24 $Y2=1.095
r73 18 23 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=1.092 $Y=1.01
+ $X2=1.24 $Y2=1.095
r74 18 20 7.42251 $w=2.93e-07 $l=1.9e-07 $layer=LI1_cond $X=1.092 $Y=1.01
+ $X2=1.092 $Y2=0.82
r75 17 27 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=0.625 $Y=2.035
+ $X2=0.46 $Y2=1.97
r76 16 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.615 $Y=2.035
+ $X2=1.7 $Y2=1.95
r77 16 17 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=1.615 $Y=2.035
+ $X2=0.625 $Y2=2.035
r78 10 31 38.5662 $w=2.97e-07 $l=2.06325e-07 $layer=POLY_cond $X=1.905 $Y=1.3
+ $X2=1.812 $Y2=1.465
r79 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.905 $Y=1.3
+ $X2=1.905 $Y2=0.74
r80 7 31 60.4753 $w=2.97e-07 $l=3.38969e-07 $layer=POLY_cond $X=1.895 $Y=1.765
+ $X2=1.812 $Y2=1.465
r81 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.895 $Y=1.765
+ $X2=1.895 $Y2=2.4
r82 2 27 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.315
+ $Y=1.84 $X2=0.46 $Y2=1.985
r83 1 20 182 $w=1.7e-07 $l=4.09878e-07 $layer=licon1_NDIFF $count=1 $X=0.775
+ $Y=0.56 $X2=1.075 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_1%VPWR 1 6 8 10 17 18 21
r24 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r25 18 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r26 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r27 15 21 12.7913 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.475 $Y2=3.33
r28 15 17 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 10 21 12.7913 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=1.165 $Y=3.33
+ $X2=1.475 $Y2=3.33
r31 10 12 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.165 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 8 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=1.68
+ $Y2=3.33
r33 8 13 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=0.24
+ $Y2=3.33
r34 8 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r35 4 21 2.59604 $w=6.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.475 $Y=3.245
+ $X2=1.475 $Y2=3.33
r36 4 6 15.2404 $w=6.18e-07 $l=7.9e-07 $layer=LI1_cond $X=1.475 $Y=3.245
+ $X2=1.475 $Y2=2.455
r37 1 6 200 $w=1.7e-07 $l=8.24363e-07 $layer=licon1_PDIFF $count=3 $X=1.18
+ $Y=1.84 $X2=1.67 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_1%X 1 2 9 13 14 15 16 23 32
c25 13 0 7.78164e-20 $X=2.132 $Y=1.13
r26 21 23 1.2336 $w=3.53e-07 $l=3.8e-08 $layer=LI1_cond $X=2.132 $Y=1.997
+ $X2=2.132 $Y2=2.035
r27 15 16 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=2.132 $Y=2.405
+ $X2=2.132 $Y2=2.775
r28 14 21 0.779116 $w=3.53e-07 $l=2.4e-08 $layer=LI1_cond $X=2.132 $Y=1.973
+ $X2=2.132 $Y2=1.997
r29 14 32 8.1095 $w=3.53e-07 $l=1.53e-07 $layer=LI1_cond $X=2.132 $Y=1.973
+ $X2=2.132 $Y2=1.82
r30 14 15 11.2647 $w=3.53e-07 $l=3.47e-07 $layer=LI1_cond $X=2.132 $Y=2.058
+ $X2=2.132 $Y2=2.405
r31 14 23 0.746653 $w=3.53e-07 $l=2.3e-08 $layer=LI1_cond $X=2.132 $Y=2.058
+ $X2=2.132 $Y2=2.035
r32 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.225 $Y=1.13
+ $X2=2.225 $Y2=1.82
r33 7 13 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=2.132 $Y=0.953
+ $X2=2.132 $Y2=1.13
r34 7 9 14.2189 $w=3.53e-07 $l=4.38e-07 $layer=LI1_cond $X=2.132 $Y=0.953
+ $X2=2.132 $Y2=0.515
r35 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=1.84 $X2=2.12 $Y2=1.985
r36 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=1.84 $X2=2.12 $Y2=2.815
r37 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.98
+ $Y=0.37 $X2=2.12 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LS__OR2_1%VGND 1 2 9 13 16 17 18 23 29 30 33
r32 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r33 30 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r34 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r35 27 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.62
+ $Y2=0
r36 27 29 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=2.16
+ $Y2=0
r37 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.62
+ $Y2=0
r38 23 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.2
+ $Y2=0
r39 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r40 18 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r41 18 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r42 18 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r43 16 21 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=0.295 $Y=0 $X2=0.24
+ $Y2=0
r44 16 17 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=0.295 $Y=0 $X2=0.472
+ $Y2=0
r45 15 25 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.65 $Y=0 $X2=1.2
+ $Y2=0
r46 15 17 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.65 $Y=0 $X2=0.472
+ $Y2=0
r47 11 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r48 11 13 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.675
r49 7 17 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.472 $Y=0.085
+ $X2=0.472 $Y2=0
r50 7 9 24.1851 $w=3.53e-07 $l=7.45e-07 $layer=LI1_cond $X=0.472 $Y=0.085
+ $X2=0.472 $Y2=0.83
r51 2 13 182 $w=1.7e-07 $l=2.71477e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.56 $X2=1.62 $Y2=0.675
r52 1 9 182 $w=1.7e-07 $l=4.65833e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.485 $Y2=0.83
.ends

